PK   ��!Y
O�+.  �    cirkitFile.json�}[s$7��_Q�_+��~鷱=��u����F���N+F-��el���}��*���Ld�U�L�vǶ�HI~ $~_����o.�ۻ�����������Շ���%?�+[�>]�\>�^��.��a����{��ۧ:+o?~���o.+Vy�U�լ4��&����k��u��%[��i��Rت�k�9�u�$Y!�&c�禬���䫟�G��#=�:/�w<�M)3�M��TY�oj�U-�K�)]J�*�sɌ/E]g�;�\x��,3c]ř��WU;܄�cc�oT���e��Ɖ��y����WF;�\���K�G�G�Dq#F�YEzV2g��:�+�g
~ͼ�)�J��0Մ�5m�'�¸�1�(�)H�{Rז�5�ia�|��XYXU�:s� N�2_3���7���U��. ��c��sL��e�`ă8i�)={X{��T�m@��:��G;v�Ym��8���nU�̕�Ѱ��Mm���k�6���g�x���z��A�9j$� F�q�y�uVf�&�),$S���J���q���6��iV��tM���J�vܬ�uN{=nߠ^���cF
�&�7RP���qK�z�Ґ�U������GPK�̚�Ŕ�Ʊ�v@�34��&/|�Y	�b��
h-+�W���0�h=G��|S��*&o@q"kTVlg�� M���s�x��6�uSL�+�S�xX��c`,�TׂK�X[4�%vM�m���E�e���Ǥ�����c"�b�؎��Ȍ1F!��wMYyS�Q,��r
TZ��)��1��%��w�~���EQH��M����@�h�S��������eԇ�D{EĔ)
_�X�k��#�Q��ԧ��0AT�"�AFF(][J�1��uL��d���QK�5�e�ҲZ���w��68��e�z5����#c���i]S=�X���i�--IT�hiɸ��B{|E­�'ؘ@��b��M"j1 �ɔ�/a#�4^��h&��.�a���*�z&�%m?$�z"�?Jױ�k�S��"v=-��t�N�E:�����~ct�g�SP݋��A���˘�c�<����eu�K0Ѵ�D�+�7,�!�E�Z����`��ia\פ���?��5��
GuM����}4I�!�k���fT�$|Gͨ�c�5��2CuM[xhʌ�pN�f4���I�q�:#i�hD�u4A�5I�EtPV�D����3r =c��z���*@�����*@�:�U�z��uL��z��uL��z��5	���8R%��mnƬ$�O�:f%aW|J߱���S����X���7�I
���$�F�gQ��1F������]\z!2�2���r�"I ������2���\Na���R܈��b�����v8��\��g�dɨY�㛰'|��6rK�2b�]YL�_&�jLi�
|s�g�,M&�2���E<.��8��ӣ. �oB�$-���ul�HI�H�I 9�X!���v,W�;�62��[\��"�9-�#C�s(��I���m��py{}{G<+���i�g�4Sh��?�VĖ��0����x���^<ӌ��!��"�𢶼䵭	��$_d�/b�֊Mk[�U�SF�o�[k�ЇF�?	{�30�el��g9�y��������4/�3���dU�!�2��<a�V���ƞ���X�2�]乽��*^�)����e{0//&I+��{Zo���bZ
y�nZ}�O�%ޢ�k�dN���֍��f����4ͤA0Oa����)`��Z/�
[��J3i��H�bѢ�֢�H���$Q[�Ι���<	��I��lQ\;]��A�(�,����D�D�b�
�hJ3it�L�b�F�Y]�=�Y�{
e����(I������5���=����Y��=R1��Ч#fbȳ
	Z�u*�� ��[lB��)���_dU�0�f���8Yɂ��V&|Eh��䕊E�y�0G���2��X�*�v.Xn�'m]�/	w;�7�����V�Ʀ�wM�I�"��ב�A�,i�p�T�b3�W_�s4ܴ .����Zt&2��vD��F��06�xZ���������ol�tc3r��M���/6Ov�ؔ�i�b�W��6uZ�sJ�u:=tZ�3=�Mt������6"�ٔ�V63r�D&H΄��Ɏ	x�9aS���"Eج��̎6Q0A+|.J��ߛYg��t3�&df�v�Yn�)6amf\�	d�.66lf#��5�6Uj�l��t0��4�6�)���Xt��?��Ģ����.�g�XDoE̵�N,��2�E��"z+2I+*I+:I+&I+6I+.I+>�f��N,��2+��"z+�������N,�����Y5�N,��2�E��"z+���XDoeV����*^tb��YŋO,J�L��4��i��� ��A0Oa��<�y�4(�tp�4(iP,ҠX�A�H�b��"�e�4(��L�4(�iP,ӠX�A��E1:����,jЉE�Vf1�N,��2�tb��4x�Uz�Ģ���Za���Ǿ��E�V�c_��"z+�/lb����6����|��X���4�w���E	�I�y�X���4�w���E	�^ϻ`��"z+ix�(tb��YqB'�[�&tb��YQB'%@]"�A��z�O,J�L #Br��"z+��:6���ʼ�M,��2�b��̎:���ʼ\c���c�XDoe~\��E�V淐��E�VfyA'�[���XDo吗?��>l�+���~]�q��/Ww���뼬�˫��ۻ��[���p9�ΟpY��}S.-2���AJ�
���u	�"��RH��kډ�X׸J�6�32Ʌ���L�9cў��J�t�hGzF&5Q�嬱$�;��-�G�/F�9��'�vT��1ZJ���sd��n"�}���I]+Rp��5��3�kڹmRפө��&���1N�u (�H;#��c�(���i���5E�q�>��3N�guƣ�r���I�)���MS�|�w���T�����w�gt���Í<�@�:�b"�[��k��8R״+c)]G��a>R�"ZQ���DJ2>ʌ���a��:��Ty�jp:�ͅ�q^4q��ʺB��{U7��56���yE4j�Ꙇ�i��:�3n����v��ϱ\��E��=ZRה����:�ve�gJ� t��h��w-i7F��H�P��XFg���>I�(E��U���B�[J/X��)ŇЕ�(u�KV|��e4�>�&rc��%21 �329���Q��8%3�4�/���t���������?��2����5~&_0g���=�b�ƞ���_.�#�Ď�;p@L������#�c��s�~Ч��B�b&];B��B&8GzH��ˉ�̂t�4��)8�Tgi>~������,�3�!�f�̍�y��s@��I�1�'�ܞPS|�@����@M��s@���s@M��s@��s@M�s@�	�s@M�s@�J��h�B��X{��!z쀚=t2��DD�b.��� �R��bf��8�&%���gD瀘n� �H�:��"5��t@�� Mrp�T$�3��8Cb��8�LMSJ�1[i�><C��D ���ďΑ<uBmx6��Tq�G
�b�Ha&�#�y �%���1��� 1�l��3��M��3d��N%���g�\�HC�Ð��6��.�ц�Ȋ;Y��7��Yr�&98G��, {�Sf�Y��I��^bAL@}9�0��ٓ!2���n���=�~�����=^U�R{��K�C��c�R m�]l�[��g��*��ȴ�����!�E�(_g��PR�,�7d'�Y�-��k���6��h!Xl��^k�-jtվnk�����}8�����C��qI0@W��q�.�
��_O*(g#
?2v���G����?��ѵ�(�Uzl�D����c��O�ptq��pȈ�����k��N?�f�|5� `��X ]	�$��� М�hN�4b:���E�p���I�����U'*l�P+G7���H��ڤ=�6n� {�E�2�%{�Q�9T�2f-���ڣ|�$�!COS���T�-���T�-'7�0 �}|,]�'�]$0!w#������R��@W���W���8툯"�k�r�!qsx]`��\lmGW�5G�ء��"�as���X�	�҉�C�rjc(e�tc�y$����`в�GV�1�� �����C�����h<懒��P>b{j����?��a�t��� E ���k.�/t!�^s�����k.�=Хq�G�H�a],}t�D���{�Q�X��%�P�P,bz_Y��E.��-�`��[�[�(�1�nQ�ާ���]v�!{l%F��!47
Dc��?2:1�[�7:���C�dı��������i�q�����.�ÖmD[���]lM�rD���c��X> ��#�;t�Gw�b�8��U���B����"ܡ�@v����깙�*d�A��!�U�z��*�>3���d�t_Z��3,FA��f5HE[�c�I�yn^��t^���t^��`F_8:��@�*��ӚT����E�Z����Zӭ��Z��'�z'���zQ�Fy�k� Yxk�
��F�N[�U�2�Ya"�˧�P�gȀ�ٗ�� ��4�.L¤}��w� �w^�,���VW�I��n＀Q��j��i�c �=|o�y&uaK%˼��%��
���΁���Pږ����͖��*+Wd���Kt*�׵�\��[J-����zT��\U5�u��2o�ah�� �e��_�4yoYl6��
$O�)��u-3мa�4'e���UΝ�R�ʗp��XB�y�%!��Ε�5jG���Q&�R �2��K_ˢ*��%ss�d��A�J���VΘJr]m)�⎗���zkZS��Ð������氼@3л��k��2�)Y���ӈ���;V�ȋ&s� �,�fK���0�����yΡM�HW� �`��+�[JX���0,�����k ��RãҴ#���v����*}�{�ożI8�p���tP�T��Mq{(i��ؒR�)����"�RP���|�|��@�0�("�g�Y>�N�pC-c>ܼ�pC�l>���pC-v>L��ps�����qf�R}�ěvM3A�ލ�.�1<B2>�g)�=���3s�B��
7�����
7�r��� 
7�
�ý.
7��í<
;�:�ÝJ;����mX7�j��=f7���t7���� 7�2���7���ü7�b�ä7���Ì��#p3&R1]|�*��[�WA��x��vRv8
���<5��GC	�P�2Ӝ)n'�R�0�� ;���ô�ؐˠ�(�P+����P���q�P��"�-�3��l�*��ԓȰ��p�0������i����L6���<��e�L����yQ_�}&��Y�Y�g�p�������#�{$����>R�Gj�H���#�{d����<����#�v���o~4�4~5�5~6�6~7�7~8�8~9�9��������g~�L�L�L��E�E<�a8.b?.b8.b?.b8.b?.b8.b?.b8.b��b��b?fb8fb?.b8.r?.r8.r?.r8.rϧ�)��.��.��.��.�� �� ��.��.��'�ߧ�ߧ�ߧ���
%���,��*n�P�������z�YViP��''S5o��ZN�̹i�,*i�Ⱦ�����%/�����o�烔��o�k�{���w��껇�:�_�n��no� , �s�J+�Ίu�6�I�A9J#�uZj��
�� ���-��5���BU\��N�V�ݷ]������!�)����֫ۻ+h%߲�j� Z��+���7�o�~�����<|�)��Z0�<X(������FE�q��[6�q���ᱺ�}����MH0�{���I�r���k�k��܆�9����(SdZ�&���g\��]6J*U�B�5�D����]���p�50��Bi3��L��~�+���7|;3.�}�J	o��. l7���܂!�ws�B��n`I�},�T����1�[�v�Q��C��ya7 ^R��zF��r+�<��9��jxl64��=ӧ��b�v���jc��A���9�B���f��o��$Y0���kx�f���V�̩����#��!z������YU���γR��a��E����A����Z��6��s�f���O�(��f��ƀ��Y��0��#�j�I����{08��v-m�A��;H�FI���*K5Jʴ����T�O��M��3����n¿° ������߁���c�=<]���_?�������ބI���u}�u����n���Wo���������߮���ow�����a��f�����<6y��xW�M�pH��˻O��?���&+=�����w������!|��UL��U&��1��:��\H|P9�}�<~14�08TZ��-���#K �0��-���z�wVQT��ec2X-
��Z�`T&�*^��iמ A� �T~���ɰ�ԷC���0}��`U���* i}d�o��[>���ѷ�����o��[6�����}��o��[*��y�{�*L�pZ�d �HF�� 3B6��1 ����j�l`C�Q����o�l�#dc�!��P�d��!���G�ƀ=B6 9]�+ɣ��޲rWup	�ʁ��+�5��J�<��sP�:���E���0sOћW�y��	�Ɂ�0�G|���5#W1����#�C��*gv�bߋT�o�D�q83[�P8�)L�lk�2�8��������}"��r[�W{�3�d	F:˳\������x�ZD��/7Cs���h��/�[hD�>����N���Ё���n�l��UZ���	b.a�w�-�ڡQ��v�Z{.�ێИq:ώw�� 7@�M����00���{a�\�c�%4[���t��k��k���S`��u�P�� {=M�DKg���c�"4���3����^�!�b��9-��c��Z�~�7&#t!T����q4��o��K���B��$w~K��ל�U县'�OU��=^=\|wS=�w�CR���o8v�I�XK�A}+���
��]�p�)e��v�m@)6��ȋ�Uf�y�����u�[��V�[U�J>=Q�IWOO�1��'�I�>������@���"��f��o�ÄOD�g~z���I��������h�`n�!žs�̓�ۿ�L
H�+��Ń4H��L��#��n;�+)Lポ!��Yn\�i�]�L^�"�J M_�	s�\io�>q����+�d�����c���s�	�U-��}V`��D44x98@ҁT�p`���`��/dm#q>���h��F��BJ�=�l����tgB����/o3�Ӿ~}w�W�9'0Ԇo�&L�b��O�)l-y-�R�6D���F�ZUa�Ģ����D�e�E�N��xo�	)ֈk��R�4R�����J�����+,�MÂ�X�q}�U&����-R΃�w�Ͼ�o�������W���?ֿ�`�L��O<Y�k��"h(&�Bڬ�)h >T�s*�vj�|[ ������9�3��ζ��m0@u�G���k�����o�}�9�^�B�=�F?�e��;�q�ٜ�(��r��,ϝ�\ä���������E��V�n*m�b���g�ǿ�m��-�2Nb��n�B!�u���h#gE�g�1���"�fc�}^p�;��@]E�A��� �X�O&�</��å�\"��⹒~��
�8�(�����)����2���r�����:�A� �����bE?@�v���yz����W��G!&�#p:1�{�������]}s{י��>�^�wW���������� �O���z�\_}�f?uo���>�}�}	�)����}������=��33}����i�?���>�e���:�S=u�'�g��??=�z�i��ۛ�wW�S�����QP�s�E[:`��G������bop� $L>�A�rDz㙷�3)4؃�l?�Q�k�����E8�dfx��!"+X�|ԥ��k�ل��o��EF?_�/(��n`�t�3%4s�z6��̀�^���$B����	�W�qu�����"�����Q��Fk������؍9PwE]������]|�����_�/���(�/��
�6�[g$���!#+�C�&'��$r�����������ş��\\\�}��鋸~����kjH���Y��p�	�Τ�x+���<��4k*���+����/"�������{�zC��P�{%י�X�<����s"E�xE2���~�e=�����S#����Q���E�z���s��IDUa��ꅺ��C~s�__�����"���������l�^��^hf�Zi@��JXN}8�uAE�zE����悛_�ŷW�����)���U���^�p2Z(�V�m`9�6��0+O"���r�HP��w������×��g)�/������pa�2�q��ڄ$J'��[��i�P�_��>�7\|_W�_�􋜞7ɺpK�r 6�x'��^�x���1���20uU_���}��p�������!�"�gND�L^a�v���~�����J����RTI�W$�~��B��/����:�ᾅ��MBR^[�v�m��`����`N��*$���� �>d~YH?GA/�ڠ`��ހy+��\[�7�(�
��8M��Iٔ�-3k��T�,g%�[�*��4)2�yp����- ~�I�7Bl�j�W>��<cg��~��>�&��V���?~�ۃ>!m0�W2������o�`�˼�PW_?U`x{W?<������aR�Ce���À�ޯ޼���j��G~�w�]�>:��}�Z}SM��,L߶u���.)s�������
W��m����߯Bы�����V-߇���)����E�˃��T�M��`��n�Gw���na�:w�>Q���-X���KLqߣ����_�H'�U�L�0�+���]��K�[ك��Y���#���i�	����!$����|�Sr!�����ׅIT�<�R�\�ݿ""��T?�)uY���MYh���� .�� � @�U\��/`��-n�l�`֝գ��y6Nf��
I6�48�?s�@U�]��eK�<����ϲ��6�Zi{d�j`�3d�l��/��*�y9���:�,��NO����0���r�\�������]�I%^�^C�n9-`�UaH�q#�1d"Bƻq�!�+�`�%1�-`�_l}�G&X�bSǐq�7B��=�E�����ӹ�eV�:����2C��8���9p`�^�e��8p��&��C�ڍ���Rg_��w����Ӆ�:�^Q�y�������^�=1MdG`�L�D�� J�4m�	5�����٪6x�-`-�F�9hϕ�V#�#v&�Gv��ƙ�n��}tո%d�1T�=�PGj���p$"��Ve�S�F��.�ni!�R��ni�����88��#�0�����2�x��z��*��A��"ȦCВL���B�q�=u�.?ͧ9�j��{TjW.v�Sa٧c��n�O� ��.O��Aأ"H�j厠�h��R�x*�
uZe�A	=��:(�c�F��(T�L�*�]�KV/��ꠦ���X��Ue�3�}��ʸ���g%�M�dU%�A#�� ³�
?�������#�n\�0��
�ݍў�cЇT�
틨���ObLV�n���!.?0/Z%8���򅨳�T�m���Η�!�����:���L�&w��g�vYs]���'�)��>ոͮ��P2��{�P�q�0�L��!����ZL�7��b]"k�v�D'ҍ#jkX��Vr_H�+�� �RK���Blw�S�x�j��P+x���)���9���Y^	�F�5�Ƅ	mj�J�_�X{Q��D�Y������8rzD��Pm<��E�g8��v��P]�Z�}ɣ�ק2h��7���������(�xpT|<�"�TB��ZZ���{�P� v�D&A�L�̤E�<��Ӵh�q��Bq��5��Q�=:m��QF.�����+�g�)�V�ۦX�b�	@�3�� vv��L9>.2����&�֧:��]0�I �@�.�$�=J��NӢ)��E��o�a|sDD,p?/n}*��e,��1t�S���1����Q1��5�bҺ����6�
��M^),.��j�+��MpO�/���>���2ܰ�_r��t��c	o�����^�s^;M&��]���Ȏ��#��w*4�J��;2��
;G��ɰ&	���������"R�w�Lu/�i�@%�%D}<��8Y�")��~fuj��<{K��(������Dm�",���r���ZԸ/0f��
�e P����n��0ѣ�A���.)$�f�yrU�w��8�Hl�����jԧ_i2�Y��T� �Qqc�`6�B�5��f����H�&2����R�[
4�Y��T�i*�3n��V�O7b�?�E|AXhoɠqT\(S���O�t4���O�>�7M���ƥQ��~�txK�#o�Ci��ڶ���$4�THs�v�
�~���/H�^�[2h� mQZâ�FK%�s���S�QT�Ag���y 5�N_,�-4�;}�,ƨ�QE����8��Xߞ�Ǩ" *�K�[Fwy��n��.?*��q�R.}���¶���e@����J�mL�$���ܴ\~T7��`�d1���TL�,��]�v�s�!�#�4UR�9a0�/��X�[2�y����"T�G���ɰQ�ܤ��u�\ ���d�8�&��}��(Yl��6!��i��'C.UVUi-����NR��H.�kp�]����"��l{�:C��.�
�0v�ڛJ�=�({����9Lv�\�^����@�d���9�d�����.��E�Pw�'���[��R�n�֍���b��2�����액gN�����(�ݨ�,vqk��Ay��
Kƽ�����YX��;�`r�D%��x����I.&>�����e���P�zk$Y��b+�!�^%�4�I�$�`C-fK�6-�-�Z{ܦYO����dƯ�,��;c��*�I	\��R��\���2�C&"Emz�@�E/52����Wh2���)|���F)$�,�-�Yw\H���q#�T|�V���%k1����Y$�Q�
M�Mg½���O�ݻ9N�����W�E5~�P�=����B�K��܄�~���8la�}�2a�Ԏ�L[ I��#m�1dލ�P���xK��2*�YYV5Iըĭب
��^��G�����]'$�W��{�IA�C���G_3���SG|�\��g-U���(��٠Nq�,b����ٹnzG^�����Z	�o��sGs�_哩��]�9����sl��V�7�)أ�{dQ�&�d��J��'��E����Z/$C�Z����zے{�A<I���9;O�g�!"�zI���?�G��k�1��NK���r:2��	t�d�4x��n��w��>�u��h���E�!����Eh@A�*d�����ZT-��*:�v{DW����{H2	���E�8�ȕX�pǐ�ߟ�R�2�*r����Uqu}�C�����ʯ�Wo���_�������<��_�~���x&��?V�/PK   ��!YG�~��  � /   images/0739a1b1-a163-452a-a325-ab452d55b136.png�y8�m?�r�J�M!*IY��Ie�^Y&������[�d�cb�0��d�1̒,�ٲ�L������������|�|�4}��>�r}��|��mn$�_l��mۄ�o^�ܶM�i۶]&{w-�����A���{����� ��n�m�&�I����em4�6�l����
�*y�����x(����WŶm;����5��9t4Gb&��Ȳѹ�}��OܜΉSٱ������b��MT�}�L�1HƸD���?j��i͘�ǰf�	�A��{�ξ�[_����J�z���r���٢w��/5a��t�I��ե�EnhǶ-?����'m�ں-��Ǔ[�n�-��v<����xN��J�h���e3��2������7��=V��)u!";G?�� ��<�|K0�yY���I2,���^)�Ϭ���Ev�p�����������d���4���dK;!-�L�^�$Cx�䐦W��k��E���9謗	* P��ϕ�����S�����0C���~�?��$Ǖ���φ%mXJ����{���w/�y|
�T!��;��G����쳄�[�����⩧�U�6}3���6��{�[$��ab1�P��~z�3������Y�q(�V�f��¦�&	�� ��l.Z��s9�2SH�W�ơP6�[��SnT�QokF!s�Ǔ`��� 6rl�������fI�:�v�K�|l��%����)�m����}gw0�6=y�dk��?�/������<�w�}l��جJ���s�+����������6����Í�͍{3�����"R-33�	a\yoU+����̡-�߶~�S���v�ѯ�f��nY7�߼�K�pE߬�����f�J�\t���+"D�,�����AGf�H��X��i���&���oց���A{10�^���l����UL&0���ٵ?���E�)�Q�5��s�=[�,�8�v�Y����>\��>\+sS�N��88y��</�!-Ot�HS�/'9��q�ZwuR��
���ӝ�v�����xS>edf5�Ի`��Z��/�j�3�QM�/
�1Q �wH����G�h�p���"[�|���fi�h.��-
��f�:�[<?>gh8)�2d����q���j�GZl��Ϩ�4.{��F���Hq���5�1͸�m2�2~�l����]I���J�&k�-�x�T�/�O�z�5�k����8��JdX��a9�<��V��\�����R��9�����0�TƦ%r�hm�[o���b�Pԓ��YپQ5Y�� �>[Զ�f�UG~����bhA�A	���6��,-��:[��Y����p���m���k���A��p�ʂ�K��&�{sdJ;?=3�O�	}�Ij�>>wE�Ws20NJ]=X�uq�g�j����bN���|�G����Q�s˪�r���W��ӕ������7�[����v�ЂF�K^��FY�{��s��ʻ��R�:i��D{��x�����T�Dr��j�M�s3�����:u˙��[�.�[Im}�v8��0��d�Y�S�ܷ�BW�V�F��V�E��V�
���355;����҈�RW&/�+�'��]W�e����v�@$�Y��=�Vܲܽ��ٳ�6�tinb��[s!ޞ�C����<_��iG�Gn���_a+*�� ]>��-u��{\lrǹ��x�|�b�ߕ��?e��@�㕸�����[�`J�p-��i��m�'���n��:l�xm�pd�l�em,W0Q�:��"�A�fXDyP��pOTG^uPiN��c��+l����~ŭdyώ�ȂrZ�����?���A�Xc|O���/�Pc���>���tx/��g�N8^xai=���
\�ΟNXi��@�l��]Q�0��!a�+ץ���q�����`Vq,�o"�B8a�i���Itq�����1C�06�J��J���
�<-VTy�����kQ
�ɍ������p�F����Ϝ����r�}��O��u�~�Ar�u�����Wc~2�ƪ����@�m�����
&�H�;7��.2g�>)l!�(�|�v�z��[�TJ�й��#�J�:F���R���:oȼ�>33�w��vå"����P|�?{�&��#�H��+���#��<o��Jڐ(-�������&�Mt^��R��|٢����q`�g��c��j��02���)����F�;W������+�xR��:P��/�ސc�H���\k�Ý�/���d�����^� u �Ƚ���c��������-6yK�.�d�j��܉�x�������7�.{��"�'�>����K�۰o�g����m%���UY�> �/��
zo��X{_�v��Kû��q��Ŧ�ү2#G�_Z&�k3��x��r��2#zל���@�[��װ��^_�L�#/=lql�X4Xm������nq�p�7ME]�A��J60��e��ogU.Ė�FՄ�W_Ћ�[cT���l�hze< &��x����/{�"�Lv��
��= з$:��Ln�_�|_�!��ɬK{U���G��Jak�6����������R3Ć��S�ۿE$��|��ӝ1��E}��q[s<w�R��.�$����V�P���Lկ�0e�YK�9��qO_L���p��Tu��/8�ˊ��Z��]��A�@(�^�1���s�z��'�l��x�}u��A���<�� m������j��1õ��B��iB��	�A&q��6�t���+�cQ"M	��յN�I/&�'9�˹��Vv�t�R��FAD�/��"������N��+�',��Z.����xT�;(a��C��?����Drɴ��J@a��m�e��h?-����b	���M8=�^����=�ӽ�b/��Y:#�3���rp`��$G7��0_��s�N���vo���B��
]\�R�	�e�1cٝ)z)A���۹����E;DO�V$���t+˾C��@;�sA����.���8yQ\��Gwz�O/9s>u��ř����e�5o��e=���qפkx�t������]�o�O��V��f(�\z/�x�@P�p8��R��fU�j�nL�`v\�\fM����qY�cGr�?�������@�W����:��7[�zȏ����{�N�ND�v�bKT�
{���=��s,�{B-#+�Vx�Z�%��/�(?��9&s4]���5���3\>�P(y
�6*���+����&�sN}wT�$�8���/Aa�ԥ5i[����x@�� �`��������4�nc��,��R���1��q��a��­��[C���	�~n���7a�F��G�S̻1[�#ݹ rŀ�}�uNʂj*�6I�VU˕��UP�����h�1G�2�Rs���Ծ�y[�J�梵3d������A���i(Β�����~\@?�,�8�(ݙ"�i��ݤ�܇^��g�ms*$��ESפ�#-
!���U	�����lQ�̵��K�1u)�ױ~Q ���16������	���8@qY�&C��.:!�6��;c0߷s� ��g��"HSK�P
��10ڂ�|���}��([��`�d>�*��I6�c)<���H[Y�ғ���,~ �lvЧ%	Y�m�[��>+�8U�t�@�e@��v�AB�a������m����p��_ \�**�>j۪��q�E'|���s��}��)��Һ���w,���n�b*� M���1?VPg�>V{���M�|j�:`�@�������x��Ox6���Q���s5��I�a��P��'��C��ݽ��(��/(���Y�<x�̶H|�d��kѺ>�Y�G`���*"�r��l��$-.���A@<��E��u�#�n�����,�=�bB�B��^ͧځ[�<C��^� ��|�C$S+��G���.Ԟ�*��� AP�	�oe���W�\t ��i����� �D=CZ7��<���?��1����m!�����;ZЮ��|�-����;����ٱ��rO"���_�yF�
�`��!�;��U��X���t��(�JW9�~�#&�M���j�n �I=�x)��s�Y��rvHYF|>zBf�؉P�":�m��'(����n�?0 �捻Dr��Ox@{٭�Qh�BU��_FQ��(p��
�zk6=U�E��+��2p����v�)��Y��4`�n}��Ƕ��.E�Tes��q�e� p3I�k	Y�պ��ľ̫�}�Q�@�i���u��<��mЭ�6�e@x~_�"^X��$Ԥ����txY��&��_�/薳�q�1:z�3#9�Sd��V������#�����m8./����V+}����� ��jm�*~Ԉ`*P�,��\aK ������=}�������1�c,��s��E��J��3�2doR0�e��&��}
�)@h��}�G,;�`�͉BJ�Q��ib�]M%�%ᖝ�$�3���0f����9��.����l�O�u+6��,w\μ���� j";+k�Q@��7�HDi;w��d�N�Ž�͊�BX���+z���I��Ӎ�R��2��q�:�r��Ť ꛕ�4�J�\Dt��>w&�����Q�)�,m�k�b��	�KM�PA9A����C�T}�v�٥M���dҊ-"�Ҧ�^���o"�.��Jf���Q�^#��B6��&���(t�f�4��g~yŪ�Y5����A�Epq�3���Ĕ'�Д��*�AT:Vb��|���-%�uw�e�I��UU<��2Pl�SF�׋���t���ޝCɶ]+�7���Ld=>e�_�T{�+�F^Tx'M����DE�o�-l���P�G>���Ѐ]
�?�8a\I��$��B�Aِ�"�n��P�j�����Oy��eDH��t�k#�AX_�&��O�-���T`g��JK�7J��"�Ÿ�(64U��]'�YP��D���я���rZ~�xy���uu$|�2���d~���a�sa�w/���������&���5#k��'+��}PkH,h�d��v���Tϴz��Z��G�_ZN�ad$	c���Tx�4�nʤ��6�P�����ʞ���|�uxP�[�+l��VF�߃)��k�~1s��Q��"���c&�,�Ƶ�ͦ�X���ϠoC��l�I�v�$Fc�I��2!cY����RI����-䋴X�Za+K�k��Z��\�=�Y����n4a��gT���SQM����܁G�"�]������ ��wl�q-��/\y�u��f�ň7'�
�l6:�9��#�!X�Ě��b�����F����w�:N[h�[�n���=��C1;����M9"〧����;/Quu������� ��N�ۖ^$b����|7���V�Â��a��s�.X[�H��M�K/�evTv>�U۟��gSǄ�E�|���Hr2���}U{9��y,{�hh����y� h9��&5�Pg��X�s2� �b��ͼ�tzer��;�4O�+NfpE/�ݔ��(BW��r���9����(�oB6������픴Lq�K���xRtJ�?K((2�~^>��npM��Y��#�)a��ݡ"�#�|�a�*�*�j���[e�G(>�D/��(�|y�W^ x�m#�]���h��0T[fLL�j�~Ԅ�jo�u��9���p���r~��So��}�'�ť5^LP�1��
IJ�p�C2�����IJWC&� ���/��\���=%ݰ�){�����{8�ގIR�v
�Hp*Mi֪�X;����SAe���x$��V+<�$���s��\~�z�}x_a{�x{���#2'ͳRl"�/=?�z`��V��s����8�>�ȷ��k��*98��е��zy�i��S�h�4�?_�\;���Yմ%�V%��b?�����ܕɪq�ꑝLO�t���RT�^d.��p�*�> '����'b�CU/$mް�Q�ql�[�3@��pu��ToV�@���Wz$�jIgg.��]bT��$%
�?�H��4(eh��Խd�,�m��cn��B��
�b�9�uLT3��	yX��a�*O��;۬&����Ⱥ�6Kо�S��`�\�˙o�
��Z�d���%�����隲��/�@,���z��҈��I��cW��f�HЈc���h�|���Z#��Rt�Kj��N�\%�����n{(�ډ<��3�r��AI��֞��C����Gz�.Zm���J\i/��I��)�k|�c����l3	]݄K����'�q#��+��?_v}c�1N(��ߡ��~5�(5�T�Ӥ�O�!��n���0{HMWǥ<�����e��ؘ298���i���|IT�VDb�*y�>w����$�Om�~W�z�n�W(���r�
�z��Kȯ���'�q?Z�X���U/7���3c�n���e�����հ���e��Ym����� DQ� &5��}z)t�ȩԻK����k<�q<�2�1���<79��������8��в��u�F�'Z{r��(ഏ�,5O�o�ܙ�v�ʨ���Sn)ړ	h:ͽRj����D��j<s���Y�H�5R��z=�B���㼌��a�}���UZ�6�@d5�b��	��sV��5�n��7n�:�m��!�'u�	l��1*�Pte�
(���l��U��<$u�{�<l��F@�O���Wyl�@�+,�)����a�
e��k���O�X3��J{n6�Z���G�6o\�]ʚ>��R�,�g.����{Y��ma
/0���U�υWcnI�*%\��W�+�V�`õ�x�����b"�r�=�\����Kmk�)3��g3���	Y{�D�}<�76+7Ŭ柕� o�|feQFW�C�:?��\lS������[7tُ`@?����چ���� }zY��E=	)?YQQ��-ח�q��syBk�S�3Q�0�w����`�ӷ��FI�e�c�B�g�Y���_���x��l� ������l�MҦd� v��q�P�>@_�����^ZiE>�)>���K=��*�ڍI�t/��.%S�B@�����T ��/��GJ�{�fm^ͥy8��ro�Vö�ϿNo����i���ѓ׹F4�6�>jY�::�zֈ�K8�Ϩ]U5�SX��k�<����)�Q_���ߙ�%���sY���}�Q��*��4f�d�Q��*VE�z�5�
xI##:@�t�}��+�{�;��$Mr�J�������/�\��1x��U1y(¦}]ĤwD~���C���ڣ�1��H{�g�d��4=�Qa���M��QZ���ը��fGR�}�\��8Ғ�q��}�4;l��/LoF#�T��7����֍1�ޣ���'-�xT�C��h*��-'�I��M�ڈ�s��/�_�{�����G��L��z�����,�+����F*�޳V�����>S���D�Rg����;�m�.V<�����3�t�`#����N������M1��nܩ�7��u&�]�{جʦXO�k�௛:Rg�L2�4�Z��O�TS���q֟[� ���]�h���uj����X|��Vmwa�O��D�����K6}���n�Z��Oe��b�u��2��A�:vq��L�J�� C"<��Z��������������;��X���H���[���jB?�ݧ�#��Lr
���-T:�+�D֗��@�E�ѣģ�|Qgp=��F�uK�ܫN���Q��� B���Ƽe{\[7ҵ��H���n5֎6�~�b�.bצ�!�P�	�	G���k�눸������J�|������^B�^�Y�n����5��f]$g�(M,���D�h�t`&ȍ�f�j�7���xYg]�22X_7�����=��f��7*qKn�ֱhUr�Y�}$U��G�e��_~�T�1�;��j&�>��!��I�.�*۬�=��(��0T�	�GU�Weh�7bTQ=5�8�n��މh�\�_����+D��YZ�wr��V1Mw^im�G��@S�ɚ��� �w\E���Y�wStH���n�
H����v�.�ѥ�n�]Ux��D^����ї��ox�%��!�����NKx�#��:LۧYf<�0�W�z�4	ռ\agM�*�L��2�^caJˊ�:������Z�&���DS�zu`;%4��P���f�e�`�c�wH}�*6@v;���9_�ġ%�]���gƷF���S�T��0��o����� =^=�
���"�����P8� �ױ+^���#�3*d��T`� A���F�>�o�{�҅W=���ʾ�3�yq�z\�S�Ѩt����):/���G�*����fZ�5q^�3���XRg��X?��p�O����7p*�̄\���-��d[�P	M(�vQ���nS8�Z���j� 4!�f���&N!���[>��^������c���
��Er����ֻ����۠����q�c�]G�1}WUv仓!TE��d�*u��㴧����ag�1�Qz���,���R��yI�u�(֫�^�6_kk���	h<�"��Dk�y���'�ߋ�n�)�k�K�ngX,�h�{�]5Q{�q%��:�Dв��^ndH�P�m�R��
�>lB�D"�tf�����^O3�e�z�stX�g%����u�	��<�W<��m�Y� CDhkX�� ���fß�| An�G
�H��`�h"���L,���;/sC����HL��/�2mnM�� ��G2y�d�of��;���>$�����m=SfM;��&��n;	�,ů�)�Nl�]��3잡�.[;;˦��Ť��Φ=w�^��i^���`�#I������X$���}���L���l��4
��~Ti0�l8 z�Qٚ�(�~�y��H�`i2�>a�S��U.+׸��L��TO��<��u�@����#	�m�s��ӆ�u��*���~��fj�6���>�H+��m�8�B�������l==F���t��'Y����eo���|��$��tT
n���W�k#e��ND�\nB��.�l�,���=K?����p�|[��5��O �x5�L��z�L��Z˹H������ׁ�3�F�Q�Mr���4�4���2k���m)��4e0�$KufN���'W������L��3��̡���i��t��nQ�eJ-�X*\p.22�	`^c�9ν�z,p���ş Ɉn�}# 9|z!D�!J��W+�g(̏���\w��>�����	�O1���.��p���׹��\�h�(6�3��d'�jMk�XC�ݺKc�E���$K8s�1����m0�# �
�Cln�#z��gI@�gAЅ�t���:�g0��Z�2���	�1�6/L��%���I�(.-�}�g�
�)ޔ��}��_���OrV�^���xK(��Fe���^��"6�w9=��1�k�k/s�bQ�1L1ԃ<�)�N������uac?�{kQ���>��
@������R��m+q��j0ߕԓ���	&�Л�軣����b[`�����\�:��s	��G
�� q��H����r4K�;@��]	�D�Ӹ��$�����?�	W.@���)������%Eg��G&�Z�ɫv!%�h~�=p���~xjX��(�߲^0k����W��/	��kмj��P�
ʑ��Sv	�E��1~��R�)+L�
Y�� �P��E������=���WH�zq��{�3:k#� 
<.���?O��H�v���܍�M"r�I�c(��A�5�Ŕ����،�z٣�B5��~��tI��t��X�}�|N7pf���M�ڷ<fțP^�̙\}&�"׏L�p5
x�R�1yQBxV���v�T�%+�������j�n�	��E����#�}�z�-��S��G�=qN���P��76��2y�ɚ�����pQ�XW���4 ȤhS2P��+ZK��s؝ڛ��o�'���g����l~�`�f8)���>��z�����V��������?O��4��o��A�ΐ��&�d������^$�0��ٍ�47.V����9��B��OKH��<*S�����Gy�VJ��Eu8������\����)���kYp�<�l������'��|ݻ�NA~�ֿidC�量s�Tiy�E��r��x�?>W�F����N6a^����}̶Kn��
��-�����>��ݑ�O���ܡ~��3� �(��p85C���pR�n�{D*�Y�`e���zb�1�L���a�Z&�AE|�/Q�%н��]�d'�� �Vx���X����9ݵ/��t���n}"���%c�^�����u#}tD����@OK�IT���͛S�&��#7E�bή��>����գ�$?�o.��Y����DYP1Ёt��#��d �	�F�7�o�vؙ�s�5DZ��[ �w/�E�j�A�y����xR˚���cGe�����rO�I��d���r`�#��7�<Ʀ*Rv-:vE�ُ���?[��N�l�`0��_�����/�����4`0�Rp��3T�z*[�'�L�:��{e�]���z�	��*���I����ފ�j7b��~�_	���8�)��PV�z����D��8����Wdg1|�z� �(�߂]uB�p�:�%��dS8���Q�B?WE9Tt��̀	�ǋ�v��7��,Ö���ip@���ڷ��U�s�}sk���c���;���r�>l ʾ�����K2����"\ف�{>�!3 E���o�.����7��D��vv;��Zu�b�&(��_��eD�>2�H�TA�E#��s�"FhAb@j��%Bm�@�Yz��X��'hN2>��������M]����>�T����.��ʂ�`���<!`B�ju��`5r���`"��$	˔����T�F@�m�\�(k|����;c�XS�D*�}{�!ODC!�x1W`G����a�DG�z��B0�;�]�!� �q�F����?�8K�I��0͠����0�C�0\{�>�'@\�Cȕ��P?z]�*�1���e��C>@2e_���(U$���#S<0N,�t��i�;������'z��'�]�cDm
D��#+R���_Պ�����a^�����J9�
S��%t�p�������9�{�F�N�ǂ��;=�?����_E����g�Z=��;��4�2 ��)��\~����"36�(��C� G�)��T�pN�s��*?O�͂�rd�Л�_&Ϣ�{���vX�v@�;Iϻ�^��tP�����p�?�CG������+�D���o�s~����~ߩ�Y0�4��  Kn	�T ~} T��a��u��J��}Wn���NRVՓ�v��#]��9ʂd]�,Z���̭L Ț ������E��,�/�DM�/}j��HI�O1��س��m����N+?v˶	o�LQ��6�W��@\e�p��uZ2+7�&�����~!OV3�\�Q�c�0۴9����wN]C=��%2�N�b�|��ׂx;����t�E��4L�+��j�d6�YO+n�YUMP���ɜdD�=`` TΙ$(I D�5��^8њR���d�e�ɰ�}v߸п`Q��?��{t�LF�/��k5�Y�#b������&� �iw
:S���\�Q�vQ�a�(��Ͻ.�%�X�z\]��J�K4��}��<�ư*9��isx����?{�㕙* �(��z�׸��Us��:^��]V3�M�߼?�g�皖���rS���jjS�s�g$�e_2'o�G$�����I�w^��'Ӻoh�"��^��W0��rK##��9;y����܅,I� E�ӴMa�sv�!��?�t��� jG�7ښvD��΅�����t����s¼�0�������f�t�7��(}8�"�>�����7��fTP�Y���ٲ����A�T�t�]۪�pq�఑$JF@�@m�M����]��P�7��}���˽S��@O�!�ҵ��n�׹̈́K��X&)G�m?a�S�U#ah%��	��(��+������Gyw4�L7�E�;�r�\1W�}������Rԉ؋����R͚C}Ύ<���:<�����q�\����	�d
+I�~y�<xxQc�F�&	1j�6J¾�8���,r�z�]�U\Уv��.<�M�]���6�����I��B0�a,�[-�����C�o�0�qcè�����t���m��y��`r����l;[��j�7����_�:�����°ԝh��l�k�^;�� c�eIv��9�~}x=a�{R!w&��ݒ��b��v��gO�����\��:ټ�?�[Zڱ�i�	$H����;�\3G�s�k��"h��]3�oz�&@�NV�	B(����s8�WuM���؀zw��(eJ?����,͎ø�o�����1/�ʙNك���A�]>?��bby�H�������OYjŝ�.~M($k*���AD����9.Mn�w��sۭ;��WJ�u3�j�o���� �8]�Z��Ͳ�`�:��� �1H~kȃ���h�g~ã �m{�xJ�}���f�;_^ܽ��<k��>m�&p�h�������1SEi.Jƚ� |N��0� �#�i���_e����{+/"4jS��O;>��g����rAlP������/>àÛ�Rʓ�`��r=����*�U���G4��_fx�"�Ǳ\�X�A�9۱n�5���1��kЎ��y�-��9�1t��&�=�����hN;�}�.~7o�qU�+��照E&�V8W;Ͻ>{PB��ދ�z&'�������	���t���LgO
�,�9?{����@��`�7��������!���[�ʔ��H-20f#!)�99R�4]���IQ�T��f?� �o�3��>�%X0{�}�R�2�GK�W�5�l`o�AK�4H/����dwh�>-�)��o�C��.�r�C�f�����^�b��,9Gc{,^�9���9�u3����o���&�����j������-�T����،�=���t��������`�T����=q�����bff^���@�ԧ�m������_�ܱĂ���H���vr������=�q	7�Rg����_I�/-����|؛�>uɯ��BQ�o����Eþ�e�����A�!�;<�uz*}�wa�N�����&wr��?ȟи^�v��`��ԺP��͂�OB.�,r���	�߲���q��9�?;�Hs1��s��#�U�Ӌ��*��2�o
�n綱� �7g��J�-��u@M�q����"��ׄ�v����Ղ���vW�T�$������S���N�:~k�m��Tr��X?M��nU����a(��̅��o��i@��[����pj�rNpX��W��?�h�2�2-���`�W��/��*����؜Ps
�8 �� @��ݙ_�c���5�FL����;qA>� �k<~�Y屼�G���ōv�Y�7\/䃧�F�J�8O��.�Ҭ�w�;^���ӥ���64_�����
�Ƨ�g�l�N�]9�z�N$Pn�v6 ��ƤK�@���PZ�N����fM�*!��}]��`v����

 �)!���2CJ�����L���Ӭ�>��뭠7���;����@��egXa�3��ay4�w��)��/|)u�4��3��]`c4��<Iٰ|ԩ��T��Z�#�l���q���^�������<r�3{���;"��
Mw�����k���L�j{���i1ڕC�ch�3J6[�#Y�
�o�i�f�u�Z-�@���|�.�g2��L>�	����ʰX������HreA_�pw��[&�����_�{�Wq��pL{��U�w"��RMk����2�zœN<��>�4,M�z�B���~"�_�z|
j�l�T��Q����?{4�����~N�_�ƢE�v��H���ϩ�#��GO��M�/�֑�k�.H�s�>\s5��I�&ڇX�̒��g�0���u]^;��d:�����S�K@�#L�{�od�F�,H���c�\1sZ)5���u}�{B����L�5�?�T#^�:G�-z�u=�ь�FG�C����s�u��j샱�'��|��{���C���|���<$11��];����#Ъ��]4;�V}s|�f#���|НS��� ��m�J(���t55��E��8���K�=�)N&�}���U(�ׯ���w��(����;�%�RWu��J�Ś�I��~��KA��;OV�@�~>���TI9�cz ��*@���򈌴(��	������{��Ps%�n�E��轶g�;*$P��U9��5���_����wU������޲��*�w߬�P�D"��f��"��\v���i��T�ſ�D����'л�?�?�c����������!��*�r��Z۶�+����8�W��N4K����0��P�=A�Id$u�ߪ�-�S�y���m[�aT�����Kw��x_�ȷ��j�������hg����=���������7�0�4�1����@48�Iix��<$���1I��gb`/�V��R�l%��'�H%F���m��=����[��=N�\|��(��	/K���J��γkpۆ��ew���&��r�1�Z2���@`������lbj��/v>��y\m�@�J�0�,!�r*o��)<���QqaaÝ@	r_˦K�d���$�����k��m�=7�8�a��.ľ��S/�F+d�d��]���_���9K�9�ڼ�KO��D��sh�����=}|e[�K9{U��햲>���v���8�O�ʥl�U[�Hx���$��Y�/\��Y�$N����F�	}}P�!���==2�:h~]����y��cQU�ք+�5����LE礮ŭ���
�&3���O�R��u���`HUE����;��:(2S0���1�|�Z�RTW�[8{0M*���+Aj?���!nm�4��&��9���CO�ZF�v���|��.�^�kz=����V�ϰi��=�։R7�|�!hR�� �Ra,�7��&՞Q˺��.��#�vg}����2��B"4C��/�̵4�}�QֻXل��%oj�@�������h'$ЪX:p�¸�wh��	���t�'/e.83}���<.�;���8�U�z�������"���==���ӳ�?Β�:+���=u���oS/������U-���?ǳ{�)9����:}VL5�)���^��.��Y2ri�g1~��em/�{�ȅ }ȉ\�����ޤ����� ]g[�M��޹ժ��q��$�)]����(������)���0��j֧�Q~֟Y����A�yוGEwThe1/�67z�ظ�H�J(�''H��t~Ş*���Ҹ�ϰL�̐���!U��"�Y��f���g -����2���j̞�(�p��0��]���v�z؏X\���̫�=.�jk?��[W�V��o��C})M2_x٘��-����|1�<��JU��''�y����h�P�W�#��������bvM��e�����ְ��2~��N� ��M��F��ͩt����ʼ���F���U��y�\Xp	�Q��uչ�0Z�*�nԔ��;�!�k_��CN��x�E����PM���<��i�AՓ�"
����E����������^��7-�e��ƙd9ʇ*��x��JcJs�>�ԕ��M=�EC?x�#\I�g��3U�{7&��f=�Vwh� �l\l�h��t��+��
8��l�e��h&���7�<���)�'�Kf	����ːDz�r-m�C*d�dl�ou���"(�bV��_���d�#��a�4�`��O��%�lӑ�:
)����X�B*���������RN��
��sƁ��� x�)�+�����.G;�G���q�_����F�(���G�~��>�~_&�6��0`��(�[�\�N݂]\����t�?����s7^���//��s2�PK3��� ����C�FC���K+]�)��GCi�H��tG
���&O�ݕ�bֽ�:^��6�R����$�Ԇ�Ig�g���Q�ˣ�j�W�OX��W<�����DX|�����Uu���qu�	k�Je�Xpӕ9��)�d8
�Q�a�9"=g&���A4��wL�|���g!W�<�fJ����oh@|��|��N�`w�;{�>�r-W��nN�	�M"�}i67���#Uvß���+����eI�~�]�3}�eC �ؤ�qc5�
Z�:�z@��5(.�Ƥ}k�Zs����J�?1�7k����<�����xf�	����^���$U��.�Ս�7���7��q�gV�g����t��Mgߛz���j����Q�?:��������;l���0�l)�J@�@X��'��jwx��پ1`��p����~|�<�	>R-��鞬G�M$�_x�i휱g�i�
�7$ cE��ɸ~�O�T�L�I���o_����´�nI�y�/$J�L��ȆA����2�׿�F�GF�=�I	��a�_r˟ ��P��j��3��q�iL�N�����$��/r�J�o|���~��bMuuC��E���%�[�*R�{�����ĭ����c���όI����K ����u:�45��i㫴x���CM����8V/�,1 F(sa����j}W�I�{ZH@ڃ�NL��zxA'9��p���PJ���`|ĩ�֒�h���CO����t
ujL��Y�7�a����6�����w�o�x�3R��J;���t��h E׸���z���7�KX'�x��ڢ�ULW������ipw���x�M����^]��;:E1�b3�6��t�'�OB[�0B_�i�6���,���Y.L��y�ܙ�F�ouZw��O,3$m�r�}��6�>Cx#��t��8�����QM/_ߨ�c��X�
�DzWi
�;��^#��HWz�{�� ��.%AZ(!�����9�G|����u׻�k=�יٳg�ޟ�e&|gB�/�!�>��	[�^l�I��۔��<$� ��rŒǅx
-V�-��T����T��h9�	��oXi�&��I"���yEH�;~�.k��b��MԊ.l��d���u]���m
��3�����8'	�Z�s^eh�����<9�hW�!j�S�w+GǪm����o���%��#*��x�������i�]Sr�ytfh<Y]�4��i?O�R�/h�7�$]��ث�f��\W�=?.-3Z�X��e�.5���'��8�o���7�zj�3_��g�E-S�a:k;�o�3]�Q�j�����������&�y�b�kJ�:%�h�R>��9�!j�+���� r�)��(�8}�S�۸np	�}-�hI� RT�L� ���<���fH��n����``դ�+�r��E1l<��
B���LrB����G��X�c�[Hd��<6�� �/o�M�R7.u�����qt�i��ǰs�3��\��h�#��ʇ�]�k��|~;�L��y`�0'�D#�L��J�""*��#r��6)�^!k
�����`O�Y�0�m�[����Z	>'�g���])7)I��\��6��*��8jO�SjB�6�ȨUW�m���Z�=��6-g��X4OK��K!i��@mx��=��:@����"r��CE��"��i23n��FƬH�S�U�Ca���m���Nc9R�i��,2�Rk�4>�y&���H��^�OR��cl;���*Z
��Y���\��&7�X�s�@��w���Yw�~ W�Wǵ:���E�B2�s������m��#��jz�}���rV)�|+I�յ�y� ���7&06�5}O�U��/�a�+�~�b�m_ �f'(��޵_i�OR\n�@`K��p����>�ACf�d�<�j�wgC�_���B�)��6�ͯ�ne N��_�FA�sRG�{ô��� >Qį����U��:s�zOp����551y����8́�����G�������.�k�5o&���(�Ɖ&dd���F+�q�=�Y�"L_�G"2,�T�嚡�'��ܵ���)p�`��p*o�C�EB|s>>���!}t�挿����qZ �\���mK�W�G)��|s�Ɨ����s��k��s_���d��#�B7�1�
lBR�EH�u
�|���ǝ�Qe���%�Ñ�u���J��%͸�4��O������~�"�͢����#0�OHK�ǃā�8�ǀ^�B!}S��F����Ȭ݈��j�ykG{�A�P㞣x
�o�USu�Q�[��ټ��!�
e�T7f�<bM�īvk��ZȦ׀�Ɇ�j�$2��N��&��ϛTCۻ��o�&�k/���u6���[,���6!�2BjK���x@�轅+�,;�2ʻ�n���úL��ب���:O�Yq���5��+]}�0�b>M�[��V5*VRɄ/���ARՈ��o	��<�v:|���`ϰ^Z�ƹ�I�C���ܝ�:�TY�$t�Qr)��}�jM��CTS�k���v�1�諸�[�b��nv�;VQ�resK]�\n�dG����'p�b�V�L����k��m��_���[n]4Wh�gGi8�"RW�h�n�ʷ�!���Ş�$�3�n�w�-��"'��4��o�	�YWB�H��#�3h�D��_�mA.���9̳%��q�Cb���{����Xrz<B��f!��E��[+tX�z�(P�rZ�`��z��*68���E�m�NY&����n��<a}�(�j��Od]KA�vN�>�e���+]�
s���'*vP+�>	�-�6
�[d[��Yj��oh�*�кT�:z;�38߲� ���ƒ�8k�vW�7g��[�7B%�c-���M�M,�*�q�L��.$��$�w�?���=a�Q���5)�$�
ۋҰڞ�}��s���lU���^Dg)Ќt�q���[��������)�&�>��K���6��FrY�`{|QU����=�20
 �*6>��$�O0=�U�Mbّ��L1%ios�<p��l���ot6�m���oI��V3b�xҠ���W��Ob����A未c�[��zq��8$�����:Ӭ��\�o��Bܠ�z'|���I��zẶ��[��5D�k��+��
�J�'W4�����yߚjYE�l�%6΂��{#��+�_#�{�?�9���X ��}�U���n>g��͕�x��C���Z�~�9��ۮ������DX;h7��wH���~�@@��d:t���@��%�P���i�Z�HLLY<su����u	�⮦1���}qa<o�x�9�e�?n_�|�RQ�
�gT�>�g9z����j)@m�T�V�]�l/&�~�r.�*�A�{#w�dլ|�:D��+��T\}!��³���#j��� `��:�$k�ڎ��>0$�<@s�[�9}q
�K5M��$�y���"�'�k�Z���E��M��|c��:��+w�e�@�a|�;l���V擖�:]X�b>TVw/�2{��)��5ta��U����.�k�3��w<���ٓ�ҜD�1$��σVk���k����-�{������#h��6�ŝ��LqVuSU�`kN{�嚰_�M�.��}�@}��ul���Li�S��g���5]�+�-��`YTu��x2.��e�̐hY2�~�=�j(���UU-�7�&|����Z�"[�%���dt��W%Me$��ɒg>|��U}Q���h��{�=�4G_��x%�1�w�^��R�Wy�[�̩h�h��B�[�B�U�r���Dҝ͞��V��-0"(vߍ��X|�����*���*�l�DS���d��Ed�L�[�~G;�f�Z-�ж�%�Ȁ�|�>�~�@��Lh彈��6z��Ͻ&	e��J� LOot�:x��Zg�Ϟ#��(#���.�Y�L[� kC�ի�.������|�륟���a5m^�:V��Q�T�c. ���X�	�BϹȂ�fe����99
/���YZ�h�c���Щ��A�ac�fӢ���ojA�_�b͏��������ߞ_ ��z��I���:/ r}�,��C "l!w,d�{q|��Ǟ�������sVα�m>�Z�D[�N�85�
�m<Q����)w�������C^EnQ�S�w2��X�D+��J��0�Ub� ���Ė�S��r!-f�X:m|×/��R9���7ƽ�4u���]�&�/i���Ѵ�>�`�rX��,�,����q�ߏ�����jk�4�������$S�t�Œ�����o@$�q-��L�`6�L��Aig���gc�ᶂ��p9f���:�����F�i��}|�.��E��+�ɴ��[}�!�377!V�W��v� ����(���fūj1��i!S��w�x�=x<)���!5����~U���)Db�[f�:S�i�4�+Ͱep[5MS-[f;�/-�4�S�mX�g���e�8��E�nIV�߶��<�IR�D�+��s�
H��ZU0���Q�㙹��%*�D�r����-���G���w�����׊h����a��-R�U ^z/�_-�]y�e�8;�M���+_S7B�4�
���Ro�y�m�+?	����\�ݫD*�_��&���NI)�;t��&yñ][+�"թ�!y��˙�z�Ֆ$YC���0�e��[|ح1ʽ�y��OM�zܭ��|q����VΦ{U�Ѻ�z��֘��XS��y�"|��;�i�x c&3�ڷ��k �Oi��[ׯ�6�m3=?�U4�ݴu��x��#1�x()=ׅ7��'��B� ���Y��idr`�X�oH����5�2��=K�hla�h�l��MY�^��$�N������Y����*�� �R+����-;��ؕ����kƱ��[9���{o�XV(����P0O~����NV c����r��S�E��"�6���@����w��Z݁�#"]�b���)�(RazG-�UC��gp]�9%�dw�r^)6tt��pҷ� �7��uX��g)k�5��q�x��G�
���6����^K���x��0�c�sQ�&�H����a'�7{R;���l?��X/����
Q�^*ik�����8a^s<e�" ��N��-�9�t��u��!P-�����'�CAէ�W&�r�+��f��]�߇%&a�k>���>֯�����JW���U��Io�� ��^�������޺�ni�o��t�_T�u7-����C�$�H�l�7w`�k����Q0 S�[�f��~��I�\��Q��'�6���L[͕6eE���*�#��	Q���3�R?ې�Q��"4[�3����ʘ�Z���eM"��\����.�4�\E��s;Q�i~�%X��X��@�G��?�9e#�~ �N�DV����X��&;a���L�)��6� b���w�9�����:��>z��w��7���C�5�&_@�	iI۪�|���F=��lG�2R޾�wyJˑ�{{�̱O�_U�S$z�3�O�qЫ���{���E*#1�x���P$G����GƄ� 5�M�'�<��|����9�SLf)�Dn.@K�׬�D7o�Љ_��6`6�^w Չ�� �2�+� �D4��(�^�m������@�᯼E�'��C�șq��d�Ze����D��]�.�+����:�t��ʐ�5�>�M�w;+'v�pX�<9O�������r-nst�o�Ho�P�����ֿ�<�H�LW��Z�eN2��4���O����ؕ?�{?�id���;�9t5|�0��M����'!�O~���ᰣ�	����E�>����)c
KV�z=��v�cv4Qm�]�%l{_�/���J�z�DԲ%�������T:�G�� ǂ��-�k�=p
�h*_.cr)���b���n��B�����M����ŝ�@7wT�
�*�u}��ļ�>�Hnd�m-��t�S˔`��mX���?'[ǭA�64�3Q�E��u8Έ~t5xխk-h�3��	���f>�9�r��i���t�m�W��x(��;N��&���C�ig�L�K�yeMHJ�7+<��T�I�������U���o�,���[U���@l{�zh_+��~��y\T{�Z|
AA��S$:w��	!�YUa�|�u��C�^U�Ms�����Z�Pqc9c��V�/�a)�
�~�F<|'�6%�jk�)��@��v��x����6�E��EK��+�rx��u|PH�	Qq򉶵�{�T����O�ԽOڵ\pL�Ś�%��S}��pKqE����'	U��8VP�s0��\:�T��5�(<��'�K�Ι���5.�������"��U\��H��"N>X2��f�p
[�e9� OF��4�(ܴ��ͼ���)��t2a���(��R]��*�
�2y B�0�,�
�I/�{_/��bsw�y���??~�U[a%�3`+��կ�DU��ǧ����>��1Q\��
�l�����<#u桅'�G��3�������@��:�[��Q���a��N��м}�Ĺ�*���&W,���.�8Җ|�t����%U�Bk;ij��gpM�̅�v!)�\o�g*���bm#I����a������P�!;�X��Qvn3OU�L<;���tENe�[�@fv�p �%��s=yd��ѥ�~��]�]ҹ��N��k<YZ��Tl��c1���1e���\@YL�Pop�R �[� *�솆C�XS"��R�O'� +?/��$���U����N�z詡����-�Ƀ�-������y�z ��`o w�ne����~s�>���2��Д����R��+K�M��]��tų�Ӽ�%(ķ,a���5)n>5ޣˡM���	>��4���;��N���R���2��R��&�b`�\� r,s�����e�$��D2�ɑ���jUG���{i���XOmu��[���T܋�3V��%_ҝJ^�:K�2�����ƻٳ�P;\�~ϔG�)�Н �|���R�����m��r��[W꼟�Fi���ɯ�6�|�^�^ee�Ʈ�trL~'�݀���ee؉)e%�X�����u{}N��:�!��l�4��n�c���b�܉m�?��CN֖̂Qq�?��@�^>�f�&�ȃ�[o��M�B��M�"xj�O���l�=�������ǣո��x
�iǩ8��|��s���׶8iw��L|_u\�����c�"��il�1�>?�*5O6O�@�����H%r��M|P�6n;o���-8�BK%_	I=~܋�ۂ@HSVAeU�LV�򛊷�y��t���=ҫ� ;_p^y�T)|Y-ϻ����\4!>��z�B.�|��҅�<3{z��Psv��Y[�Ϗ� �L�6b'b��:ې�싮�,����=���7�$��,'�1w$ׅ����C��6
@�9�J���F%Bt]u�*�+���4�#@��߿t��*0�iZ��!a��I�VjOc�т�qq�K|9��'�Q.4Wڐp�~���D��9�I�)�y��N�
Iic��  �A!��n I�p�`�p��[q��9���6�HV��`�WF|	AVMw��/��H� �QTJ@�˶+�Zt��5�f׾�y����8	;`��H|���a�zk����'ʧ처�S�v �Z?fIﭠ�1��k� �X!��e����^c(D����ߊ�y�E�A������F���)%*J�H~DR����K�I�,ѢU��A��;a���j�]��-� �0��6�%���YEb=xk��5�Bt�h�$��R C9���N�����ҧ���&Egc�)��7�:�(uaU/(=�H)<�ꂊl�\^����L�D��JS�G*!��Թ����6�U��O63T�����R�W��NIt�z�sڱk�`0�-3	 N�1y�S����3�"�꽡Bg�B><4�d{�$	+b�Xez���zԞ$@�	K��2���9�:\d^_�݃"�u,Օ��n�UV��Rd9��s`6w9[�� g�?l���R��c� �h���cB�b�������^��*�q��9N���*vLZ�������e"	�أ��Kޱ��$Ia*g%��.��9���mXj���/�1�j��@p��d�f񑈂�dʗ�X�S:�l�.f�w�e�u2�߾�dr�}�<(��1���k�}��sJ�Xm�̩J�.��`�GGr�ԉ��@����]3��������^LG�e��O�2G�n�"�� �7��aʬ�ry��7�ۼ��}b!�����Ĕ��e7�WW�Uq{�H9)�ޤ����O�b�G�x�T-�gK�'Bh%j�2��>i�����ȴ�cJ�/De0[3���c���p��'����ȳ�N��&���%H�o���3s�u4)9}|�=�*�,qV����߲{�+�[���_�L��XGY����d�m�nz�ƽ��%U��2�Yʹ���c%$��Y"������C�=�`���Hy��*�C���@���s*R��CDÉ���Д4��� ��9|�)��׿'I�.���/�g�}1���������,����j������ ������~������I����w^b�����^����?#���S�Bw`�������86�L�C���0����^���%���|q���9=d�4�+�ލ�l��!��]�dϮ�Y��5�:���-����%@@f[�J��'����@`�Z4o�k8gԋO��>�F��$_Uy��D����L���o�soߤ)Qˍ�1k�T*���Qd~����'��<����c&%>�:�=*�k�-�2[V�z�>�f^���4}'Xh%�3���Ĺg�X��~�~0J��d���po޶�ŉF&)�CZ�&�'H��JP}�<��f�*'ihV�����w���D�2����}����C�AA���Z��U���{�3��߭2f_�N����7P#:\�`�[�Z�ïa�8�}�+� ڟ�*��Y?���pMv_)��2�Gz5Ri6��t���:v1^�^D��lk��Z��$Iվ�WJ�܌�v^K��%li����~\�x㓈�v���(�!�8���w;�E�&�T�������
����Z�+���^��s�c�z�A�Zk���[UM{�����{�a~U}	�g�0|���RH��^��� A�|$�x�*�Aά�����"vW�n}#��r$Q����@v�&�4�[{���Y�غL����M`���Q$�|xq�xR���#l��#J6nf���̪�J����7�V��g{"���@��}�-|*�&	��|�y��
8����s6�����e2%��
����X��C��}�U{�T��
khO��
1���C����9�p��
^����:ع4O(�mJ�A��g���!���{���+�M3��fP�w�&�OG?�|E{Y(B5\m�l[��'��l����Zo�ը��
�����aJâ��K�M&5�-,��H���md���<�j||>"�>_�T�r����~Iq����[�}��Hy�(TM&�`��i��rGn�t����,/2R��!c�V���{��{��۲N�ǈ�@6p��&���z�F߷ �=���!i������S�c�2!��C�%Ȃ��;z�b��c@6X�=�j�ve8����4i�2sF�೩����(��"C�À����a���`�����pn�NV�H�p��C�FDD�33Ծ���h��AO��+��e�&���ѓ�)��|ȉ�B�rOxC?��D�����9@��햎ײ6��c'��y(9�a�v�hV�黎�X4d�j�;�����+�v�T�����8�#Q��d<���õ���-��C��&���cD\D��O2�����+�`��J�VP@�́��Z��!��6�juu���>-GkX.&ᙑ��0�hw�¼TRp��W �W���u{
,>MaB$i�R;2rr�Za岦HUϖ� 6r���-Y�tH�;+�e!�������wH�@��P��|V#kV�ݬrO&1���8�ٺ�Iص��$���?���o�lg�I��D>d"���L����hM�b�(˚{
���ha�\Z4\{�*4�@n����k��i�o.���8	[�t<��q�(C�6"��T[$��$�d�~6<��RL�(��Ob��)��\ �J�]CB9��e���n��,��4Rqp�b����gٿ���T�=C���i��{�l	�Qv?��Ņ�W��r_�C5��;�K��V4���0�ј�[�﷏�=�[�٪�����ǻ�Ʋ�~=y�]�9-]ћ��f��f�i�̺!�	�b�E�����(w햾�w�Oy�_iٵjﾹ;)���}|��8jt�Qvɦ-� �����OD�����gt�m���'�䞻����!'ݭ��ok���W��Z�N��}k�L|k6' ϻ��~�����銿P?v<j�J����?k��vtH���J��x��*D���E��.r_+^�����D���+���$��[f�;SvW����J����t���5�����U.j�	' �nw"6�@�����0�W���,�+>
2��씎E������	���QI���0��>�ik�N,��U#���p��r�p�ũ�V�}����o�������� 'q����,����6�kLW'rx��e�>'Q�u��j�����S֛��������a �7��
�t�Y#>��#�5}Oj!غ����ݨ*�*%8�U@Yp�έ�njg�ԝW���a�q1QG{/�-0'D��������/�������L�/�V7=^�{:��R����v�cJ�h|���\G�,���SSo��*��Y���d}���iX����wT��&�0��M����� ��U���jq�6eA�����|�H���B����� ������!<.���@\�j-$��%�^�9�M᫴/T ���ơ��;�}Z�Eҋ�V�9Mm��և��ߤ������TdDT����i�0��9�(�U���YH\p�f�ïL�<��,�����NU�1�bg�>�!�7�W��8~[��!҅���<o����}O��А�]�������i'����:=2��m�^�=�E���4;��z=W����t}���B��#��%Mb+��k|ޡ���	��@�PuZ�l�ע+Wv�y\�eWf0���:u�i��b*p�}={|2$ry�2_�ʊ��7���5��1��&�ۯ�����uK;���|5�=y��4�5x�B��]T��y�(B~TOA8��6���$N�p�ˬj@ZyvHh��jrM(b���i�>����(���-kr�TŖ�����u��Ğ��*��z}��k�6� ]	K�~Ř��p������=�.O(��~�[��Z�����\Ӣ/́��/�ii��yը����O��%�[A?�H�>��䞿N�%�8&�IW��ү~m�Sǁ/���ܤz��qG�Y�,Y�n��ք�zD�!�����e>+P��vʫ�~�=������T_�e�>��|�wJ�"��z`�T�+�;Ojգk<ޱ&�]o�Ђ싮&Z�2Y����D���)j6��p,*��֏�|(�@���E�?��M_�[ �*\����缋��zE
N6���s)1��6J�6�������rDG,���x��Y�Jջ��iЂ��B�|n�E����2��4,�iN�Ep�݌ii���T1҅T`���]���W *����oUS����ʆ`��<X����3 Xx�b�@�!�7�\����!�!�4��3T��hF�Չ�bx��M�}���i�K��+��
���<i⦛I6NCwz��m�v�F#�R�r��5����y}ҥ���7��N`�*��½���s�O���3Z{7+-��8��ֆ�V��Y��7<�i^��;�4eP�a�hi2�2���ᕧ���~J���<O��%�Q����%M`�ƣ'��9c��)�.Þ��Z�*NÞӒ���g�6D��z殍�:;b3�ӊ������n�e�秫����\N�`�9��������<v7���Ƈ�$~o�y���ޢ�:�0g�y�%0�w�Ea��9�^伛��a,�M���;���P�T�)�3l�%���q�>�S�߽ݱ�������]��'�?�)�g26�7���`���D<+.��ۏ�?��L����)���DN3�����79��<�ʜ��%�pjʤuֵ����	=�n}����M�S>�O5'���k�1v�[Ke�vkS�.�����ݺ�)(,l�1�����h�5',q\�MgX!U@�Ĭ���5(��{m���W����9uSS�A��������k�r	X���A>�<+�U@��tБ��=���̵Y�WB[͛�$<K����EL?ui]̺Ӝr-f����w|��*��>W'V5?>%��c�F����LR�u��4ۍTa;Af���G���*��n:�R¹/�|���8������[`u��$�-���,�������ӞZ�0_���� �RH����sԲ<�<���GaR@��y��+	�Wn�?�ʜ����%h�!��(�l.O~��Z��=�*�DI�]:�S�G�`���Nd��������kVb�&gm� ����'Y=�hO{Ƽ��}���N�X���
�����[�\�����?t}�V�M�0C���o�\'�>�P�?��d�Qʨ����1�y�[�)G���j�n��8jf���z&�Q�ityr#�Ϯ;@��IׇV���\�|ˉ
�|!�$"BWɱ.׆(Y�Y;+/�x������^���z2�U9�V;��m͸ں���Z��+�Y��8��>��-T\^��T��Џ�䝒cq��R��m�\�/�5a[]��m,lEJ��Y�Э�4�9�ǲ���c(����_Y��[�d����B�}v{�x�f��?���Q�������r��FW����䙩��r��`8�礭��kK
=��t'x���-�p���Q'</�+))Io��N���O�b��A/]����j'l>�^s����Jٔ�hy�ONӽ�g����ya�f��A�C����'<�.�� �Eq茈���O�/ӎ���%i���63�����e�c�~}o�>ͩ__���i&F<���W��i�;��ӽ��J�u}�6��Ox�衉L�n}���>Gu��(g�ޝ��[�O�D73�jڇ�����?��L9l`N�~���@�J���Ldtt�#�^)��� ���`ϵ��G����՘A�{~�]i����z{��3ix�U<1ES#{Ү��Օz�E�i$G�׉j��5��ΏlG��� ���QZ���B�]�Q}�~��Դ]4bc��X�s�����JK)X�y�ݑ4ϬfEۈh���Z� k�iJ0��6+J�~��I9�3�1����)������E��(�ds!F���pv�쌘5���^���y˹��4V@��f�b��#\�~mmm�di.��$E��/��;i~dH�'���kЍ�&��K`0��Ȅ��$v`T9������iJ�w���]nz��?�9�iv}�c_D#�#��� �:�����N�>���L��c8���Xdd�ܑe>�<k���MrV������P�;�݇�9z��`�Vs�P*�ƳcQ��=;;޾�5�y�.�;9bؔs�ڵkĦ)^>>#E£iJ���-����BQ)�T��Shcy����]�X�&L8��M����P�@�k�#��������QUMmֳ�d컿�q�<1������5S_jSߍ�_���@��5���1��!�6+�MS^�!�V����f�L$f�/uf��)�n�a��]�_`5ݹ��3�4P���:&s��۞$�#�7;e��t�5��\���gmy5�5k��$Tf"�C�'ݺ/�w�^\�|j����K��5-�*R�@�7ä#n,J�����p�NJ��� (l �!�TU	w�^7�t�KH`��l�%9��_?;#�+ ?6��N��g�Nv����u4����e�d ����uj#t�jCG�l
]hQ�A��陘�\io>0�244�Ƹ�O����t��ׇ�\�Ħ53X���1���dB��8c�O3��,�ç M���K�����0B@�!��R�GA��۪|Ǧ�� ��T��$�۲�w�G&� @Q�m�!D��N�.�y�Λv:���`0M۵��ݑ������@+��6�e�7f�SRRz�R�(�Gp���L䔖���!��e���?��F������FH<�i�|�y��n�%�,/�.�y��1C�-kdj�/x�HR�ABH+q2�;��}]A�f��<�:_���jW�/s 	hӯ�B߾���<ӛ,�ׇ?و>�ݞ@�_E�n���^�1����E4탊t
�O9�`�m�h4xm0n��]q�{�`聑��z穆`��mf8X��w����!t�;ݦk�w5�1?7�K��������"�[�SJuL���#�c4f��C���0W@� u��y�ޞ��Q~%�X9�!�~��+°�gv�k8T��y��<�"�i��xe��z����i~��>)""bfq�������ג$���`������?��������Z�ciP�a�-jj��s����Hg�b�e�8��4�d�FW��ו��Wk
��.N֗���</�{7���B��<�#[��wt���r�4�Hp�~oy��Yb��)\s Ja����a�!��K'�!�F!��ԿkN5��5��f9�~���fW�A�B����;�q��4��#���5�%��y�ɺ���ݼۍ������,.l��m����Gwc.ǜ�>J|� ����̧O�0U=����NN �0ź��Ͱ�wu��n��������i�����\j�+�9?���ܻ��.o�P�>|k��33\�~��S#kQ#���ܝ����@��XǫS��aL�!��g�ai��U4B�	��e�c>l�1|I�N�X����7�1}!�ߩ��s�{�������xえ��ʭ@w��&��-H�w����[I���΁?����.��~���j~9�k�_�\/�:�Fs Q�#{l���3���.����us��=dJ���J��á��GVN�WjD����"��O�?ן
=�ރ�0�a(P
Ŭ�f4�72u��F��4�,s6oJ�(�j�� G\�%աV$5�cI�'�;�� �#��A��i1�[_Hc��G�N�`6�N�W�68���!�� [�q[��Ą[� U0���s�Y﮻3��̑�3^ 7X8�:|bpp0P��� `�����fA̛f��/.��{_G�����:��*ۀRpv������	O/��A"1t�]��JO�ز]��׵�k#�#]�ă��*�@f��� �6�0��U�u�FĕK���~7����y��0`��r�գ�-��uu�&N���l�T���B����>bȄ;����*�s7���s�K-�#�K}H���V3E�B�w�q2�1��o�\��^�4:qFu�R�̐V��iAd2���%�.|p���S��[�}����AT��Lp�]�#!��5*��pM��Xp����#�rt�$���Z5~��>�	w�e���C�B>�(y�i���|�ږ�C��ߵ?y��[�D�`�(5�"��i;ފ��̯�@j6��i��V
��_鵌�Z�o�d�{W�<~���E�#h�l��$�\jTS�8ɥ���Lpв/����s�QGBنPQ�EA��7!�����k�ZD�+B-�f�c`޸��t�"o�T����'T#8>�F�
����W8S�����([U�F 8J������k<�o'�n`�����3��kߍV4B�Y鎬��ݻ�o��A��7��N�T-�F6���g��PB.;�*��J9�+r�/��yF����X��8���zn�T���G<�QA�a���ܩ�a��^��,��
v��/��sFiՇH���s��>�q�'+l�J|�1�d������B�xvv�DyVPa�R�e�0���6m���M]<uȱ4J�c���X���ɽ�eUs�dnGAv����p�� �R����9E��z����fEw�W�@��.�1� !6I��b!�HH�R����5.h��K�0;���1�wO�"À0����N�s&�1��5�F]�Y��Ai,�Xƨ���2�ʉZd�&F;{^���}iuv�{s�3Fri�?r0rf��$H[�0ȌX�D+O�;�B{��#�6[3�x����V:�@�Vz� ��:��X0�r��2��'��
˄*{Њf�x��	O�gb�N���O�t���7^~f��B�|���l��o����D�*�R����l��/�gEWk$��r� t�OL��˭�9����i�w\jN�\ҫPS�4�*��6y�`��CM?ɛi,B%$� ��j���oȥf�@���x3���#�;�Ԝ0�A-�.A'#f�VWW�b+���m& pU)�rt���f�I5�yp�<@r����� P�O[m�un�D��v����$�Ù����v�����*�I���f- H��v�Gieq�(�xfZ�8��ˠE��w?�a��0�������/�������C������xV���X���R)oeH�D���>�7�D�ĿI �f�������B�P�_��kte����
(��M ˰���#<ѵO���Ȉ)
~ix��7�]�]��a=�p��������ֶ8�wx��r���QGy���/S��	eh���TR�_���,��@��@�u��31a��~Y}���'p�w�^�����`C3ޕ�~gL�swt�%5�H3gۦ"��2����܎G��.�|��?�.��`�/�A,I[�z�4��eʯ1�+�s����8WY�Ɵ���IE������	�i��+�R��p�6y���N�Ǌ97�Šo9����!<I4bsrA��+h]k:
��5K��J�L�S����:�y|�PF���O?�mɓ�X����_�'���yY�/�mG*� ���$�d�T�p��d4��?(�%�nx,��)�+)� �o�G��d�F�E����;��[�*#���s�L�~.�%���lu}eBr3�>�t�n�h�z�pt��Ȧb�vK8N�`�2<��F��3���eƺK�d�te����6?�س����{�G�7��e i��x�r��椄��Q��$(��P�}>IS���%�'����� 	A��Ί'R�q��3G�`϶5N�bHT"�	��PWJ��A�/�RM��G����EN������
ZX�X�^�i�_ڒ��`�s�\U� ��Dg����B���3�&��&�0�+c�v��\BQ�v�`|���Y3�_�4�ܴ:�s��]��/��iǀ���|^瀚���)p3�!����_�T����_��_2Pל��z�+��?A�_�����s���1j@��?~�e}!j�B�GG��$��?Ww�O���i����E:������6}�:�ԔRO�޺����ڰY$Q�8W͘)���J;s��٢��SCr��z�h*G��@��������V����{q�j�.,��ڤ��࠺G*�j���[�>��ͭ,�V��&#��C����)�;Cھ�OteJ[���D�C�#�#I�LD~����������w���Sh���ƛ���d]kh��
�׈���F�֫�5:?���&�4���&�E�ѕ���W�]1g�hҢ���}�-�(3�#�kلL��`H�U�ss$��yh6�j��[J�~ֵ	9V�[���f�O�'�O��K���eX��Z.��ҒJn�_ɤ��aF�8C��M��@��4� �n���7��}]�]����$4S;h����Eú��]�5��_JF+�90��r�:r�͚:���s�Ṕ�T���
�l�j��}v2�ݻK����\3 9"4�u�ɝ�\:E~s$Ƨ�}P�>��K]�������2�,�+̻�a�S�ow�rG$O[^q��_0�t�|��k��ނ���'1w�'�row��H:�f{M�U:W�ƅ�"'w�;H�֜���7vp�mR�S%bg�y���J�;�rJ�y�'��6&�]�:�{�ѧi��{D��azU�Z �yb�ۃ�:����'C�[�8~ћv�Unx�Nϣ۠c��_w��s�=/��r
7���gs.����PMfQ��#��)�FP�)�;
�(D��4�HE�A:""-(ꠔP(]�H'�z �$�������]�w_����Y�q��s�>���v���\lUu��n����p�e��^�i�kWJn�b��4-��/z:����{�y���hK���q&�j��|�{G����e@5���mR���ni�q"n?~pb+��cV
4��� ���58�w�����Tg�ON�-@nn�Ȕpt�hB2�>Ι��^�m�c:���f��n�x kr��6��M��{��n.���]��	�^��;����w4������(����?�D��O�?�D��O����Q,w�}��t��������G*�a�j��8��ess3������.S>�.�6��E �M5;ח�fw��<G}����
,�KD�r�䕏(V�M]wi:��Qz˽�w�ƈ[��N�}�<��HS��ȃ$�Ra����
@:e�I.����x���pj��E.����͔p�4(ES,w�5>5S���_��Q��թ.��:�q�d����*�]�O��_���(��.��k��B=�!���|U��5B(��t�X���n9,�U�P�0��f�O���Fn��g�WW%����{��}n����W¹��~��O�
K�����=>����V^<�${�n�۷o��~5�T�P��RI-��um���dP��k��9c�4qM�;y��^H�/^��@��gyp��2��Í�Ύ��ן����.���<��}a��dT�_�)/]�F�r��)D��oom�ඬBH��<QUES ��HҾ���k �=��q����;Z��j�[m�;F�����	e�=��%-�g��V@yG��*�_�П"���'��FH	���\�t�α�[�Ł�2���<K���w���~���'kO�	��Úl�p������Y{T��2tJ���H������\$!g�7v���1�����#�#45��^��@�!�j�5ߏ�Z��A��0z�֤�hȔ`��LW����`���!Ͽ�0O��No0�65���]L��X�ʽ�&?���ի��mi�j�,� ޣ���D�%ni�H�!��r�cD�`4)A�љ�<��n�����3�a7l��(pUY��u�8��"qi9��bBi;m���IF֖�J�?�)�:�G�G�r ��sjϏ.�˯΅���\��2A�i� �咱��&�=����DG���1��_�V�yɸh�;�<D�x��y����It�����0�#��xM,_D�*t)�f�K7op}�%�q���a����m:6|
��1
����
�?z��Z���!G��l�y��,��b+><q���@\}D /}��~4���1:\ӟ�}��h��?rZ)��u��4g�����u)Z_M�zN��; �E~>-qͪ0�>u^X�M�M���Z�l�%&�ż^[��lME�Ѫ��PNvRMJ#�F*[ :#'Kp�?��yq���l��g���$4�1�fu̪��*������N����T�ՠ�'�k���u2�د����[#����jl6��p��+���u�ܕ�A��Q��oȺ���E��L�����?o��JQ�BQ�ZG�
�[�UK�]S��#2���H�����x<�.�8�5d]��{���
�zN
�覻o�����\*0pjE�}�@v��}c R?W��w-�p��v��8pbǥ�};�����������_��y�����/�<k��!��`-���Y�l��dԗT�������{�\�דN׾���6Ɂ����YJ�vk?>HG��sg �0yQn��k�4F$�5Į�b�Gx��U u$H�>�]�k��`�<�c�b/o�D]�^�����7f���������1?(|�:�N2����1��wא��{'جn4��>R�:��#�<f���L*|ϒ5�x@V��Q�k/%4�
�
�uF���'�$��n��A缢zE$T���������f�\C|���P�Θ��#��RY��819���I�<���o��C�XǼAZh��+���Lq��M#,�X�8N� �4p&N}}������-�m��c��+X{A�������>�=�F-����kLh3��X!�����m{�p�{jf���c�����y�BE�f�#E\L�L����+K-Ǝ,< {n�0�Cz;��\y�L����M��2�����:����Ck��}N����������TmJ��h����u�W6���߻܈���1��E{qa��X�z�*35�	 � ��C���}��E�jʜ7�z�LhC"���kGN?�x�&'��+�C��ܷq�/`���
�������y�J�W�@��EB�_�#�&S�����?����
�1F����ӉK����"�&8�S�[uB�b
�T�2C]+�I��ty����,��@�x,@̺��7.5v�/��>* �/%.�>�V�^w�J�#�x)�����S%[|�/��;�o~� ?.�,��&>|�l3��t���Y��������w*�=E���� #��sI�ƽ��FD)9�k�B:���IS�ݻB�]C�W6��;�_����x��r��y+�I�0���ɩ���o���|Ȑ�F�]��
գp,��Yn�u2r�ע�à����K����z��R�,�tEҾ)����{��؍���6�X� �G�G1um%$L��I�j����e�0�X[Kv~�>��w:p�z���ar���p=�L2:��ݶ�풏X�d�q���]�#*\.�#�ݪ�+_+�2�30�r�j�������<G.�~���
oBյ�]+Ei�׶2:�z�!y�P�����k��]���t�A�TI�����\)o�{@\�F~����2��_�k�^%��(v�_�n|�-O���H�Mhs�z��Iv��}q�k ���mÞ�	�]���@�؛����,�w�Q�qKaa��X*�R��<:�J�S�`�W�iK���B	�C9�,��������D��'� h�o�TI!/X���M���5z�ڷ�/�Y�qĕ��\�C^�����������ג��$S�ʹ3ل#V��r�O�ؖ�p�w�f�t��}W��S�\�+�7\�N5���f�]�p�"[T�D��ۏ�_��uvv�f������_�.���{�a���W����>�5�"�KZ~���J��\S����^�zspГtGW�� 7;�#xq��7XM� �i��D�F��u+�{��|����[����{��Pp��J�����Z�?��=���4)���a�hz��GD	?ݺP��	-�VO/d*wM@M����
<fBU����eW�IYɺC�1u��S��������5���H�X2y�5V�@޾�+�. l�5�aeƄ[n5aM4�Ɠo���S�q����|�ˉ
�(Ș�����K�Ԉ��� ���/�	�v�+bkF�Q��#?*�Ԟ��vШ�~��|�����xA��R�~�T�^/oQ�0e�����Ƹ��������\�91��A�No��?�bR?]Į��)&&�%���e�U��ѽ��3�2���$�}1�DQ���[��6Å3!	9�o�6�?x�T��G��e`�Y�-+,999_�\G�͕"��.���܁\ȷ�X���\���Jy������Gp��L_;��y88�䎳 n�����*K[��+/S�_���3n�)�K��H�[���?r���u�#���<V�k��s���2�(����B�Vl4U��dqa�3�
f��ʄ�X�$;�',�����yxr�RdY�54�D�>����ׄ����O4ϑ�m�G��"��ɗ���P��}C�Q��sؔ¹
l����A��'ob�pw�>A�q�7��{�8
�hi���8A���=�d���~���$�Y6̄Y���e�^0g��}�-�˸R�ޑ��m	���8g�4�ח�ó�h�3������>7��>�o�9CS��5T�j繐G�B��\�3ԝ�����`�}M�e#�.�vK���*�]�������u8>F������e]ԿC��u�O�L4�.��H�*�nޠE{�F�uӏ�E2W�
/�+X�	R]��K�)�B���W����u�?����7�ӝqoI<��v{�e+�'�x�VU��{�h����=��:�eQWV��R�bg��vѾ�Uh'�n-\�Q�/m�
���&]f*P����8.(�����d��:3��	!��â�;����7X��>r�~Tu�=gb�Z-�>_�["H�n/�a���K�{<`��,:o�;��ci�V`�,�h*�i�XU�g���^�T�bsr(V�D�����U�_p���K��ÂABe����f�:���q�?�V@��RQ�L`na�ix@�Z��ܞ�����g���.Kp����Eb����]+kd�vz�����,�>�;�I����p,��Ç���]k%��$Q}}}���:�5��9�E�������r���Q�t-{䉵d��x0���>x�<K��3v�����0��m�� �����y��䃔��&뢗�'�����i~F9!�UH	4�Cu�1�� g�濖�L��؁��Xy�r�\a�V�Llnn���t��S�N�-l���'hӷ
�� �;���/����!����_�	N
F�zf�����dt�cFA5���^�UfA�Zu�9)i�lA�d���WTo�	z$ ��F��P���n��|�����B`�N����G�Xg�dLyy"�>�wB��߇��\PX�)z���2kH�E��Ӧ�;��#�:���t}�6����5��Kd�����}��X�L`��.��~��P��&=NPY�N�n�,��/�|���S/��g�/ʮ�vyX���]{b�滆��3T�d=<�$�Xr?��CF����gryX�ԙ��i�����*��0��e��\;"�ps;j�jr}Hr��%�6����x�P@����i��=�]��pK[��[J2�R> 0�7�BKl�/��/
�K_��	��t��C�LNNc�c���q��=Q�󆼞��^0��Oy��Vg������ e�^,N�����d����.+j/h�Nq�6�U�&���Z�fbr���`�>�&��lsFe9�X����[����5)����Q#�|h̢+� z=i���3.Z�<11QǔȨ?�4�� me�p�IS��
S���Y ��".`��ԙ��\��ҏv��_l\\���n<;P�Ԕ-�Mt٠S��(�������շ���`N͆�_������q#F%4?�:UFU������rz�]���~��\�[M�n�g���>`�S[[[��;�����Ph�67w��7�39�-���
���CX�3��yh�R��j��H�tvvf�'��X4�<`Jj����H�?�+F����^;pr�����e�I�+<]+ �	�zzzZh�t�B]���@�%SiQY`ٲN�\��R&'ݔ?h����:]�V� mu٢�f�&sh)�fK{�=<��P��-ҐM���N�@�~s�5����qxju�K��h��lv�2L�Y�ͨC���{�3��
9��S ��(�7���_�+oI%�b**-�X��(ⶵ٩I�#\e��d��u�(]PQQ���KNO�+@00�Ծd��|�UN��DGGG��V��.�����)���n�,Z��e�nL|�tG�e��fuH�����8���>`)\�کEq�F�E?�����Ō��f��i��"_���(5��׆<M�u��b�B3���<�C�j}�x���އM,��:r/YF�\"��"E���=�v����|b����R�=�W�ta�޶�璋7z[��~�y�Zٛ=H�^�C�o��)��s���=3]���_w$�;o2p�8������wށ8����GyR;@���v�ꏷ�99�������/�Uȳ��>������y222+3]=��'`���*�����CCC��&�}��:wy�?���9���������_h��K��P6��&ݴ��ٓ��̃��%c{�K"4�Z���4�~	B&���1rUN�h�td�#�GPs�MH�3�%�Lm�jӛcb ��q�t�����c��;��]�WٵJDPWV�+��.J=Ӆ?Z��N�3; �#��!��1N��iN+�TZ@����B�vu�-7������k����p�?�꯯�N��y���V���o�w����bS:7��Im�����M��D�����a�����_OA?*�<;��>�f�_��'?I�x;9�Ư��S�c�Ϝ�{7E����W\��h�	xv��ġ]��rq)Ĥ�9��t�`3G"E��$�����S�!�>�D	�%�B��|]sՇ�<����K���"���k���p1���� ��vK.v~�D���G�OS�ͪ��瑧��9�iԖ�Vw�,,縕Y���r������!o<_	õ<����+��������n�D��7�_#���NC��V��i��|�n�m��˜�6q�&����P���Ē�.�B9�����΋@7�!T}��ƊCW��Z8�۰�&F��b���\���e/�;���0a�6&$�"]\\ ��(,\H�K2Щ=K4��w%����&�%ʆ�25I.�;��U���#=�VB��°�F�^�ТT�"$�z:�5�:$N�8۝�a.��i�n�C�u��!��5���bJdVݥU%R[���s-���}��\6�	��!�����՟�yR��?_5��r'�"W����=�:İ��򻰨�/[��g��ot3�55R|!����4%u����r�����`sV�>�p'�Oۀ��M�ŵ�!"�8w\1`�<�*������g��W#�^(�k*T������}q�%��w*����*ɸ�[�Vi"J����ݔ�aQ��0Y���ɧ�a�E]��Ο���	I7�:�����ܣ�G�(�[_6Z����X�{j��y˗�g�Z�U��cw�:�1�%VI�G4:�p�
�vy���ĕ
+;��0i�_��Z����6�M�ǒ�
/�<��@;�DݶBM�U_ Z��՚Ҳ]�>�2�amu=!;��1�g����/5'�ͅ��"=�s�k���v*���G�c����9�<��?��O��s�d���m-���}zG�e��02R�R��}�*��_��5q4y5aC���G4��R����e���W̌����������#oF0����~��Y��@�~�P�vrPk�V�q����|
ћCB�~Jh��GO�r��-u�PIԅ��K����ِv�Z<�ʚZ��M��8E��v'^�48�@���JXc�	�<2"d+�c�����ҹ�4�$�{W��z���>}hY��R%��5��~�q�h�Q���k.�y5
��wv�W�g����ɗ�%+]"X����.��MW���R��3vp��t��ދ���T1x5Z�h�n]u>D4�צJ�ۇΎ+*T��\9���}���i����|�|����(^���s#Z�5�]�vэ���ĵT�Q��]���-�JL�/u|q��dKn�bΌ=Ito�j�S/k���E�^Ws�:�)������UEBN<��R��z}�å)�҅��i�7�U��o�opq�q��e��=9�NC���mP��o�󸈫0#׮È�O� �y��+�ֱ�/SF9���c}!ޯMרH�`�բ
9g���(�Ό������K�M�|q��w� Vr��$����8i��ܝ�;��W��!���@#~^���
ǖ_2Y�C�7H��d���uk�B��X��,ת��{�l�K�W)k�mPͧl%��bdi����ң�LPDs/GӪ�t�m���m����XH�v]�&����wS��?7, �=�Y�пw�/��W'°K�J>V��>t���O�	Q	��+��oP��l�Ǘʩ.�f^�(_ݒ��͂۴���9�}	��{�*��1ۧ$�g"���XW����Cj���9*T1a�T�]sv(	g��R�¼h��-\�yA~</GfKO\N�y��O�0����%�cɆ0�A���Z�����G|��4 �Q�W���q�������=y��e�zf�I�\L^jG��\B�Y( /�{�J�w,���	o�'���t��g��j�M��MT���m'g*Qs�6>��"�ǈ�xo��:����sTH�W�l$�{P9w�[�U�Mc6�of�Q�𴮾�Qu������_0c��+�/V�����[�9���l��G��5z*nI4ή���l�<?3��5'��:�n���&�B*��e)�	}�#���Zm��WI^i�a��-�+�o��U.仰�u~�;?ZC���Ĥ��l�
�D��#L`{�s�7Ҫ�b�}(�4^k �l�'[�l��\h��$-Qo2��T6��oe�����+����z�������@X��-�8�]�i�\z��`x�3^#�]Oh�u��Ls�r��X����V�#�w���׈�\]e�H8��QMu�c55dlQ�㫧��)�V�p��2k���X_���xZ�o#n�M�Br%�$�ƭj�V�/���r���N��&�^���mw��*/����M�x�c�cx���������7ڙ���.9������a�k�H�å9/�#p�7&ν�c������h�	o��PO��S!�҇Mn1�B�8W�RH���K>�_�Q�=�׍��Z;#���g%�G��l^)V,����-��yiɳ`N���Bn!G}���15/qCy=&���4�����dM������	�{R�f��Mѫ|���u�t �`���OA�9�wh�P��8.�g��{��h͗���Xʩ~(9��*�u`I�r	YTekd�qA�4Ds����ͬ���	�=�nհ���� 7�{���BU��B�����w|�gA�:��D�l#��t��CIw��ê#����β��Ȋ�e��RM���v�q�gc��c4�3s��^��b���h��n\X�@�5&��F�/�5�����S���ޭ��f������=xr��[���w�i�8��61�����!��6�%'_�kظ9	kT���;���plX8F?Y���9��Ԫ���P���)1{��� ^�YSs�B���2>Y�󎭭�y)-P瑘�m�vcU�c��G�x�����<�q���޺T�5I���Q1N������;����k"q�.#�zzzK"���YQtC7�4ٜsaxm�X��Ƌ�J*��|0Io�F+WԻ���z4_b\�����FH��f��������@1��:��j$Y�.��+�!+���c��ѹ7A��!5,AK_]�\�_1�0!�Zc�q
1X[�#�&�sL�^`Z���)kw�E�W&ʀ�WY��h����,����%����j$�ZV��x�$Er1����.���[#ۄ|�(��p�Y%a��Z��DZ�g,`�q�ڧ��.���^t#�m��'\�4�<�e�
4�<ahZr�
ȝzz�]9�)S,c�(F������H�<�-9hX�aA��#��lT���oe:Z ���9)o��f
X��լ��W9y�^=w!����%�O��G-��8L�����ۡ���-�p_�3HC�� �)5v���9�CV�+ҽ[�������2�S�u�QUz=�x^R�Sc�O�	C��u��~@$�ߕ9���<�?�R�1�	4�d����8x>�Cn�xn��l�xt�7�X�#ӷ���Q�Iŷ�ͨ~mw�ʍ;��ӡe� ����_�8C,���$�4(�V'2�8�hiZ�ϔ��� ����]�Xl���[4j�>��]�hğ�,'Ʒ���3E�+X��ي��uu��k%���T�;*�%��#T6A��NC�߰��kZX��\j���NL0��`r���Ṃ��'�@�d�����\�Z��r�v��%o��s6�g=���K�$,�ñ oБ��cG���[�l�<�#x�y\�(��[��j�YR�b������m�@B֭釋0�z�e�j����ܱ������)�f���c-�<l,Fs$b��7����69)�	�ל�3�7�1�T`��]�.{_h>yQG�2���Y��y��.��쒳��#�|/K�]�cā<����y��
y�~�4i(�@bg7�rYG��N�r�զ�e�<��E^�䜈J�=6��E�o&b���C�[_���l�a+��?+��d���v)�r��k� a9=�Q�
t$"��	y���5�g'�ȘU�ѵ���0.����f�eǎ����o'?C1�.j�o�
T�4켒e�� \����3ɍ��4ߚۯ0�����=�Z~�ϣ�J�0���A�E��Z,�F[�P�AU�؁��*;�P[�Tp�����٭C���)��������Kx�\�ĭ��܋\L��9��ҷ��{�Q\�ّ8��;�Y��<��T+�a�ǛҷP����I5`��������A���v��کk/��o_��Ӹ݃�|T�(ˋ�.�'���ߏO�\#�����{���/!�`��{�a=I���KA��r5]"��.�FJƥ����B~���U��Zv�Z»�\�8w ���U���9<h���c��ނ�ԓlmF����	Une�������W�@!�kڂ_h ي�ra���03/��w�����{��U� D��rg9�D�~2x%��������@<��T.�g�%�/L����4�`��S_-��^.T���ު �9b�8��� �����tՙ�z|�A��*r�4u�7g�Z�36�7Ns�]f/KK�X����2i�o �xy�d��0[���Q�����L$Y�JG+i��EP��9t=���r�k,޻�2'�9݋9�W]ϧ�`��F�e�/�:a��z�a��Y��w��5#��6���O��X|6��=���θ
�@��Rt�W6р ��Pէ���٘-f�����bV��Ǐ��ܤ��
�ζȖh��I%��#����*�PY��6����X$%�{��,����R��C��`zV�G�b�:�1X}۞�~5�4)XSs�]~� �|��k6D��,��R�Hҡ΄Zua�@�D��amHUE�9��?��A:�*�hQF����^�a�����@X��_f�z7a�k����ـ����d��D �#�h+��0;+y�tLP��֜��������0���.�w����m�m��}@�>���ʒ�wu�Z1����.�[�W(�l<���?39��R�j�{���Jl�����m��׉�%BCbZ�AM����D��bS�*�u�z�V�q�5MBoRԕ�,{i}ix���İ���~��'┋Ͼ��<���k }�j�Y��WGA7�݋mN��?�M�B���[Z5!�4��^���9���`ԣt3������0�z���a@��P\��bsG�����ʂ�k��H��<٢����`xu���|�Q�R�՞Ae<=3R�&�l�G���}Z�j�M	��d�@�"��Ճ�CE��#��4ݮYH�K�T��zh�[�J����(�p���7R����*��m� ��17M�Z�H�2am�O�����1bq�$mc:G�Ve�sd��."L�G$UWc�5��4��!lY�Ӆx|)� )-�<|��ǝ3"Q���C��[��Lu�B7�6��a5��Nꌊ��J���a�4�3�uQ��bQ�yM�e�����f�95u+�x�����h[Ȝ��㒪��5ԵӶ[�Z'������L� 4)j�w��T�J`������1�2£��uO��Uq�-T���Пcgq�;LR^FA]P�ܝ�Ea���[7��_L̟\hԲ?_m��c��EGPO��)�h/�*?�GF=��6 �ҡ��ߪg�y''?��]6��ز��73���*"�����1+_O�(���^�i逭���/�h-)7�(+�����+;PR�.���Ц�����7m�^~���q�7y�j��X��G��!����?��M��vJ�4���wu4��C�j��2� ��>t��7Q^@Yʻ�ӡi|��v;��>J��u�OQ3��5sV�Z [��j���P(����
br��ۮ_`��vKX�C.�Dc�gC@r$�IK���܊��D i�ޏl��>�@u��"i�/`�k�qg�d2��n�G�j�5�(vv����C,P����Q�@�5��	F�7�k��Ҩ�v�A�?X�vg���/�U� -_Mwܑ�7��op�����@��u��	M�.���<�ܫ���5�)���F�NL	 	�(�F˂�2�q�G�W�4����0F'48���H�`5��V��YTl��[���Tax!Ǥ�)�����R��(���?RQ`�>�q�`�a纼��]��.�՚�p

��J����l�����+��/\�Ҿ����L��Wy��H��Z�R�������J��ƨ������v�+�[8U�V�Q��)/!=�5ש��N��;ŧ���zm.�L�oB�Ӊ+�f�����A�l�,��3�i��ã#��WR�>I�3 ���9�$�h͈��O��j��VZhC����^~U���U����ZH�R�3曄'V:�iW��}&�Y��Y�^,�,��ʓw��
l�L����G,�l�	�1bN��&X���kX.�?$x�@b�%P%]�TO1�����P�ˢM�k!���[�^|�;<�I�h�>p��͛�;�U�RKv6�ޗMO��yj���%�K�.cP��k���
���X��]u@P%���c��`�P�%^ JH_�N/�f%�i�q��Q��,O�q������+Xь7�/}��3A���iɕGF�}F����S��u��rer�$y05E���kt�'MF0���l�F�N�v�p5�l���.0��:֬�S�霐�ˍbz[��bH�E|�^	�c]�,P�3����6:��R�ԟ&=��ZF�5UC<�֯_��6�Ar>}u�-��1Jڇ|�㿖�k�Ԣ��ÏT[}��&����4�&��yR�;}ݨ��*�Z[�e�!<i�+P�P��^*Zhw�.����[�f�M�識�1A��r���O���T�r8Y}�ՏP
k`�@.��q��z�U��(f�'�/y��<�_���N E @i����J�אռ����K��H0�m��x�����5#t6�L�
V�淐����8Uc
�8/�	X�.1��h�%4�Eh���v=����g��2�6�Թ�q��=L��j�FOC��4��N�Gծ@I@�@`@]ZI�@g�ݾ�.�R�F!շ��V�=!�#@�^tC�����ٍM:����By��$�O��(4h�n�"F�M��N�M���lm�[E��z�:��%��}Y/��ش���9���R�H���gh�!�t�w��8�D�fc�w�q�hrv}���8�Tt�q��>��V�S�>S+�k�	�Mvx�7֥`�Ɉቘ������Q��U(�!�I6[��]��c5��_�ʷj��j��+-�ǫ��9�.>�幒��s�0�YB�JU/�K<�ڄ^{{����(���Z���4����P�M��\�`6�OU�R#�.�+����©�c�%WS����,K	�m�C���L��U+*	4�O�Z?�|�8��_w�
��+��\aD�I	A��������ܒ��|u�E~?-�Z�Bu�6�A\������H �/#s �W�ďjjO�x�vO��k��7���4�	���C��ayD�6���Y�d�����'Y9���q'p��z��B�i~���S�g�33�x�T��%���{'�!j� �O
��9�4�l�B���Q��V�w0�`���Y��eM��٨g����Қ�Q��'������^g����Åѣj��K�=��j�#HS�����"�!�+�;�N�`W�U���Ĉ��D'���-�r	@�ԓD��gG�B�\yWԳ�t\����s��~cE���'*3!ސ��4�pѤG1�8u�^���P���!��e�e�k�a�9���þ��l�~.Б��zFZ��T]i��+��τ�|�
�R�I2alY�_�'��?$1 dI�92n|VVǨ��-W�L�p�TT�)<��xT���]�bƆ.�B�JHN)We���{�%򬩥�i>^П�E�a_�Ɖ,�Bi`%��ƨ��U^}S���oT_�{��7�J���-Z3��{}�CYAt~!|��Ja��`y�`�R`�S��]3s�$�(��֯_>�6
!Tױ5aa��1�4ػ'g� �t�_̛�=�����v�u����v����gl@����1��*����ꗆ�M��0�[-�lxA;\���`ݼ����1�|p:H�]5��y���yŚ`��GkLô�a���O��m�k����13JқC�Z0G��RG��e��������D%Y� �77���gxAmWk�!���/����g�s�b��8W�|FY��7�%b���
����X%u��>,�֍�_&:�7R$��zt񵒊
g|�u�=䒾/=G���������Wm	��=�ԾR���RB/%;�d$�r��s��JO,���澄��ڥ������;F�`v�������/t�j��+�a����{���_\������_�����g������V�Ż�7PK   ��!Y�R�� $� /   images/179c08ce-6e18-4019-8002-932a24469ad1.png�z�[�a�>XJ(*�"���� A�P:��0�]"�HHwwMb��Cr��l�6`�o�}�?�w]_.v}ೋ�9�<�}��|X�k-eJ

JU��:$$��HHn�ݼA�S����p�榠�w���w���wrgc7�⋴�NO�p��������{w���	�s�YY:�8�ڦ�dHH���|�畱��s7���8Yp+��~b��x#�񋈻�jIPH�i43l�q�Ͳ�SĚ�4"^6^DRd+>�[��:�[�WJ���=I�)�C+Ocy�;?(���(�x��ZBD�$��#�e�0,Y�[曽�t?'��|ߌ�D��Y��2���I�o͕7`�6`�Ü	�����`���C(�͚ɀS�@��2�͸�H���j�~2��g��s������n���������:�#���9rHC4�NM]O�~Kˌ�S8_>��C���d�K%I�:���*E�J�<��:��1�u����o�}w1^��o�gx&d�/7 冞��S[օ��*�$�o�}���J+m��1�b���~�`�Q��&k��#W�;O����s����X�tyt�P�2D�DB�Q�ș�p)�R�!ߙv���ZJtc�.����}��4�e����2w�(*1�l�j�['?Px^�h��WD�8�v��qoJ���D��e�IC�g-��'���VثJEVX	8�����d�Mj�e��=/;��R_bK)��u�x��Q\�[W_����u��PόH��m�w�!#dT�}�N�hm�]����¨!��`i��� ��}����{h�9�a3�eHud�u�4�K-@mɩ�����]���I/r��Q��V�tb엑��>*�O>_;tT��̯�.������+mD.�H���i�l�|���a�\{���U઩<���Z��JC��
�py9D��h���=��R�h�_d��_�P*2�e;VE��iڠW]�
C��	�QF���7|h���A_�>�s���m��i�P���s%N�/Ūj�m��h۲b�-�Ώ���t$3B��v�q�z��w�H7	�By�y1�i��v�S������ߺ>֟�Җ��Bm��gx�I��$�|~L�{�[R�e�G��J�������^Jo%�J~V~Fi�����������������j�vU�+R�����v�k��/�	�0x�{<�!
M���T;��t����P�6�+J�6�Il����Y��ρ�h��O1��#/�ݦ<~�H}��^��(9���OɄ�|	��j���P0c��t���4J��ω�#';��s�޾�7&N�ط58�IB~@'O�l��<S�4�N��1����Z ����Jr�� B��DlR��a��`�}i�m¶ַ� �g�!C�d��N�&�����u�t�������[B�|ȷ��6��Lb�t�ַ[�ʀ��c		f	��ϻEfL@N���qx�~"��4�j����k�n$#i�XW�^9���!��M��S)?��RP��(����a�Ύ�*����T�4���7:�e��š�[ܶ�4����FP+���d��{�"�$S��L��3�󿲋�s����g�k������	˦Z�||�ܕ�k�M�7�����?�Tj>�}-��������@����?9k�<\C.O-�X��E��Sc�)�8G>{�x�D�\��u;7�14�N����U	b/���a�)'�q��"�[�?�}����謁Ow�7�lr��i�����G��1�������]����{?ƏL�1���	?��]q�Ͷtω�#��p����(h��:*I�f�W ��3���ښě��݈:��
�$��̿}��k�4�g+G<�������y�_��4�Zz]�y�$� ��Y��Fk�>�Q�-7봃5Ph�Mg(��(�@�G��ݩ& �I��S�Ҭ͠�U]kɒ&�X�W�����Ͳ4�֎7��O�lB�|鼒r�m�]T��M��z���jP�dx���35ǚ��郁{�+�C���L
o��ezC��&�0�z��B�"��}�zi�r9���H����s���EΧ���Nu�B{�rV���4C�,\��.��)9!�[���?.��+��?&�B����w���,MC��f�_˞����<�8 2^�З��S-Y4��[����;Vk�Jl�9�l��Tͦ�z��n5܃�����i�(���B�/�����v���[h����C
���m�1�JGӃ�-�= ��Ԣ��&(	d}��� ��_u��&v�_���F�VDox���^*��_�ER�� 1�8�O��y��+G�>��lpq��ҋ,�۶Y�2<?��>`$������s��[4��eC%e��{�0�m�r*WB^�(Zr�CFk��퐶�=}@��j�ӫk�c/���3b0|�>�7��n����z&@@���5��ڒ���*q��;���e�7%2>!�1M���:�O🸈�|ƶ"ĵ��:�Q���ojV�F�!�Q�m�Xߦ��砎��|E���0����8�Fx�<�6�^�cb"���/�ώ�-8��V_�I)?�rܒ�p��W_/V�.�8���9<�����	ƒ1�����]�:9'u����f�YD�Bo+��wwz�uv��x�_܏����_L�&���L�^ -��Z����D�[�ˈW�	��n3��5��@�n����R�9�����|_�=o�9� �~���+�0z3�=��9m�Y�����K�W�HHb���* x�݊�5��N�(�%��l�{-؏��K�A�rb���v@r�M��c�l�i���_�Ħ���O�Gr�'h܄Q<��h?�I�(� y�X��8@d9���~�/��]C6@�,��ko��A�u?��cUA맆�57�@�y� j.g$"�$� ����q�����Ib�+f ��c���C��̽�?� B^�^�2˯���`ׅsMi �2�����XyFԽL�L�s�g��潓7����)!m�
a���s��|���eNo�*(�m�{;�Ϫ%�?Q�ǭx�g�a{����	=�LHg# ��$4\�^�sc�cѺ�*sgti�*0�A^^�3���Pm���������%���?�n)Uگ������Uku/V���B܅x��@}�ԶWQ���%��ZJ��3�fe�@*�&v��%.�r��]��F�SmH�m��,<�}/���F�-�ukgV���6�Baׯ��U����*��j�]��o(�I��$Z)�����jj)�]���W��z'���]&�ɣ����<Ęj]�8�p�K�SSS"�p������4��V����.I�4�oZ'Se����%�7?�"W���.2����X}xSHƹ�Ъ!Q��;��
�L��F��Z���Z\���N?Ӹ\�J�,�)I+˴�*�4��ſoJ(s��?��V��I������<����B��7��p�A�͟ô�������#$m�
F��g"� �����v����>���������#`�E�xk��+͹�U�%����Y���\���ن����~yY66�MR?p�����V����r�t!TOj��ه�ZoC�وB?�Zo ��?m���q��������l<���DB�S�*��2��B�;!a!bS�-[��(v�Ԕv�VH���5he��k�O�-p�"� i��X���풏���/˟�i�eVؿ.�=�x=3#��ŝsK֊�O�Xu�L4oH���E&l��X����b�*�}����"�Ù٪�GzhS�E	�{+S�ƥ*�1�_̾o$J�=�I�ıE�n���jI�r)�g1'\f��ޜ���@(��
��ɤ�*w�>O�)�-B�'��C��L��ŕ�&3ZY���2�=��$�#ގ��|���y<p}_�3J:S�mEE�x~�Yn�����/]\R�s����ЍMa���&x���4�x�	dR�߰y+�կ#to<�1���L��S�j�������
�ﵖZ�iFr:I��G�����Z:��P �["�����{;q�%��A��"������)w��%�h��̎%��k�:13F&e�m��>�tBnn��qiԖ�ƍ�P��g.������UUL ��i??b�g3� �*��qfw��1�ٽ]�����
dx�E�C�O#��D���		��1J�+�a��Նq�L9���rx����bRի3t�Gژt��
�����N����6~�� g 軳sF���.�:ߗ�xN��[�dM����@�>|��;l��Z*��}�V�R86R�ȇ=r,[�J+s1���~]�d9�{��V-��㞠�+V�S�D���'��3Y���>�e�������k���,�T�p&xf�oȬMı���ætAoL)�e`0G(�����c����j���뎽��� �4�����^ws����=�d(+��Mē���+�n��M _ȿ�u"��g'�ʗS���V�l�p�k[r/�iA"���1��Ϭ��o.���Y���(�	�R��4cc� ��iPP��45�o�[�B*A2B#	�t�� �gs0�PAD���:n�j�:2)Ll��q.��/Lk�fR��;3�3�������*�zO����c���.�ߙ�e�n��{2oMH�n���^'�'��8���[�l�z�3��Z��4�-�$?��P�ޢ��Ym�s�-�n/�z3��pi[��k��@W�����������)e7���u�Lr� ����ǣ\H[)�K#�9��%���m��W��
��Ñ�m��Kb9��˸e�bJ��K�qIBJ&�r��VG%��ilf\>Re�mKX)D���oS�W��1���MF^x~}�V�k�h�x�`���E��I�T�Pl����{l��br��կ[\k'��;�h�&�ۓ��\-���ĺ����#3Y�·��kߪd�q&p�ff<���O�͏���3`wtB��lEG�"[Y�/��p[��4�}+.��	����҆���TȰDE���y�� ����O�8yl(C7�e�/��(�l��/�/�Ko��L[h�aK�]8�=��7�^%�o!bx���챲�H z	6���q��O������y�}^܌�[��L��E^ฎl�νļ=��9� ���L]��=�^���J���+�&�����f��hY�%�n=gRP��	'�vc������1��b=@F˓�;��'
�};����$�*f_��y�֍���&�~jvˡ�o���ml�&:��� �.q�g�s`�Y���K�o�掉��s���..?	":^�석{��%�>F�N)��1����	����|O&�Rqd�D}��9�V��3W6�1�;�������F����G�\����Yƍ��l]������P4f3?)��T��z�����ƪ��m������;�Hxy��W�e����<���d���g�z����Ŀ[�"fDj8Q�g�=�X�	�����`�mfh�����^�v �_1�@�Ǆ@s����&���S"�r��� �>ٶ�*nw��i��|��������-c*� F���ý�*f�1���)j�Z��u#��i�l�����I��	���)z�\��ޭ0��b�(�|��w����w}�,��,�Epl��w]u�tj� >"�޲HB*no�_ ��۟!�o_۱�43md�8��#����Xկ�4����;�v�{mcY�a#�M@ek��O��ʴ���b��)�L	I3�N��Ģ�Ed�3���))�:�؊0d)�L�mV���6�m����2��cآ�V����*�'��Ɍ�ꏈ\�#˸t��6"`�s\��D��x~���+g�<h���HԻoj|���J�0@�[�,s�j�Dtíy���B۸�m�pLV��{�[�3���/h>�&�2M��/!�>�|^#4�YqsJ�[T�TX�� tgh_[q���S�EE���N��_�P�Vn�&z��~��Z>�$?o?m�lO8:t�#}���2㏀E��T�@��F�'F�R3�eXJ�@MߟY�W joJ/lr�J>�/h0���>�g��|��#h�r���9�e�Qlrz�Ι�j v@�AN�P���=U�jc(S�}k���NJrϩ� �cG�/|��Ouԩ��I�'�E���DqLD�$�����Ü՟�C�B���=x֒�K�堟	r����s�Z�cɷ�#�aPxy�@�5+'�?h/N4�c2j�"��H��k:F��N�i���J��>_k�p��A�T�]���wW=� .-<P�L�%Wa�	И+��}6��ǂ��g��*�9��?�5β=J|���7�蜋MH4�]f�Ԫth���$*��*%��W�1��A���3~��(���Oެq�=��R�51�)�y>¼LY�q�K�U�$�K���^�*+Y\�e�*	s��|*5�6=� ��^%��6o]��؍���aOsy�boRB�F@�e����B��$��~�����0��+�H>?��8U�yA3���˓� L;�xn���r琟��s�.�3���"��1^̸rriu�A��w��l�	�A+To�c��c�;҃������]9����%_�V�^�|&��p���#l�w��k$�?ܓ�[���!m���X�rj��#0�X��|���Bˢ�ëMF�!ι�s�ܨ¿��]a�.��B�\��{��44�&�����l���|�]0��Jrؑ����$c�rz��D.�MB��

�6T	�����1Y�3_��� ���K�F�ŝ�}N�R��~�jQ^�&&�-8�|����K���N)�omo�>��-��G��X$ob��@�`����n=�}=y)�=�j"���A%���//*F���pC6_�N��yPf��X���'1�}�3S~�w׿��5�����g��T�\�[���_�+6K�|��"�b��U|�B�����?�~�
�/l;�o�|�-h�D�H>��*L/�)\F� i����x���\͈D���xzs^;3s��r�G�)Y����K�+$�/Q�!�p������}q���9-M��Kk�c��sG�i�}_i��v	]/�G̏��L~�(� �h��W��:�Ϛ��\�(�8��r���#�$���4�04�%av�cZ��jq�?�k���ͧ3�9̫i��g�Ԥ�Ot��-�߰��|L�]�!i˗�v��gēe�[I����;�����n�Ph?���w��f�bE+�y��ch�����9�!7Rv#�yW�.����P$}t$q-hN�QFu�,�p��f�U���jnFѵ�ٺ{���o�4�}[{_����%�-6��1�]0P����N�c,�߽Iv���?�_^L��@�:%����'t�w�?~	<;��_�`Ys�
x��ӓ�h�O(-I]��i{OO��K96�;+��sVX���@�Ǣ4��7gc���:�@�'������f�l�Y��w��.nLv�?�s���6A����� 4����</&h}��3�5z�h���i;����V�mQ �S���u�y����Y�;���jE����ư̿�������{��b/�w��[t�̀�xb�?h�)~t��+���N�N�a�g2�l�ڥN9�҈b�(|�MФ����la{�������eIY���Y����T�%�;7Ь>%�~?�3-ϗ�v���2�=�HH։��2g�P��p����F�r�Ys���3�̉�3�����f=��E��z<�V5q�*X{s�L������W��2����5�q��D��r='02|>� �ڈcP����V�	�]�
���T�z��ޭHQA{�'m�4���&+�c>�n��(;Xp������1�v�m�iIH"4�	�9����}R�����a���;�?�'H/u��(�R�ꬲ��d�p�>���3TM�X>4���g��U\ⶳ-dhO3H�N���(sl��<����~ ��k�:Q�E��G)��`O�b��H�XIP�H�f�:���~���Ox>�9�OQ����Y����K����o�_���r��6�� ��K�mZf���xq��:�o4��gd�i��pD~����;i���{�u0N��=Zy�[V,
�"� 2u�R$8�������N|~�Fr��G�0��ar�A���5�|�<#�2D�ͬ�LL������f.���Y)o�{�ڊ���;c���XQ."���LЪ7��߾8U�_��G����]Y�Dc��D8�׵���VY�Z��K�Y�A��X�R_�;�>j�K��VT|_�m���H9��y�J�!�L�\���7k�ݫE��ۢ�b��;?�J�0����\��ۖ"�\���N��{ypd�nx���h��3�yJ5Eg�)��VN����{X�_���3k��<?L��w(e�BD���S�]<�cZE�Jo�:��jC��Z&���x>�Z�����ǣA?r�Ի� /�6�ԁ�,m�������_�̱հ��� M	��� ��G_�M2����+�J������e����ڎKe�k��Y:��@*KT�\g/�7k���6F�;��*+�777׹o��ԩ888؃@� P������TIR�U�d]++����oz�C=��I���_�WL��Y	� R�f�n��~��wTK�������(�yH@%w}�W�/�����SWL���?����~�.`���ݱ�Z���-&,�6�'��5'�)�o���)�Z���ȑ��t4��r�"2X������"۠ʬ4�����`m{gG����0�t�D��ۆ�b���|�@��/�_���{��O���f���)��Q\�M��=h�y�'�*��K��7O��Bt3č�Д'y���JFC�Qj��H4;R��L&�ԭ��H�k��+��Rg���_6JJ�R#�0#�X&�}�r���}��ƵJH8~�AN���CCC��W��;��m�p�q��,�ƺg��o!xg@~w�H�A�c�r]DkE�wZ��³�zE#3��[����~V�#X��4R����۴�oe(�*���������ǡR��s6�R��߁lg���_rs���߾�'ƕ&J>�gv;�[/��Med���������R�L{Z��bNC����6�#��{�^�L\��z�qn����\C��F�߂9MV�"��[�L�ڊIH�dJ��+�GSEl��ٝq��7��'&
��I)o���bt���՝�$M�6��8���&=Y+�>R(bS��ȧ�U���EC9�	f�O(t/�r�|!?�f0z4C�b!���)��啭���ܱ6���D��� �2���-s%�"�b��-%-u�}��fN(B���a�J�͠�L˻dMkj���'[I���jΒ{fy���f����A���|I�×cL�
�W���bf.=�2���L��ܞ0��8�� |�=�Om���u$$��ú�n� =�۰P%��mN��� �������Llvƾ���6_ؔ�����;�cƻ�Y%��Xd���i�1��A��IB��"�d��</��_���cF��>����+�g�i��uN�;SG)��;M�����O�	�w�5ݷj�����|�	�R1+�5����C:��:����HE8�� w^��$�]Mn������H�������<]j#ݕ�yac���,�,?,���
�����h�j��P ��ŝF����*<��7��$`� ��77q�@_�I�k���� ~�f���aQ|�EGfYEnv�y���w���;c��E
p��(�U��!Ov
=[�q\��#t��&祐,_��?�0Q�[�,P�!TAٰO��\P\�L8�E�в�)�ʘi
�^��^���]���i'�dm�f���*t��2&C�~{�m/bT�HP=>f�����U�<�h7�1�P�R.U�5��>�*'ҝ�J����3큁sk���0m�W;��}�����f��_�ո-^~e�X}�1r�v�K��c�|�2�����ϜӁ6K��W~���[ِ�C���5�{�x�T�@gy��V&{:MF�Y��	5@�Fgy����5��\k���o�R�Y�6{ �:�^6w�+$���t 
��N��*8.�p#%�,Y����zB�o=\{��,�g	A\
����R����_�X�tೲ����V�e~#�f8p�.�^j��c�6I(|����͹�w( ��i�w�g7?���Qv�evY�@,��r4�S{3T����c.�JJ��S�L�f�� 0p�4l	]�����$v����lbf���&?q��vN��$C��2cw
�#k
��6x��:�UT�б7Rq���47����S�~e�����״I��0K{n2.�Q��<?5&�!�J{E��dd/�c��Y'nb��k!��~��v���-u�P���Rއ.B���W}b�E�]�8W�8��^1��#��7/�@	-!!���5^k~�!vq��7�SZ �s���"�?F5-A-_�[�^�gZhz��4�M�9f*��"�P��J��g�X�Q�;���ĥ|������*Ͱ�і�M������]�eJ�q�\G��80���ӟ��H-����RSS�%��xf�Yh}��b��N�m�U���0C9���;��U�m���ڸV�5�p5��5��������0N}�A�*;������8�������)fg�+h.�����2|W�(�|Y����<�g�P%;��R�
[�p�����������;^d/Z<�H�,6WD�ͧ�>�~�K�uZFƸȰL~;�>��j=�Vp�@,�fJ�`��c��{�e��׆t` Y��o�6x|���ܳ瘷���:��	O�\�(��W&���ې�>��q�n�,����/�u>yG��y!i$a���٠�j���!K"?0�O���?3����%Of<f�W��y!o�
T5q�K���p�X�= ����|TW$���A�������أ��|���t����Ψ�s�˰��k��uH����V�d�:�����n��0ú���l�4TS�,U�5%�5nB{i�
Gg�R�tR�`	N٧���m+3b��i�a?���ݢe� ���~��_<���ɔE���aͭ�����&�81�IU����8+�
�c�ȵ�H��h��Rn
��=�,��:{����z��?���}Lhl��m�0��-�r(T��<6*Q6o-��c���@#c[��oO��~q�*��������S��Ui
s�?���Vl)c��Ǥy���w��Y}���ċ�����ew�3��e�7����R/{���D=�۬��㬭*BO��y��9NhpKW�:�f��?5�rq x��p�m��Ż��#���E���i0�~���A��q:7�Ct���,�l�&�����d2y�5���WO�k��c����o�zE?���9�O=�(fƼޕ�#9��x��]�/�GÃ>sIE���t��\�<�ǳ��Ke����(������@
��eU7�Q�0�H&�5�)]�o�g���t�[q���@��E����Y������ѻ���1pU��(:樔GO�#���)j^����Osp��/��k�:ں�� 	r�g�l玌���A-��9���k̡(7YG���k��5��6�1�ZT��&�˛��>$��i	�~���7���2��U9HI�<Γ>y��H_+7V;,�~������z07�Q\�߱b뤖c"�lb�o)�Wg���Ò)J��+���0>�3��&>��+����K~ʗM1��ù����n6v�p�Mf,���r�4́��U�Ù~yeR�_[W�S�ŝ'4[B@څ��"}���������/,"7�].�m��,t���X�:X7G�]��^#�76�'�1M��Z�I���TyU�zn�C!���x��9���'N�H���gq����7BZ�R�[~	����"�� UC0'�O�r7���;�,�x�<���c98�/�r����O���fV�r���S��!N)?��`�'<�cX�@K[���/�2I���vB�8@��K(`#�������s��<�(\���'�EjoVE	ک�O3(�YS2\�����?�ҙ�ҳǣ�ۙ�A\
5���syƌ7(���d�,r�ʰ��E�cH@PiJ�;�Z �����Zv�cwVcw�-�#ئ#V�� T�Y�A�E�ak=�>�Оr`��Y��aZ��!��[�i;t�N��"���)� �c�r�oZ/��1�z��wC���Rp�c�^�.���ڦ?Y�%o��Zj������+Q8ʟ�}�`��P�^eE����0�����[@@ ��㉻/���ys��~tq4M3aX��s�"���U-��J�#��Ƭ�E@��^��,�r2�4������Fa2p�~ᡩ���\���qUYYy���-g0]�ۜ�r�s�Y����]�M�K��Н7�i{�sÛ놬f�㨀�-akc�j�Q�c�z�n���J���ٰ���	z֜YĄ��7wn�� (�/�P�������t-�~����u��;��.X�	�$9�E4;��c��n�[>Q>=]�f
W�ݎ�,�'�Γ���8��t�����1������;�9H�Þ��da]�sY�y)I}�6z�?B�%��������]�Wks�����1MW0��1 c8U�䣉�3�l'ƍ`��L�X�b����z�em�+2�n�-&=� =���ɠ�m�-�r��Lm{�4�D����ҏShK���O��M��f��T~�*�9��U�=����y�&��p�4?��/���e���l,������g��ڳ,�6e���VP��d�of>��g���S��o�O�T�KZw��Yx�����az���3�`,e���"���+��|z9��^��k��,� }�{� ���hP�Jύ֚%ͤF:�E�j�q������,��)��3ulz�����������F�/�^�/�p���5R�r�����Q���r����<Sסp�ʦ�)�Ԗ32�D�v���m�, z���π��J\1d��fj���<��ڨF�;�adDXk<Bw~[&vc{�w�ۄ@M���o�qpx���w���ښ����d�4�AV%�L3��I�)a�ih��OX����&�J���p��'��}�-��o��5��>Mop/�\�&��|�mՓ8M4�9�{��*V����<;�A�U�<[7�����S�ǖ��̡'�a�-b�n��M\uL�l��F9+��!���ǫe�UH���Y�aZ�7�T�Nao���.ޘ2OyO�Kw�3�R�5ͅ��.���IO}!U.9�FZ��17%�=�������,�� c������u~�����W�H�
֝��[V�lC���V߲��ɡP�V��q���e�ǝ`�L��S���g�tu;ٶ�9d�t	4��=��G�xܯ)�yم~u���<H3��?����m�0�Ur����@�����#�öK~��֤$rG��,�:y�_������ ֣&o�ң����~m�x&�K|_�*����f���s�X�X�Ywm��]��i<S���O�&��CE*o�X���x�l�/L( ^�&���1�p��8#�S,�l��qo�u�Ot��M]\��4��jeV=m��9�T�����[��~���R�rxV��{�/����y��t�L��u׻�]ކ�#���n������?�����@co}��N�O���[n�,��+<?�5�<S˅����Q�2gۥ�B��}��{ukV�����7��>��v}�Y��B�aM �y��ܮ�8��'\#q��hq6�a�E����%�Jp��C5�P�=����qq3#����TN�����u������=��	��f�]���n��ƨ��&t���.��㌷㞺kU���)�R�n�>�6��F�߫7lm�+�xϣ���7���Z�����[��C<�O��<�7y����(C��'dni���I��3�W��e<X{�M���yx��q�q��1�^N��U�U�<A: ��K�,�v�uJjj�n9�b���0�����5T��q3%r^S��j�1�i�����]zɧD#Wxx�{i�&���_&k���QL|
���i�Au7�nf\:?����7N=�2F��2Ř㜍��v�����,�����m��}ZT�%�+�K����/������w����'(���!��追��tS,A�Ҟ;�.֝�ܹ���5���"6KpSJ��Y6+{��Բ����5C N*ך��x��ڢ�F��1VIS�B|%�rZ�n��!�{;��P��m*���� /t:��26��8�͵�*��'W���=~�u��̧#�=I~�t<~�^�^�\B^{8�5��Ű���8����{���*��ۀ�����[��Rfւ��BY�z����?�}��P�G��g�7	�P�zr&c:2�����Y��V;e������!'a���ϫ�N��tb�,a�5�u����t�x�ݶ� '�-�������C�i�k6�I��4t|�m�*@�����.�r\>Lp5�0=õ�L�:�(�p\�6��A��î{YU����_�x��͔��-�ž
Y�=mp���~^�î�}s�\�cQ�ٳ�������q�J6�R�,X���{�o��&�£�V��#�Cr%㖕5��� m���T�j+d����?%k���?I���C��d66��x2���f�)֘=��L��ϦB@u�>}�"�Q���vC
�����ʚ�n�pB7V�3Z@�y������<h �@ō��ʉ�
���P�X�a .�8`�w�.�XA�����H��ǖ�4!��1��(����Q&�PB����|�`�K�;��gw��נ��-/�G9ٶ^*ޜ��N����#�<h �q��s/��ϟY��^�O�ޗ�4Uf�Ou	�8k�*�LM��,���+����X��0�h��0��ؑ�:��>Z��]���Y����!��U<��j>\��x�?Pm�S0[�M�1g�On7P�5	�w4
��Mb��I;���*���n3�Ά[����mN�N�J�������V���qZ+��}am�] �mi:@�M�Է��ThY�r�L��c���g%Ir�_����b�+X7~�PvJ�k|�#߽!��a�>m3>�<�ۆ���cn�V��O�$O*��=����6G�`�恉c\3���ɚ�S/�G}�ǯ�F
���]�	�����|v����^���\������&h�H�J�ox�U�v�l\�A^e=">�A�mH�$�<�i�5�}�wL[��B5��
�8�^ �K���w�ʤ��:���S�[�:+Bհ}k��= ��U6�i�ъ����Q3TVM}5�%�z��O�K�!�j~Er�{��mp�5q>`	Kwe�g��g���b�����,��OD3�=�Ҵ,u�D'?XLT���@?�zw`�5ͬ-�W�A��a��_J�������]Ǻ���L�~_�I��)����i��ֿ�1��/~��r
�����{ul�m�V���>�I����,5����*�O��&k������`��w��L8��e�����
���ȿ����>}M�h{�?#'اrɇ��W3�����
]��Z��Ms�E�N�c)����S���ק��*����R`��ǇQ���V��N�M�)!�����OVټ+Mm��2��BP�)���@�ؼ�B+�$(��z}��Y�vV�0��."K3����Yߩ��~([�,)pU��,�(\����1���,��ۏD&ݙ����R�C>]9;N-�rU�5�"j��;�1�kv{���O�.����8�U���^��vL�U���tS֭�d���
C�22��]�)��y��
��K�K^��&�>/8�����b��^-4�5T�1ȸ���,��U�6��Ń��㐹<�*t�b�ʡ]�eb�������<�,i��p�W{,'���,F}^0�␿>��e����;"��^/hii]�uy�+ך�m�)lmv�7���:�@c�ѥ����|��Bf'��/�3�%K3����L]���e���k�%��"�v�e�R��5]�'#�cx�z�e��S�|��쎒��O`���g��pw)-K��O=�
��n��� �(E��&���7E���Yϵ$��F�>1-���n�y�y�2��7	FN�WUpa>>�T,N.��Һrf��8I|V�)ا�\Q�F�k��G���3�������x��d�-��l���SΧ��g�Q��O������&���$�f��6�x�/K\+E������xrV%�y�q�D�O1�q˒�bD�t�81�N�+�h��!߉ى�3?6���)ei����;��*V��Ff��n|+�����鲹��51����U�R���= e>C���lA��b�܀�₆�?�OF^��Y+&300�YuG7��^'x�k�NYg�������i�$��y�&�d�`)���y	���_)E�+��H��_:k3N�m��k�ٱp�|�\Ф��ǔ��h�oM��������X� �����iW��%����~�m3ݕ''<���g�W�����:��͟����N8L�5 ��r�*M���>��4� ��t�[��܇��AE�mOM�$�S�,,@y�}���Bl��@��<N�a��%���V��/�w��>,�a�&��hk������2Zۆ����%DZ����chD���a�:��������q��9�?�\g]k���JU�?�y�9&ȥU�Pښ�*-�D ;�Bd�$d��J�v�����g�x�
ߡq�wt�{͘��%�{F�ʵ���Lo�,VE���%�����������C���J�w^e�8n0!�ϵ��i��O�n�V��n���;����y�e�HJYѽ�̀����5S�c��O$���G���[�Y���d����R�խ=�>�f�O�m�/z��4�A��!ϧ{>��͕�?ܜ�{����~l�'����{y;h�L�ˎf5��u4�%p
�69ٻ������Wo/)�
9�:F�>�Yڸ�q�z�L�c������Ҡ������*�o��}N%�O{?T"c�#c�FaW����H�V���}���h�k�-=��(`��a|�o�k�t�_gT�O��,}P vQ�p�+(=�ٸ_Le���gRtV+��*˳�vD]K~������4�-Pa8!����������/��k3���t^�2��3!UӮ��������M��gj}���;�T����v����S��x9�ي��w�OC�#�68P��o��󦐪4�G��X4�I�?/�SVcy�c�����C	��1ڼڎF�i����"�t�)�J��U=꩙����O�HcB�O6����^�=����
WCf��Yony��*
1�xC��Ť��Kү��b�yE�+�o���gM']�)�PN�J����^�����������GF��Hǎǫ�a�~]C=�D(Ҫ��,�a �����K��T�i��ҕ;�0%�p��A/�0��?�u��Ms���9g�����[�
�|rj,!|x
�`�ǍV��6\W'T����V��?&�|���]�!fb�:����0{{�Z4H'�����=,s+�6���'�A���N:�Y��<~4���b�@aQ����H�:�CU�{툃��o�$���g6ob�}���Eڸ�{��g/���"o���
a�Un�'J=ɗ�)�3���A^]ǿPx��p;ֿ]��G�|�9d�9i�j��7�M����;')����� ��)LB$�de7���v���lt���.a\�5��q������$0`�r4�~{ᤃ��l\�[r�2vU6�&i�|,�����ȯ�F�:=�m�?�����x�>��{��4�&� ��jo�s�����"͋�FNwF��l��u�=+�S1qY�+dC�$�f_SB�4��u�E��~����4��/lGǳ�c.�`:�>�q�����r���_g�gQoy��U�sI�;28}�v
���������,�F�/�\���s������);쾖?Kfk�y��ZQ���j�x"��C�/�u'�G�� RB�{4{#�[���Q�ͭ����%�ʩ�8��s��������^"�xk+H�\�v�X���N���X��b��.ƞ7n]%dk�#���k?d<���}��I3��k'��}����s�+�iWKN?�Ok�.i��I��(	��Rӱw?�Vh¢q�4����Djp���C��C�g|�@T$^;�$n��>���kM������ok��fρW+#�gbt~�Ǔ�y����y�Q0�b��	b��#�����Xo�]$�n ޖ���L��RE\X��D�(	i��u������dЙ����t��oe��=:�����}s
s/��V�Ju.˯��u4�����:������$����hiAOߓ~QS�Jx�Y��ͲM��8�k*��I#\244<��;m�=T���q��zc�v<�m�ے�M�r�������NZ��PSq��Nr�����n�>�F�(I�`c��R�)���gaZ4�Y�D��8t���в=0�$er�p��,G'[x����@�ֿ��RH�놕�M9��Lc���=�ݘd" ?��Q��`m��n�U!��|��x=��*�$�瞇ү.I�ʽ[�I���5���5���s�8��s!�V���Ե�J� ;�5��U�*�!K#1;��[s+�\�[݆�p kMN����䎏��~���~��3���H&<�=����B�*-Q��\~��xk�sr�ق����Y�0�ywY)n�9���R�����C�G�:T�9��l��5,��[Ѯ^�^}<7q�k�@j�
�U�]�.�w��4Ɖc:��-(=l<pi�~����b�'A��	�DL;�����װ�QLL���&'E���o7�e�܅b���74��(~�8c^�'����@[�yN(��,=J�/�K� �� �/5��J�7�0ˇ��;, a�����m� 3}�1�։�ܚ�Q-�ޙ
;��ϑ<�ݏ!������K"u�LXZV!  ��(|��縒Х���hC��jW���*6iJq�[�.L�w�d
�1�n���a�r��Ϻ���/�ey� ��2ǜpX��0�.�!�n�y;�|F,\A��)��>���4F�x%%�"��>�&�L=z:�w���JM1�n����m�~�����M����-ⲁ�K+���1�++<"W�	�Φ�qA�O��Lb���ZY1a7�]��@ ��ɤ�4�pɵvrR���M���WCQ���H�hz|���>� ��%n<����+��:y���7ee�^�ZS��Є�Up�,��3֗ QI�I	�1�>t�>A�������>�s��n�5�v��-����@3wQ�p�g�����+�^f�Ѣ�d)v��QC�S��-D�O��I�0ON��-���_*J^V^}5i�N�ɩ�z��s� ��:@`�:�?)o��+�Q��� ��i3^�e+_`�"��6T徯����D/:�7A�������(�{��#� 4�������_mm4��Ʃ�6�,j��D,���W���(�� �"�n��6r�P9���_*�/����f�)s����m(���aM�\�M����E�(�A��֎����L�`���SD	�航����.�h�Ƥ����e%�Fa;N�oP��0�_�&&��\�&��1��8�[�@3�nF�{#j܀G���s|lj����?�(߭:�q��ыF�ef�Ч�@i-�� ��N\ϯ#��}}����EOHT��;��0��b��ܜ�xF��bH��T3&y���՜+�1Q�ΒrT�ؠؼ�B���s���xc0���xYV�+��bO�Z҇��X���P%S�`�P�?�B����mBڞ�T������xX���y�׿t2:�_WFM�l�'w���o�D���H�/��#��qv����N}�OT}Qu�T)�,!2��]�(�I��0g�>�ݳ�g��Oy��xٹFz�B3a��{�:Γ�g�V#"W����w'��"Oo�$�5���Nf��1�Ӿ�T&'��]c��m�Ej���6��p2g��hFA��d�����l	��0W�k,3Q"t�~��Z�+SX� �~�-�#� ��<����r�F��+�\�����|���3K\܊�
�g�RE�X,�2I�$y;��]�zS���朋�.�v�i�G�9�_Ŝbf��y��Y���u���3�CܯE8�����V�TV��-gj����S�fc��T��9~��~��G"4ΥK?�8��@ �y��R�6�]���g�^~^�G��~��9���qTl�{��C�!5�̏�v�*dR,��<�H=�w����{̗�0$>� (�T�;�S�般:���Ws^w��S<��ү`���HF ߟ�>���V����l�]����\��@�â�}#����\��5�Z���5�~���'¯�&��se���J�b�ܬ��,������U���) Si�杘��Q�ms	�/xq�^�&b�;y;uz�]b����zGt���@i��\�^?W��ERt��㩂�7t����מ�鎋k䕴�V���VF�Հ�L��^�I�U� {�1�Je��ˍj��=_:��\`�yN�o�x��W�fSo*�,�����4��T��&lU�M�W��D��x} ^��,v�����~x�u^���M���fU�$�)0�����h�Q��7���jă�z�����0��* 䗗�@�Й5r���*�Q�éW�Lh���4��&S�i��ǫ�)��o�!�;�'�1z��$���=�)v"��V�J�����z�V7_@gk5�+�Ƨ�Ϭ5��71"���\G�_u$'��b��]t��8&8˒�<�Ͳ�KJ{c ����"�Y�_0�D�)�n]A���+�&�+,6�����v���+i�\���8���'~zGAdǥ_�+
��C  ������a�����8�w���@"!�|�Շ/�>�����


h�x����1��@`�����K��n��Ӧ�#�M�3<K�^s����)4k��������<<����~��MA�oO���&މ�'w��۶崂��_�%�#<j��"טr3-J�C��x�"_���(�r��n��]�T��(B�)�K�_1��[����- ]z�+�;S�<����T��x�?@~����6�%�GF}�����X��|+h�yE����.[!P�YNy�!wCh">���9��@��]E�CK��E�m�'=$t� n�ӡ�pr��������x/x�>}�?����H@�J%��ٖb�����I�uDY�������o�T1��dZQQ��}����ζ֍�&�M�����z@��ژ��
c�l�����L�!H�n��R��#殞8O�]��-�l�̘���٧C��Y�1i`h���-h��s�2��UZ}@������U�v�K��Z9��څ-j��6JN�[���o�	����*�-K_��~��Q6NR*��"��o٨!��ڪ|��K�rO_������F��;Yj���y3�?�ƸH��@�2�'N����6�Q:����^�����x�J�f0��C�r�n��l�l	
�������[�Ҋ�X>#�8���F���s	�mN�w�,�!�Ζ�}!e�1����A��&���:�y���L�m�_T����N��|3��g��h2�߻]�9�~����G�z���t��$��(�x:-��&G��L�7����Yj��
g�򞉪���[��]���SU^�Eҗ���Z�ۃ�h��&C5�2͢vk��R��_�K�TB|ַ3P7�D��!��;O<��q}9(��r3@�::mE@���^��6p���$|jc6)ca�h9���E��+�Q�F#��]��v�/��<�Y����A�������c�\��~O���j��P	��Wy�js�vǲ�^�±����wdŷ,t��Q�ם�;�/e�(7��m�6!1d9��\�+���p�d^uǕճK��wH�F��ϕMj�'�D���hhp�ڥƩE/JK�tl�CEj��#]�i2]������v�N�+��N]�6=ӛr戓�V#���pXFrϰ��}P�sg�~�'牎��<�2�»F_)�Ϸy�~'Lن��4U��D�A8��E{���q��<�_�O���lmm'y��_m��^\^�-68ؤhB�LT���A������㮴��̠���!>�����]�� k���Q�-l���ypc�I��;�ni�:����X��Ĺ]K��I��&C'��#���I�<Ж�פ˴����Yn�C#c�����,W�rΊ	w�I��3T�r>���/Ge��kKo�=T�m
���5��b�ju\G㚻`DP���y^�g<�����%6���w'j��0Oq��V���Ĵ�|��g�W�t�$�t.���_�#��0�Q��I ))ys�ґ�����F=Y��K`0�尼�E���v�}qW�fa���b��hC��3�9�÷��m[�Ѕ��VT@yj�d?�!x�nQJE���$����nװv��q��7ݷ�.a_��+l�g�7�>�B�{����y�K��ܿyy=5����6F��aۑ���\�y+�笗.K>�o;K�˪>��R�}l/#`2k��Eo&�݉<D����Jk[kc�'])�u/���q띇����7�%��N�[N3�ֲV���M\n`f��5(���+������𚲼����gN�O�Ua��A����.8P(/W�P�X����	�zq}m]���tD�fݦaL9�5�Ay��i`m;`eT����\������3 p!5!�������Y�S# y���U|��A��:^ a%�dn����}�{�� �/�A2W�
R��L�A?Y�'������No �����'� ���aB��i�;I�<R'��q��]Ҳ�EM�)ݼ���;�&�|��}��z4l�)���p:.���q���`���|�"���b�$�%L����!{��\SS��UU�yy�i�ܻ�Vv����\P�C`o��a�DEP|b��e�����w?䑼	�5��֞`3a��:N`��x�u�H�.cGw󇣂ȣ�n���L5��G��W� ș�b��9�pj�p�#�K⢩`�:��<��$ݵoCo��-�,�8'�9��T�D���G����Y��8oweV��9�W�]���䁜��P���+{1�Rg�n���[�U�V�����R�JH�����J|rrrݰkU�ݝ��R3����:����Ȟb�$K)p�1+'3��bh������0�eK�Euyl�x�%鰬 �����[�>�u��_b�v@?<�1f��dH�.̢RK����b�h���	ͤm��Vg���f��1�h����'h	�J5,����"Oĺ�8ҡ���1xSڃ���F���j��W�
2����L�\�'��Q��������ϕ��y"�#���g���l%�۽��W�ڴF�48~V�^;�Eհ�Q^K�G�4��(*/�+�,����Bgm�J,Z����+/�.v�%u�sM�n/�먺��X?�
:yȩ�;9p��@�	U����\˅u
s��1��CܭO<)�ү�����l���`��I"��J���&�G��zG��{���0�q�R������	s
�t�E,��u2rř��~��'.�^���3eaf=��0*��V��]��{��Q�%�#B,��V,����Z�v�gG�a�x�m>_������i�޴6F�rpw�����]���/�x�xpL�&ùF���Ař���oK���A�2M��[՗Lh���A���3�4$�\H%��1"�k</�L]��HZ+t�����y�[<���@�zYD\���8���� f+Q7o�:�<h��X�n�6f�#�V2R�sנ%?o�9�gּ���b!�
 V۠Ôk�VࢻFz��nY͏��_"O�p��f����< ċ�@��O��E�|�����U��1c�Oa�?'/mh�.`s_�\��Ee,�w�g����z����w|�fB���i���~��ax����R>��2&MQ��ƕ���+�ֻ�Rrrg7H�F���׎�y��E���lA��e�֜��2����Zq�#Da�(39j��[|;�S��l��P�(��w�Ǚ��R?]hՙԼ4r3�Kd�^�+KD�t�������r{�!��8����,���Hnj�ғ��h����� 3��Lŉ�w��H�3��~�`k��K��v߳��[���,{DZ/�$'ȴ��N7��}^�#++�H��E�~��#�K^�3���$�k�ʐ_�!��]�;<��L��W������;�&Х���Q"~&(Á�V%2���P�(�ϼ=�	s��n�>`�}�+����d~�M�䉌�.^�&N�T�a��l/�4U`-z�Êz�i��ZGy?�[���v��B.e�V�k��Gs����B9MpMF�l���	��{΍F+���Z���j���E��5��i����7��v������v�)���#a0�U�D飞�q5�
�K�T���$�`�U%5���}���j;�����i��T���6T��-�p��/A|������ǩ��-���=�jk�j򹏖[�ү:
b8�˓�
p��"�5q��|�^L���ȒLx����5��Cl��͊Q͑W�@CR�o�4#�4��_���
@r��* j��]���I@�o��C S}s�>zP�nYګ51Y<}(�_g��W[���I����'�����m+(C�㳟Nv�>��c�t�?e�7�(����{E`��&$88X���G��������eg�����O���[�w�,�B?1l�i�G���k�Je���h��w�`>	���Q�G�\�c�~#��9A�C���nf�@�0�\� ��g ɬC��J�#�ט,��8�@�Ӷ���q�i.eΫ�YVZ�������l��zɷDkԊY'&}!a�c�MCk�x�ƈf�"�x����-��n�yDp�ގ6�Pe����Qk��l�� �y�&��� bi�´$߶������?�`�7�\/((h�a3?Yi���Uy���)2�$P�}E:��=�eR/X#���N�4yo`}҂�\�{�@�;��@�tݩ�b�6�^�0���)⁇
{���29�&�ߧ:�F#(�Zp�vF�;5�h:*�Z��Cdmדm����W����r�G�85��ſ�G�%g�]�njڕ/q�l��,���E���� 4��1�8�:�ܖ���@
T3�,�qGR��ppp�^�z5؈��fy�y�.ԜY�1��{y�<��גr�d�S��3�X\j��hs�I��I�%`�ώu�0��}"Z`��aǀ�+}�ž:�����CǭtҮ���z����G`9j=�}��4��%!xZ�����Z�e�@v�+�s��G�i��JX₇f�LbEz����U�<ә^ON����7,�X�g��b7n� cD<Qd+ RW�%`[�M��1�kt�[�h���U��\mYƊ�yK��ˊ�bRy`�U��ܨ��%_�Lj�/E�����5Gr��ǈq1_v ��Y'k��Ϣ��K���ٕ�P�ﯭ���k
�R֧_Ϻ�Go�U�HIt�������N4f~�5Ln1��C�d�.C���:�GC�֧��w��#a�Y3�E��oM��(��Tʦ,���Leg�*]j(=�H� �N��^�o2�� JH�}[�ކ�lO�H8!����Lk{�®ɑߖ���U8U2tg�X���Ga�6���L��}�Y@��?N���ד�K�s!�vܰva˽t�9����ZcccWМ�Z�+��RӾE��, �NL|ÞT�����F ��ys֟<�S������K���o���L�- ���d������FKr����;8����{� ���m:��tz��{<!����=�]��L�e?�&�'��ʦ�OuW�ڍ$���:�E�쬰1O���B�����9z��Ծ�����ᝡ�� T��Axt��z;CØb�����_�\����6#�k��Y�������n�9<I����D��	���W;P���7&t�<����u��ta����-����Js��9Mk��GtIF�7$��~���h�B���Ǆz���-�M�e��~L����G�9E���,�b$��oN�~�@�)�ad� ɸ�.���[����T65��87� ��9[?@�TvL�>��nq38������h_,�����yKG����y��q"�a�Z��JW���G-�$�".B<�x���"��(�q�j�㗭��O��<��RL�;�;�.��lR4�ɥL�D6��5ioj��^V7(ћ����D�zO�3=����ui�-�7"L��}���s<ĳ���V��-,�����d���JJ ��}S����%cN���[��#�E��d��xd:��l��L�hs���oZ�a� Sߕ_���_N��_��n�!�Q#�D_���i�8�)��zޢ�r8�p7����4��o"P4����^��Ru�&뿹9R�ٴ�O�r4���-		�f�����k3,����l�!Z���(�)����w�w�?$��ɉ0������Q��b
)��?P)ּU�KJ�Cۗ4�0N�&����>=o��?�`��l�w��d�?�u��s����S�X��E�c�+R�%R/�R�7Z�R:��˫�'�����K�pk���Y��tU��C
i�
{! ���+ާ�ermpK�����E�����
GY9(HU�����2����+��t<�.��sɞ/ԟ�.g�����������9���"Nz�	�S�M��
�[��jA,�b��Ud-KR�V�q�y�̎)�n��`�U$x~�p^�\�=�?	���_ iFD(���2���{���#1}�k�~����m���s2V���c;U:us�P���B'Ɇ�@0���Ds�G7r�$h�8��%x���p�fW�E�R/�Rꜞ���+���i� �c��j*���h�I��a��ᚿ��I(1�3�%^m5��4%w�wt%��/�(�j��X�(x�ۤZ�?iM�/X;8�e�����J�I�I�**�3�ړ�|����S���z���g�l�N�fnO�InPQU�GZ�l�#YX� �4�!u�C@� �� � p����),FĄ��
2�暺���g������j�"}⋳c\2���s�뼻��Q��9ћ�7�7���0�J�Hơ���4�>��q��#n�9�*��+��B��!�'����[\F��q�m� �o}7(�J,[aC�_�ՙh��S���l˦ꪅ�,�	��$��,&g��j����[�:O���^t�.}���M�M��հ8�%b�7/ۯ����^�u,r� ���X�8|r�	�pߑD�7��p�Y�+F-ᅏ'y�ϭ)@���5��xNB�ۮ�R�˂D��E|���}�F�!?�jG n:ռt2���CkV����KM�N���x�,Q�y ,f `��:�v+$����.��uz�^ۀ��b���*�
����E��!}��/���b�觺@�h�͈�7	X�d0��w	A����}vT�IE�UR�"ؓ�	�#)M7�h��>s�Ya<���]�w0wi�fp�.�fׂ��?�ym���o׌��=e���t��'U���Յ��n���2�D��������M�eO�X.'�m��'�H�nqG�t�0�����վ<��I�f;#i6)k����s?�	H������|����WdA��1)n�h�v��X�N1�|������TTqޞЅp$��������T�B?i.q�""�?*�s���!� ���`lM�M�}�7:w2��h�ˤ�&����s����C�;���I�@��c��A�_ʖ6U)��rE�5�l��!ݎGB���P�����R���?l�AS	���M5E
�V�fң9�A�G� ~f������o�il�	��ʬ`�sf�w+ �w�F�F�w~�B���E��4��~(���<�,�_$���Q�#@.s�9�p��TUU�o��M�V��&��D��i�9��hLf�x��r���N�>��K9���_��߿HĹwGA�]=��F��R��?K�{��Wy!%3�����Sf�C*��vwzu0�S��KG��Xh)5O^j]	7%�q��j���C��A�X�H���x�߮u�o3K�z.�=h'�����B��POe �80�S(PE��d\�E����
2U��3s��w[�E����hN"�f?Ju�jn�XTvv&�gސ���P�Zn��S���g���I���=g��;�������eNo�?�6Nx������6g��/��4�K���pU����A��~G�"�9�#��e�1�Q}�����$>���o&��M�>��O��K���n�gw̷'�1��-Z���@�r	˩�:w�g��nt`�hv�^�Q�\2� M�!zfV�\�J)YK��*���FH����_W��c�5y���Ǻ�O�k��o��0����}�|la��4r��NtLG?m	IT2��ܻ̽7s��kt8]�1��P@YlC����h,I�ƻ���z�3��>z)Xo�n&:u�;"9�����������iGN���D��G�J���
C�͜pe��i�a9��D2`��+8�k���e�ECV�W=�TѓXՁ!�����?ֽi[ZZ&y,�?�gKz��9�U�)�3��?���3����b���֭��{�lzr o��À�ȵ��Er��B�*oء<�0���~����b�Ԓsq6鲛�We0����f�"J.�	.έZ�*�[V㠛�8,�t����n�V�ρ���`\��E��>��ֳ�FJ�}ܨ����}R	���݂ՏZ$1&Wx&�D3�G�ٚ�O�}/�u�o~�3�％�,��.D��: �e9�g���&X��s�&��WyϬ��t��4L�q��޿�ߵ"G���v�<W���.u}/�������������oT#{��M�z5P:�n|'	"9����?���8F�8�����tv"�ZM3��\������a������%	u�R�6)-��2�[^X�a�f������A�:s,��S�[��lG����k���Dq;��,xRSyf�Q�����C�n��p���?��H�):��<9� &�I�J�1��@���Y©F�"��H��}��Π��Q���B��]q�Ӑȕ�XJ%�Ӽ�T���ت��=-��EȔxd8>x��|뗦ο�qބ/Lu�pr_w��utG̻��пO�q7m��%k�فxTr~~���}������P���q&־[R�g�>m��ێ���_��-tZ��WԢ�LP�ԗ����h6_�����^j�k'S����s�"��<k/�/l�M��*��l�.0Uj>�0ѳ^���:���
i�AÄ���(�nY��]�'x{P zȻ�|t�ΰ�#�5b-f>DF�e���ʑb�eaq�y+���u{6��W�U�N�S�{x���eJ������ĨKJF-�:���r�N
�I�U;(����Vm����"H�U�̲J�ߍ��U��z��H�*�½����h�.��#Ű�^�����V�|�N۔�/�R_��yEY�h=���P��;nG���N�����E���Kf�_\\_�&����~"f��-#i���=�}||`�Hx�����,xlL��n*��b�}h?i��ť��J9w~N�y~2-x����m=��������K&r�a�m�3\��E����!�fFlt��T$���!�c����l�$s"����T,.2v��T�+,��Bt�l����Uخ�*�yA�S����6h�!݆c6:��N����T�8~qR���s�X /�ֿ^'#�8F1�b�]�B%���sጉ5p��Ǜ-�������W2x����l�	�Bf�&w���M+����r����f�'Ϳ��Y�<���Z�/������y�=\mއ��:3��C-,�k{��0�dy�&ؽ�W�l��M��dXu�?s�|UY+�~�F�pA~CX^d�d��?�i|�q2ƒ�K�ڰ�0��pMScC?{I)�a�ӵ�T� ��m�x��O��gϨ����y4�+-ⒻL]�t�#�f��7�k��w^��Z|
�Z�e�ծ=j�c�a>Ԏ9�錡� n�����:Nen.�4ĞP�%p~�e�Ap��rq�nY���C}�m���;o�Aź��tǙA�Dv.�����D�\�^R������z!�`2�M�tL��q�,���:����䧏?a�Nnd��V�w��
���/ �;��J�z��I���(�鉏&����{�)bB�5�����2�֑�6p�oS�4�H@�y�
�B��L���yOu�����
pjո�![Z��7�\�T�c��h1�ؔ�e:&LYj��dp� c�i��G�6�qMn�-�V��!��;�@LĠ���t��gC �Q���Џ�dl5�����N�E�Y[6�fX��3|��,�W/�[�y�W�����0{�æ�?f��T���������A���� �E�+�r\�j�U)���Лɔ�w�
��S<]�M�جM��t�{
s5_��b�VW �݉,ǳ���*�@ "���\�� ���	��FF5k�q{�p)th���>���&���p%l2V'�Z�9/��>���p���Gڣo��W2��3�2|����us�j�"m<;��⭄��.ڟ�`0Ե�uF��E>O���YK0�M�u��a�-,���c�^^+^	�C��w}z���q���gk�`�X�|��]�K{&|]�F�$%0�S��t�+�����[��rZ^)�������ۥ���'+m7w���1�>�εV_��S���>��z��;�7v_�g�����V�m&Hg)d_�3��wi�==�1����������;[�"��k?)�j���Ύ�ׄ7ՙ(Ů�y��/�RBa1��]��6f���XJɨ���S��h59D�Jʨq䃌*R�VzH ��-��Ր��iJ�tr�s��:˲��r���(D~�>�e�I���Jq�]��l�_�����6_ z{㜃T��K"��{��5�W=�7�nP$T�sB"���U�l�%^��(�2�hTv����c�%7��[�����lEbh�B���XV�K@����[''ޙ
�9��%�����5)�r#�Q!avɗ[�/Õ��;�p�W�&��O>���8�l|%�wk�.��[�V��}8�ɉ��h�?ο�n̝p!��Y�9��8�­�^�F��#�`��ϪDI�����v��P�#��J����G8�_�-A�K����q�@X�D�����f��,��<��H^��gwj5��\&�uC�y�8�Ȟ�yB���\�ׁ�`Y�+���,S�v�{�:�FZYE��e��Ï�\DH�<:����d|��7'�?�����ʂ`]ht��3�̽M�ӝ�Jd{�1i���X������;���^3���q�Iݼ��-VoJ���ʺYڕ�	XG#��0jB��{J�`@/�f�.����4t��M:�R�ŃqT���i�EI���r�ܾ���6`j�D+@º�b9븶�x�4�0�i
p�5�bv���Q#6r�Uh�Bx���O:lp0�m�-XS~Ȟ���ʹ�/�s0g�&��~H�a���Gq�zh3<��X��N��^�̯]���k����H�O#,{�\b�dہ|�S�@������j����~�����W�_�\��9r���v�=����������94�i72��/]���i;����t��r��w��M��R� �E|`�V(���8�x	Ε�f!d��VQ�f����a6�d�)7%�\j[���TH{Z����7}`��k�k��p���]�Y�w�6��������0����=*���o
lC�T���'��"\Kw��O��}�S{+_Q�L���˲>����� 1Wm0���h�I�9]��K�zv�
3��3
�Tx����\�5w]V�:}�Q����[�߹���="j��v��)�8ߖ�W\���X
p>p��h�0�ZG����x]��-)1.++������:��F[[[ ���=��y���Vy׵����O�v?�@R=�Pu�;*���5S��`��B�B�/V��O��QuM��ݰaʎ�۫��Y5Ĉ^(0�hm�<&6Q쟎_�z��G�yb�.�-H]?��wZZd���ű߹��@�=�zu�T��HCҕ!o��80�����4�Ѫy�*dDk)���_�\��f��GՎ R��R�}�kY����`�s�=�3K�(;�;�IEs�x��Ip�l�޲M�����2�̯q�X��'*��22�Hy��*����� '�[P�3F���4�a�.�������G���Vђ 2�6�L�4I_�1�g������w�x����]/G��1�_M�lD����A�!X.S�4i�$���o�lÓ(���~
ϩ�n�!�T��n&�C;�3&��8�q�7c��J'J��f�C���*���'�(�r(��֙h�����l�T��Y��a�,�m�jm�������=�K���-{L���3�r�^�ʀ��+��M1n��>fc�?�F�m�?�v�zHҦ�:G�H��G5��w%�JFOV���&��e{�$:�NbU����w?i��h�������0Zd����q;6� ��IE��բ�SC~4��X����Ug�@�.]�&r���):��@h��|\���r�FQ� ��ۀA:;��
	
o����m&i�G��5��Y;K8��W c6����'
:{�jd*�+�.�H���6'�h�,�p����z�|���R�@�7tc��P6o�qGA���U�A$��!}�J~�
��Z_��ob�Z�C�߮Rc�<Ē9s)AWs���Gr��ީ7��ZO��'���,��þ���̓[�J�sH��z����=7���^���V�k,|,�7xv �����!���D���T�
�?�VI ��m�V{_��yu*PT'���lI�B��>�	��v�/7c�vK�"���P;W�6֠������cY+++[���K�K.�,�f��"�-�Y���1Y��6��P��,N��<X]U�^�&(V�C��O��e�u��Vz��ă6���&f�Ku���_�m1��.�2�CEt[r����T�A�H\�Dڿ9�����?0�+k�cP����_D��� �H�" �!�!"]ҹ"���"-% ��� ��H	,]K�ұ������=�[�qv�3󝙏�sw-mW�=��|jG�O���V���¿��ZN�ۦ�=�=��[�۬��!K���	�������t<A�o���XX�;"wKn 1�7�	]�k�=2%w?�P	z[�6/�-[�A�e�l������'x(�	W�S1�~���~Ǒ��_���	��-Dh#�I=�,P��ڝ���M ���K��#��b�����sB΅)P��5�����E�1 �%���<n!��2�,�q�c9��W	zV$k+=D�ݨ���E���-6��'״�y_-7��ꏐ��fu}qu:����1=`c�U[��8�Rַ���֩�ǒ��s��.���u�-��X��D�}�7�kq{��4�^/& �R:}�
���U8�?�*�dE>�������!WϞ��� uTT��X��nA!�s��);���\=Ǥ*~�T�����;�I~`I�?>�]/_�!@��~?(vzl��`t��0�� ����d�f��er����w�36�-��A�����'�����G��91��D��!a��DX�S�xZ�vu{V�VZ4�n�|�{�1�K�[�7#�#!�
-R��P�j��ɾW%@A�c�J�W�п���@ѻ<�%�%���G�R�O~��o�+�نw���?\�)&]�x���Er�8��TF�)�2j���kk��0	Ǔ@ Ժ 5BJ�[�ѿ�����toUh������u�?y�lQ�b�!��es��q��]bo.p�xA��;f�Qj�Nɥ���i�z�)��R��1,�"d��؉3/�_���#�����!߸q[z�6Um0�m<�Z�2�?f_D[�߈�+���_�d>U�6��	��� Z��Y{¨n����9.	�����o��t�~�C�q���i�W�ITǻ&��8�uDA��e�?�,|�?�4j/��3v]����t�,K���D�ReX��a�����Oнkm�SnsK)y���J�T,$�Fٶ4�ԝ��g��5�܈�'��oؗ��Թ��H�
)�,}��S� 𥆮iD��2)������?anm&`� )�8���4�����ᘜITG�Ɯ�q�O,��B�����"ވ���e��S�[*�R[��GٰN�OgO�F�X�G�iFP�۪�z�c>�V��o��D���&LV����
-n���L���ֱa�lKa�2
{��%�����NMX}q�?��f 1��O��f�hV �ɧu�%�'餹2ǃ5���MıCؽk	=2hX8�G�j7�1��k�(|iF=Z�7ĥ�w�������Ės^E~���!��h��X�� ��q�ښ^�^��� oSv�r8���r�i�F�jKH!�t}�]gt������13䵃��n�񃛋�xz ����p�@ą����k$t�����v6������/�g�j�W�����+ou���@!�GK𛼺2��Q�>[�i�%�)�,jN7x�:���������!�>��໮�Eѕ7X8�T�%�\w�1o�ϸ�=����e|_'J:�j��+M��6?c��#��8�֭g���;�aC5�m]�� y_����C�%����ɞLt�Wz�tB��s�ns�|g�W�;f�2~�jS��o�3�F�3�-p���>����a����ك�T��.�N�) _��w΅��Dޕi�����m�*}?i8/+cY�ZʡX�qt�%�؉�/~����� ��������)r�ga���A̳�y-b�������&r��u�+�`_y���w�h�hp�[咽<L~�w4BK+s$��4�"Y]�ݱ�Գ�����a��/��Xpvљ�:+ٖ��Ðǌ�°�V�[��"�f�"ӛ [�ٲ�����>߲���?þ�X�?u�F�/��i�^���ȠԮ1����T6_$Lu����)�[���x/,w�&��tU�kr�[B�NR��i)�h����zW34^�s�[{�ġ�T�y���k��?� ��e�����jA������z�����o�b�Lt�6��C������j��S��:�g�V!�@�5/Ft��ܝje6/��!Q\�=��a'���h�#6]����"^7ƛ''1n��5�V�0��y��u�r�N,�Hv��mP�H�Rt4�.���&�`9ۛ_�*Û"�پ��c~��0ؑ)��|�2�DD�U���B@D[����E�y�M��R�-	�=��ÄǓ��6�TV��r
xT�7���2h�x������;!�<r_�e�7�CL�|��'��H虈K4V̏�E��wW�]M��eS���n������r��؋�so�f������5�H$�æ�#YMsK�CS���Ck�`J'�y�_荊��o#��T��z`]�lj!��Թf��1�W��9Y��&��l��,�
��$���((��q����y��
"��u��zH�[ޠW,#t��0!�D���c:\�P-��-UԬg�����ej)�o�Ι~�ER���s����oʢ�������%�6kf�ڣC
���1#r񻭈ms�����)[�[Ǫp���CK�n�[@�k����x�h��T�p��S�Vя+�B}\~�ѕq�<�v�3���Hk��������p���<d�d��[�~$�V(-��Ȟ
�l���{��%8?����Σ��W�pd��K��:��\��:�Hom�߯��1Y}�.S�҉�?�?%-;fg�8Hf^wf���Q&4iٮ�s)ϴ���Vyo��r%��Ā�ILǬ�{٫܊@��������W�&��|��Z�R������טQ���+�0�4�����[7;vg7�3>�1�� h���j�m=��1�5�R��h��}Q�&�a� � ��D$�j�w��� ͨt��L��W@�Xؾ|�����1���W�� '9�����tc;ZHX�kz��X~��',M	裳�H| Ј��M\;����lV���N��,E&քw.1��r�ҫi8�Cr�95q4V�����V��Zn�3g�k�iV�FL��q������˽:��>����4*M��o�����E-3���hR鹖��5&�fD�0CG~d��֣��"_��[�&�E�w֒�Y��SN"��|�!��;)���y��D�b蒡U^�	 n�R�5��Pc�@��:^��c�ZQ웣n��Yէ�+��J��+ɓǎ�Z1SK������1���\>���5o�7��?-<�\�'�pmU���᭦*z��ΙE4[�c伩��E�����ak[��O�m�/'��tXǪ蹭zY+�}Pȋ�q$oe#����^Ѩx)w}Ѡ�ӂb�e��H "��i�ɋi��T��KO�Z�'��q����G�5VY6<��K֌�a��ͳ��iՒ�C�^�ȱ��w�c	��9p���S~�~���l,�He�wf#����b��'���+eR�j�S ��L7`;��ųU1��z�*�O��'J�a_D���K�	I`v�0wDG����H������pSw:�!mʦN�#�o"UÎ�EV��;����KOJHטu�^2����0/��t�>k}U6���(,��/T�l����W�Iq��~X�ϗZ>�N:>1�h��1M��g����&.�jA"I�T����(����W��y�.�e�Y�-�Mx9�iDt��%H7+#* .Ir3q4 �� �̲0|}�#��A�L��y�m�MG�Y���Ij���p���>!�F�V��r�[�(;M��]� �	4@�[c��⦧��)l4Ĳ@CR.X���qRׁ
 �4I��RFu#��fL7��|gwML�v6�h\���f���W��&�6�x2ޭT.N��\(���Az���,>"�����K��~���E�����/�T��������l{�I�	�@��//Ɵ�ހ�c֝������X����1������Xä�L](c���Hu�1�0 ��Q���6�����cx/�C;|�k��yv=�)
���iS�]�~����+�墥��9�J�&x��a�h/$*U�I�>�D7�����P}�x�|8�W��a$���<Q�ٌ��[P�?�G���xC�a&�޾�ɛy��� E��5�=}G[�Ւ�"�u�^�=}!y�?Yq{��)�̅�~t��1��4���Jr5�;?�f��a?t��ܐhd�w5�����!���Y0n+OЖ`k���NCմ�3s4$�A|BL/Z?�xYj�;�Ր�W]hc*q*ݳ� ��C(�����m��0ʵ�-w��/������SE)�\/o�2�$�q�S�ֵ���O�����F��^+l�Y��*�6 '���#1[#?����5����U
W�ߜ)K��)#��^_�Dа�kJwO��
ҭ��-z�7V*�����3�
֠�H��#o���L���n�@��l�����Z��A>_s��>��9��!�a9�c�ޯ����A�I �]CG�%�!.�5���	BoB;�R�c�g-瓪���獪�nD�H�Ǒ�� ��X�6��,���*O:���ps嵙����5�~jN���z��;�O#:��B�=�|�g{��P�.��%���{4o��T��za?r��$H��jCs֊�G�=���Ā�'�V>��E8�P�q+8y�:��@�뵞#�X�^�~��1�m��4)���J��q�� ��M����S�^�,�döe#P�8g�dO~�	�F��G۔5��\I|6�e�� �f��hzL��2t�wja�׹ҳ��n��[PL�$@�d�����W����e��ng��|��7w��Ҿ�y+�����h�=��AN4����C�;;;�:֢i�gg��4p<B�M/1>j�Ư*�9�p�6y�Q$��-�\Qʬ�bl������浌��2oIk�CU��$费��6y�^�H��P���=Nm/�cS���<i~�ν����,��2�'��%lm����j��E�ל���m��+�9��'���v�D�<wN��W�M�U2y���O� ��?[��*%��ӭ�����^`���;��x�/3ц
�3�eEy�o�500�ɓy��!�r5��/p��NV���4�z	U�xߚ���w4p&8ۡ/��d�*�v�C������>�l�ݚQ�^��y�N����Tr|;??_�P���?�s]�P������R��l$������kX���>al��_K�W]��`�/����h.7���S�8��\�F��!�}0��2�i>oC��1���Fs��w��u)��*��&)>o�П�׃]x�����?
��v�x���!,�AUq��m�ZQ~��L��g��\'h�b�e�/	k:�G����[�'�ƈK�����)�7�{�w��&6�3�4��M�?A�'#"y��'$lt���
-�fꚌ�.�ӊ��� �S���9�^4� o��[���؁��0��#�ڒ��{�!n�R�$��1�)�)l���!7-�69IqZ��:�VVR/��������)
J+~9G����9[e�4OI��s����l�Ih�tP���RF桎�ϔ\�g���^`����d�Cȃ��bmnޮ��Gn��qk2��D�Rh!�fZU���-|2�o@�q��t/I�Z]�8��
v��ŭ7P�h�����K�2�W��8S*��7��+*��rS�k�̻�5�'S���f1:�"���d�5z�}�ӫN����$�W{��ƼK�J�s̮�o���b�eBmK9�~HR�t<�׸/�NŎ=20��f�FqAD����X����=�<�T�]���/Y������{�q[����&&$����4����LƄ-��$�kD99X�^N�?^���R�OlR%�u���3�J���7��s3+'\J�6�f�n��.$�Ev�Ŀi]3�l+5���Yd�.�򧴷�(˼�C�Q����� ��z�B���8]�Q��0�Q�������6D�I/XC��X�v�_Xg�m�nJ�5Y���+�K��܆FЖ|aE�w֑R�@��*�m�KFx��t�E�:EQn�x�V�=E&�|�B����M��p���o�_���/�Y\��+&�O%21=����bY}�nk#O2���"���<ޯؾ�0?_�4W>��2��0p_�}��0������ā�U,��o����1�r)�a��s	�8���D�c���F�n_��ژ���
�✪i�%Ne��u���K�0Q���ʤ�\_#�'q�u$�c'�֤��&ӥ~&����v��0�*�����n��H9���g�:�g��pv�[e�O^�Ps���޹��OH��k��v'����߼(A����~Z��z�ş���6�����ʳ!�0wn�b	Km�ڑ�k�G������.|Q��qG���׎u�?��\�	�-aa(UF,yP3_��-ď��>3NhI�f�<��|_Q/������Ў�S^�W�ƆX��!9�=������K�C��h
�c�Tʸ�/+
ό���;Q����Ճ�MQ@���ۍac�s�ؐw̘�"σ(�#�d���\�Z��쒺y�?L��kG�_Zd�&�N6�pt��R����W奋.�扷��<�
:,k��(�����\{���N��ެ�|wݰt
�YȯSh�Å�~t�6�aybA�.2��G��<M�.WC\	[��v��dN�K%�#�p8j���yc5�<�÷��e�����!�3��*����ӕYK��Ye�rX�^�懻$��'d\���._���x�f�P|.+4� ��j7�̍ʮ�������n���q�Bv~TA+.f��?&��B��h����������
c�>)(˕�I-l���8&�a��'ς��6�g�J�*x�<�(�������4�~�3�o��^�D��d������<��G��1i����p,�������I֏S����	G���k7���K�����t�wA�v�����ʇ��G��Їųj�&��i���	���v��@OB��3+�[��'��9VG�Oc%�j���A8�8����~�F|?�<���
?��$�(���<�"��:����3�(ݖ�S\�!�T����݈�P&V��^�Mw7�8>��"����io�n�H��k�]�����Sܚ">kf�pdGKv-�'���n��-��]�w�M�21��M=~�HF`�S���!�Iz�!׫�{F������0��0���'[���aG�7�y���ӳ��k˕�K�OŃe<Y����[x���Q�1�kY�f��N�zn��4��=X�0�S�F�)��g������I��uD����hݥ���Y��b��=WI�B��oJ�ZL�:B�1�(l�C�O�3�������JRDw�F�7o�|@��B�2� '���1Zb"򽲿)�A:���9-��ەK��=h������+˒9��P`��o�����8��]?O�p��H��o�����F;GԆ���2Y����ݣLtNoE�Xa�N^SBF�?��G�U#��3��X����߹�b���w饒s��e�˒x�!�yv9z�7Fm5����Њ��Y��4���Z��ȷ�0�_���*2	tU����(�ڹ
[�^IrB	�v�����La���.���O2�j��5Dկ�d7�n�z���(�L@O�O�_Z"�f�㒸���_�QMIS����)�V�͵���o" �����Z	�Q�V�b���[r%Ha�|n��{��;.�U�9׮�i�A���J�4"��/��G���p���vhBXʃEzr->�P�Ah�y�^�)��Ũ�Wu�P���bE�ҕ=����U���X��80qߺ]�W�e�5����-�5�ţ�hDX2]���$�=�o���E���(�>�,|��W�A;��:+;a�V@���8:ʧ�<�Q��A����F{K❗u^!�H� y���������b���q�1ek&�Q܃���:�MmP�(��HpXGB4؛�ζ�����+�XXLO�'�_���
��{��*�\���I�G��$��\Q�K<5�0t�,�:�/@�ar�C�}��q���37","��T�8����x$����T{;���X��3���E���~�6����n4�b;��r�×�6����ζ��"-�3$K=3��$;�`�:��d�L��U��b� 4����!��rl�O@6#k�/��tz��ǌ��^����b��������Mw>�J����&f�CT1�"�u�s ;�8�tPo�.����!�W�a#1Cd�[^nn����SX���'�\^��~��N�T��?O�������T@m�x �53R���<��K!���fkä����{>�Ψaˮ�h�>���J������΅{¬W���tiS����{撶���d#��E��7��V_��E����ް�X�|b���|����f�lj"��U����]]�U�IF^1h`t�F1���ZM�e!�Ipԟ�k��6B硎�!�@��̧:&�crJ��i8��1��L ���^o�]���r>;�^����%��N�2�b��D��*Sf��m2�_I�؏�����N�ŗ`(*�GI��/X���ׅ�7K�*&�w�]:��he��!<����)��\�d�/iLq�~�I�o�>jc���wx��agyZ,�b�x���{A�p(��xu�d``0_**�[��Y�D��������d����.���_���S�+�@��	x�=q0#�"}+mݘx )��J�BQ�H$�����Bk�D�`�����D����VBgA�mv'x�r��3Br~@����~��f*0jw?q��桢�S�:zx�@h�s<����j��&���� '��c:x6(�ABT�4��)��0�,�Uh�~�V������_��em�KJS��\&A�վ������?�V}2Ƭ�7i����6+]��W��*)�D�JϺwa��׵'�}bh��W�����a�sZ�Qgռ}��mo�Z�|��l�s�3�K"?�@"G��!H�d'�/.c�g-��/�)�[f��#d�EE	`�ܻ�x+r��������<d��Q�;1Nq�_�7P6Lx���\�0�|�+�GO��O�W�`d��Y���@#� LS]�,v�����b�t��9�IZ��|��� �v�J��	����b���ox?@�v��:u[?�men4Pa��wٺ�A�~(h�6ۙ�����N���
�`V��r%2���Lf1]��)y?Gx��}�DPn@�=�5�֣���gh�r�dBO�+��@	��=Dnd���GAJ�gK̆B����3�{rm'y�zz��a��/;�vfv5|,���Yy���m�)R\S���Ǘ(�@�>�GѴ�d./�K���/�$S=�؀����a"b�?D�$��+R��A\�7n�ϱ~��^�q��?W
�Jt�Kd�&T�a't\����X�f���Y��s��odH�+��l��@&�r���x�	�:�E&�#�����f[�:$�4Cw�ܚ�����:�[�J:hM��O%��?H<~ם`���VBk�OX,�Q(Zwd��0����|B,��D_�K�u2��._̶l�<9MMB��{oS���'��7�&�H��܎w�>Y�r����L�__�����/�>C�!��a�?>iY}�F�3�>�w�i�o�-��I1�RC ��,gI���� |��(:x��?��	��=be���y����,AY7:�sغ�x�	�H��ژ��w%w���o���r������v��ں�<*�d�/����s[��|�4^g��`+��Q������S���.���l]yW96	�b�Ǖ����!��}���<�^����|����h~��8����}
pbb��&�ևԑ�9K~���j8�-Ol^g����B��Tq��H��uzn���Q��2A�,qF��`2?�	_�bn]N�c
����N�)�JP��2B&��eE�~N_�¸���g�T� ��d]\[l8-jTe��:d��i���PXGX���|��h��|��G=O��xf������[-�I�/	�4��;z9OW�˽��P/�=��t4	K���'ȲH1ݦ�`H�����h7�����_��VO����_fI,I���]��MK�.����Q"+A$�k+���I�~+�>�#�J+�@R��SyL��jj}�nv4@�c;"�\Ph����'�XeO�e�?<t�w��ߙ�K�MW^
M�ѯ|WZ��|FK#�g��kd��;gҵ�+DYik1[<��&�U<�X�J �2�K�3s""!���X��:�g�ځ��PS`�ؖ�硧F>�>h���5���/��_m�<&�Z��q_��6�`���J�䯡�Oh'��or-�'��y�:P��7#�g�$�'��z ;��'���=Y�*����ܴ�yP{��a�Y����vi^�:$k�x�u&�^\ u��U�d�&O�GvEy20�|Ur��Q�?lЗ���o���G�z�-qS�GL͚+(�$?u�f��܌I4vK/�a6󩈔��{���,N��.]m�l�W��b��$/*5�����؁U��K>4y����΋����[�����f�-9��6>���V6�f��_(��J��,�
�zwh7H̾nhz}���QZ��%��2�[��*\ĿQ�n�@"!c��ⓑ!U��ee �>Z��t���I��7)����V��׽S;��صQ��p�v+ʁ[�3���9�{>��y����M���=[+���V�'Jl?
*��M%̆P����H
K���((�~����<����8��d]�i�4�X�Q��\�A���C'�m
{�(�'W|��j�M������pG�	v<��u>KM	�P��',��oɐD����1�A��	��HT�>Mm9���x�����	陋��1����7���Z�j�8��Ua��?�����h\ 7M8»�����ڱ�X�2@0�=|�u�#:}N��#�n6�Po�:\:.��
\�qX$����L�����݁�q!#ugR��q���9���b��G MȀ�D���n���ੑ���t��z���з�K�y$��T��[��dR^��4��	�{G+�5VT�ku��k�T�ReĆ�!��Բ��ʓ?7���OB{���Ax������wt��a�$������ ��*�ܟ(�ٯW�\�C�!W�����`�ۮ㮻�����2q�1���NQW9k*'�&u�����\CŎ��Z щ��-ߪv9+�����a~��˲�uÞ��+�w�+��S��<�/?�b��g�TJ�H�[xK&�o1����)���x'.��I�\��k�kl� ���h�Ê�Q��V�E��ւ�BdH�h?�M�D-2�nqNƗ�C.��i���� ��:1�g?d�l�M&:������3����^�c�|Pa�mH@9��h_�e���=hO�С=��ى������%����1Ĺy�׌=rT�'p�μcWݵ7Fa�SMZ��םD�|���">�=�0������c	�R�-�T��Kn����S�t)�p�;�f@ Z]=p!�v/�a�)�[`B�{�d�0�w�[��[1R�o��'�'�d<R�+��@�~��iOe:S��a���(���*%1�FJ(ߤ���~����	k%Q5�-C40x��cT�Tx/q�pw�X:��fE���z�?�Օۺ�x�S�a��{�=aT���P�L_B�ˆ�E�an��pP��&1�lW3��&�n���������ߘҟ�%׉�_I���}��FN�z.��j�C@�����������A��:�z�㈃cV%�7��e�F^����^	�ZR�*|к�e�g�WÜ�1��Z�Å��+���& "��y�v�X�(^��:ڝ�*�v�����ʣhʮ�nt!Ao�F@�F��O��S�+Y+��ػi�1��_����V0:̒����'Ԭ��$�'M��`<�_Rd�S�ym��mL�iR�Ud�R%/^~�5�<Wܼx��i,m���C�h^�~��9�&Y��?��!�]� ''�'�XK,&�	�=��$`���^�F�t���=ޭ�wl�L�D�]�t�9��osu|�f'�#�Z�}	�i����l��#��ٙ���Ϣ�B�f����m;q*Y���aM9�*���S5�2�_�W�-3�?���.>����B�E�C�,~�|D�md�ڔmhR!���������")����]jM��L��%@��(
ſ�����d���TӋ
�����UO�8�	2ݘ��;�2^�-eY�J�WJ�U���6G˓�T��S�+`�Gx�J�D��SX�ZدF��
(���}Ʊ'x����9hG����a�v]�؟�I{b�cN:�e�KW΍�r��YlP��V����-���R��x�V���g�m��g�˺. �LC����'�1P��4j��Ax���$��������SӉ�ϕ��;ʾ�%m��:	o�)����B��������u�n�CӝrA�������LH�~ʴ��4}yM�p]��Á�"�tS��1��6@�V���ۯF��W9yh�ʯ�Gz�v_a��3+4�zu#f����q�g�o&�;����:�l�Xz��x�����~{n���C�G���A�|�.��ڭ�/5����R��)��$"]"�fŸ?�y��庮l�);~�g��b�.Q�St=_���&�O�B~��SD*ae�E-��z��G��L"�ymC�Z)��a��Jm�Vy��\b�ѯ?�1�M{�{ϑ�E|�HK�{�"���\�����KH�����]u[�jרC c
�.1C�WX,�K��t�gB�}}��Wo�G�i|�
ݓ�X"�F���hvV��A�(�9 �L�#�\]���G���#OQ��W�}��A�{ �/�8h��p����`���Y��j��h�����c�j�m���p��SA��X�����a�q����l�ʲ��?��Ћv�ҙi>ȬJ�|`Gg�����:`=?�+<=`ѓ{���4KV��3�W:���dL�k��,jR��3i�LQ���Ӹۃ�`_&+�D�w���~�ڿbYW/�4���T��´R�e����- �<�o'��Eo�~\6�j~��K�:����YxBᗜ𩬥�;�l�ҕn�ƚg�-O��d�F���T�ŹXt���\�C�L/��^ltAj����
-gE���J�u�v�����[oL�p��8��Z���;eP�:W�͚����}�0������$I����3>���8��4�y�{P<+?�p|"l;½	D���� E�s|D�u�?��W�lU��x�ט=�K 06d�6�$���E	��O�(]$�V��w����D��板%�j��B����طv��z���痣a����\���p�$�{S�a
�^�f '�j�qX�>-4$6%��K���g��
ؿ����.5����
Y�<p�� f��>j��K)��N�����Zu�鮊L:)�}2\e:����"�Hx�
�Oz�1�K��n�	ZP�g� ����f�v̺�?����L.�}��`�&����©�*����i��$����߰Z*�)e���НZ<��r7���h� v=��g���_�˓�����$
��:nҩ��H�NK��C�9?Q�,��f:��c�,�� ��OBQ�5\GVh}�ܳ��e¤���n�f�F��J��
�@CA#�:j�"g.���m��X�p�#Љ�3� ��F5 ������������%�oG�E�^��&�!!���-���I c����7[���~V��&�Uړ*�JQh�T?�8L���}�kJVK�O�n��gM��%�u��$5f���i�a�9���t���l��wG̣����%�f��5�$�(�����g��f��N�~l�E�.����� ~cfy�52V�y��'1v/���_\�~-����Έ'�#)�)YR�����7��o�j���s�q�(�J� ����$-k>�8��Fak��mR�?p:{A$�A
t/"��a�5U��s�;-ʡ]��S�A��H��zy:w�ې7���&�a~���V}1�|W��Owl%����؟Mvb���b�3�X���A��\���ǔ^��%�<����(?�!�k�r���4��v�뀰b�Qm��ok3}ۺ�s��D4�^?��
\�u�D�^�a��Ѡ��'Q�G>ܤQ$,s���5�����=�=�1��}=o�%3N��oCy�M--쬀B
�G}��0�%�\ω�Yom�ٽ��m#��8�����������%v�ի0���iQ>Rg��J��vQ�X�����+J��UȖ��Z�oUf ɥ�$2�o-�U7�6�4� GZ�q��ʐ�[y�"It���I����
�Z�ͼ�<~�R�=�B���*��y�ɝݷ�w��K��3��,�`5�����0����(�u��J��Zjp�k�!���<W��_���1#Q=����t���˛�'y�l�n�a���7��b�͊f��̈́ٗ���]�/;�����%� ���$�N��V�'y�R<"�������f�'.���8�����ê�FW0Q-�Q�6���G|R�F��u�z�7���!�1�M)���F%}�z�W<bS��W~�G��y{�K
��)��#}�j�s�|�j�""����S*]=y���\%��f�!��B�сiVO�j�>[(� �4?��t�j�����A��� nPR,��HF����~I�O��uF���2��^-��l���^�s�ŧ6��	 �7��o+5�s�x����<7d�D,̶�^ׇ�� �ϔn�JnlN��e�7��a��^V-�M� c��r0�L�p�i��:[�$�Ч5��""x�0�Nc���m喫��*A�Z���'���������~�� �P����)�;䓄��{�R��i=���n�k�7C��`@'����8��X���;z�̻Tn2ei�Si�+�4�y�o"����+ڇ?d�|�b�v~�$��-��Fݯ �����N�;��h���,=	%�G���s��1�{�M��s}��ΧZAV��m��;x���l$a�D	w�h�B���50��o�Bo���ҙZ��� [��~�y��h������S)�<�^��9�C�SE#��OP��(�}���b�q\��a������j�{�]�=SI��ajM�W�}M�@�uƾ������_�5��t���p��(���ϩ=I�����o�fo����\��Xչ�<!ݐ�&8M�v䨐K�d[�!�Q��W.��O��OT�w��wv �St�V<@�Ӓw�n�E�x�S�� �P0#�9�q�GX�Y��B焷c�4T�����6��)ah�j�l{�}�ջy�Qo�T�k�'�h&�A��bI�f�;G~m��4l���et_��� i������2��,��������p�9I:Ŵ�O�f�����4%�I,�9��6�Z0Mu��"Lu�w�.'�Oi�a���W��XT�2t��,�*A.߂ǐ&���	a�B�/�݋���*p����.#�6��ʛ]$_������tm��+�K����ª���t&K�-ʃyr_}�nDB���_�G��s�+<e�	k/�5��֣a�������k[f�j@��
��:Qƌj���{�ݹ��H2�����~JD�b@S�c���~�uwԤ!׿vVv��ڎ�М�@�	}k,�����3+���Jj�1�9��&|@������A����W��.q��3�<)"� ���"vHo�t�LSA]Z�HS�zF�2�'�a=�՟Ĝ�҃�)�چÏHw5C3�ܝ����q�xA�=xm(�D_E�pmw�TЅ�極`ˑ���H�[��ϙ�Dvs��&t�C�w�&��-y-b�o+l���+�Y��҈^rT#�ĺ������w����<=))��M���IS��PA?��Un�����S���z��o��*���mlC��|,��_Ȥ�]p��C����Ȅ��bi=</�1�c���]w,уS������O�ʻ{�s��'kUu�|�;>�;�Lo� ����_I5�U
R��v����7��n��W��K�`^���%2Ϳtf��7��@���<ۃ�%&�%U;օ]sMc^�I�}�+��kc{�\h�9	M*T����x�J�N�E_�c�?�]�3�S#hr�0!܍A�/E��KtT�����D�������P��{X����5��@�b/Qs-�Y�g���`�m|��g+�*�Fa�l,��\r���;埊�8*��5��9S�*!���L1�~�D�x�['��n3uV2�l�K�lf;�D��N��;�W�u��X��[t�~T�y������D�e��E�x��W�a�X��ݒQ2�՜'-A�w�
T��c�{��#vم����'�Ť8�1��*o.OA3��<2�`���C��]�t"�=����4�"�Et�+�=��T<ŦA ��>a��"BF8V��pfq���P��`�c�#������Xa�C�RF�*M�p}�D�P:U��+��p����)���v� ����6�w��d�-ſ����j,ތ��[�7W&��fKx��𮞛�FH\\ԝ	d,Z��P\��k�jSA)�L:�vB�F�݅d�
o+�U�W�������[xE�}a�H* ��#"�%=�4�%�HJ7��ݎ���20t��w@�����޵�>��������]tZQIؐ@4��{W� 6�J�9��}�_L�����%�� ����:*��������A���=8'�F~�����R���O��r���Ɖ��8U���^'T ����~"��4��{s
|�'/9 >�<;oV�bFio��Q�<�G�?绩
ֈ����KtʥI�#aC�)����w��|י�u�>�f�n��<�0�����4�1�CF�c�O~�'�o64���#y'���F�2��M�/6��`[�78Z���˭X��{�_�-5qgz��83F?F{ >:e��&�Hϔٷ�.�&�uD�W8�������<�.[���s�#�scG��K��2�����^c�8cu�	6�Z2�&
��
��`*��� �Qf0� ��a�[>^�)e�N�v���YZ=�:w����H![�dU�NtH�$h��g��+���l�s3��+�'�����:�l��N�����7(��J���O�(Z@W�)!�lb`V��Ʋ����� j&�jD�����\��7�2k�͑�ݗ"9��Aρ�[�ߪ������07���\��T�lN���^~�����'�Z^���Sx�0�ۃ��NL|�':�f��t ]j^���ʸ	��W��d�;T?\�ud�L��_0���R*����ΉG$'F�";H��p���9
N���M���(�ʖ���}�N�Qђ$Y����U@O[z�z��]!��a@��Bĳ|<w�!�y�|=i�[|C��⣭��:	s��X؉��WC��<jY�A�6"�4�uMw��$�d��Oqyi��
�Z�(��0�Źݺ.��]�T�e: R���}_ �2�J�6��r�cD4�o��(�t~$x��	y�F2%i���Y,Z�V���K����f�|��9�	d�L������9A�<��(�� �ψ��S�i��.���VL>l5i���]���
ȋV����Y����U�3ޠ�|!�9��f:u`���i��wh�釐�?���H��AZqq���Fl�	&��8VR3AQ����{3�¼�v���S���~yjYGa�q�Q�m�saۈu�8�ĉ[��z2�nT��:^���q ���*?��^�)�PÕ��ViKm��؟yү�k�~s�v�r�#�\b-P�|�$���� � 
"��I�����a^�
9�nx�p���~�O�M�[F٣���7A��AҽZǉw�\̃������"�Hb��A��faԊ@�\dӾe/F�q?1�pF�㥞�\����5�K���=Y����!�x1�E�Rn���
�pHekzy���C3l���8�5OQh.��X� g�+�C"�W|n۔7��+�y���|�8�9&�$2#��/����=m��Kst< ��v{�;�33�fP:�E�<�OwW�����z����m[��ц��>h���e�}���Qt#�-��T-�
��k�=v��"}��F6w�~_�@�_�0b�?�z/!������7Ǫ�`ǝFV4�\�����;?��Kue_z=F{�2U�C�! jD��OX�oH�۰,�"S���]͐�(Vs���Ȏ�o]$ǿ1��ʮv45CLJ��V�^��^XS�֟}��v��yyBzV�������I�E�
[,?�0��"+���&`X���2��CPU�_`���d�M�!s� �;���c�H��6��˞y��.�&�C{D��69���;c���p{�ո���C�A<�T�-��;/���i$���N����˫���b���`k?�}m����}��83ԣ�[)��S�FV:�w��*+'ɗ��&lyl�#�� %3?p��	��4�9�pѰd�D�»�(]�3�f���_/I7ӈ�J�q<�z<��Aq���oC�9Njӌ��۲�o�Ө]��-m�A�F�r�r�=�Cy�.������c��h?1�'b��׬���O��WF�/ńC�ܗ��#��0R}]l���>ϥ�j�򵟟` П��prpg�� Ņ��>��Ҹ7{��w?儵� ��w���:*�;3�հ���ɒy�M���U��+�*D^<6_�y �u�i}#E[�[mKOA��i�Y����Q�U�geV�k.�h���H-���>�4�u�����&���"G�u~���ƅK������]F�>��h�������D�w1�\�+�#�g������]t�-�����x//G�pi�ң��`�f�/%����r8nI���m�ʥ�/�QvP�:rM���֓��%��]	&�]���4q"z�������<� ͓���y���K���P)�M�\>-�U�C�?3b	8&2��F~���
M�2��ZI:*5����'S�1�]��@�y�xቖ=�n݊�~���$6��]���v�.���!�[�?�׆�j7I�U��m�4Q�\9�c��t�*Os[���Aw�'��խ���={=�Y��n;���t�%^�^����E�J/��ŏ�H�K�`���#pO���c�`G>b�l�KA��+�y�/��~§eNv{iB�h�i��b�L}��3@;'u�vBXGq'j��5O�T�Xhn����,���;�GW���4t�|cU�.��e��������;���������9K`P��~.z���܇S1pp������"��8�.>�mJ�lIQ��J+d�;��X�����MF�~���<lt�h�ap���oP'�
�++�y��5�W<zR9�1�uj�,aenE�@�W��i���UMv<�3+8H�Pn�z�T׵QT[h�<�����ˇ���o�K���Z3�/eI����4�=�r�Z�"0����_&ɼ��b��PJ2����=��-9��[��ͭˈ�u=6S������co��ɌT=p����e��0:�5�4�䊡~�e������8��*�J4�����-�͞˯w���g>�~��婀���{�,M'x��B𠪘��|���T�/�e�<�y���'�Y+�Ś�����KMh�`p|��o�G��~J����z�����Za��f=J��x��v6.\��~���]Җ�4�����'q�B��-H���H������%��/l.�o��y�T��7�_�p�5ݙ�u�y[�r�|��A9���r5�ӥ��Y˟�|v}D|9P�O�.}P��X@O��K�T��s����h�O�l�u��Vy��I��������nvYY���DW�Nw��y(���"�WxH�bԣ&��>�S.�0���JG���꽡�r�yI؍��-����CLڪ�׻��e��;�%�ӹ��f]yu_k��� �S�?�S�}��|l��Q8"R[]�`��$��Ua����=C b�\�)?������ګ!_i؞����n��v�ab�-M���s�:����Gp�_�)?�(�	��#lo=)�c.�ؓ
��C�-���k��!=�/ɲ�Dݰ�Zi�de��������h�7�U�$Fs+LK�p�׮%Y�>�<�i�`�W�O'ߖة�f�r��w	�?��}�n��r��uD�N��3񋛇Q5&��l%c^]�~���qĿ3�G�E�-�14U�̋��Kĥ</8��;�\��H�wGL���d����!���=�����B�kﻨ����ca3��Q��G��n@mI���F�iO|��cY���Uv��~?�޷o�=�Rh���ˊƭa�`vR.��|�ÿr�z�1kV�Fc]�v�/��Z��]LQ�m�Υ�ߴތ5e,�m6D������sG��Hy�|�z7�F� i��e>����v��	0�F�ްj�q��t�l�%򦟮��W�<���K(4�Z?�*7����>ר�<��$]�����?q��[	���O�����Ĭm�R��մsC�ݖs`�\w.����O<��3W��TV=1�x�h���[��r3�7;����=h#;�|��Z�B@Z,���[;��T��ƙa=&B���+󢌔�w���[�&���2?v�g�u��)Pf��;�\��HH�A��I����wn}�ͥ�<�w���_~����ר=�DL��5����} k�-���%��6
�����<��7^�aIp!�ŗN�M�Û��׻�C|�9�;ą6sY�^���DG��n�f>�}���&'DC+��e�s�q�>��6r����a�f��+����m
x��B�U]C�]]iŝ�Q���v��y���>�ۻ���ޢ�ö�Q�>�udP5jͤx�,��',IaT,�	O���WzQ:��䞑:���ø7@��#X�d �@�!}"Y�T������}�)��V��u��1��w▝���Q���_}aH�G ���9�\|�!���X����r��F^�i�c-��w�!�q"p#�n0'����{��0��i��W&9g7ǒ�K��Hn�.#8�7\9"��Ȃ���S�0/�.u�o�(�_��<`�r=Y���je�"���w^��@���]V�0��4kHDR�����ݸ���{�<�ѱc׬�A��X(�@�:���xF�7`|;�D�P��2���̧�7��%��C�3��QM1͉q�|���Rv�k\-|��n DVK� 3����S��q�����#]��UAL��0���c9����?xD<�d��b_�Qo�E���|��7/�[�����ڼ6�P����L&�~��'e��-5ֽ��lc�!�y���OiL�}ص�s|"���:tK�]A��x�n��XZ����0��t�d_0z��^E��W�{MB�
)�^���F��o�
���]Ҽu;3<S��e�&�,�n�
���e9��[k{4&#�l�-v@E���a`�I�r=#H�k����e�H��`|� $ѤK��B1I=4����J�T��
<�u>�T��Z8�6��N�_ ���
�҄���Jꌕ�iQ���a�Q���<��J"��2v�>��G��T�ޏ%j5���q/���H?��f�CE��]�[2�zzL��M��\ZN��LHhOP�E�s��c�dT���{��D:eJq�$#���W�D�$��*;ޯ��Z���(��(2ɪ��Q�<	M�{I�jǈ��s��+E��{C�j����ݥ<2�-+��
�l�2�4��W����0�M*Zӓ�П�UK��6���0<�Z;���ΘV�I�ˣ��c{ȩ�T�|I�|.�/��~�#��k�k�+�r��h����$��2��-l�,bd��I.�^0�#���ɖ�J��L����fU=Β/����B�Yl��Ps�g����fj�=H�`�N�:�ᇝ���Od1h_���ɞ8R h��_���9���b��i�I�8HW����|0R'�-]:�!M��5d�(�iI��m*��Kz#�����o��H�
�U���e�����W���r��8�@�Ŷ��E����	�Q��ە�$���/ɺ+�w,���y��t&�I�=6%`}�_@"����y�-�V����\�|�	8��1�)�v��(��I^�>]<I���+�=O�h��ֲ���DH���ۊv�ws��ö.����Ӣ��l�6��y!��7��^��D0�gZ_wE�_-��RN.S�P�EW��oe��������°���M�L`�z{k&���U3W�(�m/�D>*P<�8�V'֘�����/����yC�6������]�e�yXs�_M�^���k.&Jb�2S/IX5�tt���-*�
ܲ
C�D�l�C&��~�+.%�oJ8N�[�
���g��h���_�Z*-��џ ���.��G&�V��-��[,L
���U	x��C��{�S�+,�7���Y�M!}�m���y�~�N�����:�����y��:e*�� j��5b��{��-"k�Gz��C��4���A�w��«�CBR�W���Nj,׀V�-�}bS���8TmD+D�'��(z�����
�N�.�IE`��W��Ɋ�9 ��ؑ��I��W�f�,O~�m��825è@>¡s��-��ֱ:*Q�2�`Ӵ @�����q}�'���!䇈Ta�7���E�~�?�yn���q�Vh��g�\�;��^��DN�d��c߼j��kA�Z^L�G�L0������]p���1�,���Xh�Ρ�v�����mԓ������Ԏ��{C�1mJz�nF�:DEe@�(�q����IǨ���p�۽�e�~�Z�U��׎=���6�!���d1B:.k N�[��+�^H�Z�Q����a�Yu6�\OҔ�}'���Tܯ��Yϗ� �^�ԨX�>s�}��)s�b:�v�݌pf��\���<t��MvM�������%���$uCX�9��k?���<�&YY	���xu�7k|u]ɤ�֗.e��i�� ����^����42d�[SЭ��;<�o&��郺��˨ފ�cd�e���'G��b�X�c���$�r�ku�s���e��y��u��~��~�ֈ�`@��.���pa"0����w�q���1��ix$�:�[����Z���f�o�����OEt��7�D��H!�(�k|a\87�������~�8+�n�n�E�E��*^^�z@���������d�r�"ć�T�I�X�>���=�l�1��G�k9c��^�Yd,4\��ښX;ʧ^�E'����闒�2=q'v-V:jF��;�Y���|䨼Gs2�M�B��r(|q{SZ�J4����auYZ�TP9�+��?��5�u�����|{�����Bq����+˰%�����퍜3�V����|Cim�^���k�s��镛n�b�<Dza�T3�")��Tq�]��
����[�+5��ӭrC�˩��/�|B�#��
��$�+�	I���ߖU@;z�#VN�=�9OJV����)�2�M���j�_�Q:z��d@g���bX�2k脵�W�]W��ep�ا��0���]��Ӻx�P�g��M|x�wLV̓�{�+j0�����vJ�փͿ��ٍGh��Y.6p���.�i���,�GC㕽��:آ�P	<0M�}�a��X�#.V�"��8BkDK�?6� 6�V]�l���T�&��/��h���=�s�����TXIݬ`��[1쳆�T���a஝���V��G�>
�zt�`�g\G��o��7�ʊ�ah}WpK�j|����yS���'=���ɱ�[,H�NW%YF�eke�K	���-!5���	�繖N�h�1��3���*)I��'ަ��W6�����vi��H���W�f~�O�����dv�����lEuj�b̀�.�UqPur�_
ͼ:�^4G��Eu쿶���<�"=H�Ɔ�Ol���~�Ã����v�D;�ja��7�&[o+Uc���Z��xdA���Q��n9?�i�t�\jF~A�[��^Rѯ+n�f��2�e7�|:�Yo2��%{<_��TalP�O$&�N�� ����"i�W [�φ�\�i��.ݕy3�&�P��.K��Zr�� <X�4���P�6��u���#wߙ�6����D��i��;{����_n�'�������%�J���[�y�\���(��?��>�@��b���E�kKa����V[���s���
��cp|��F����OQ듶g���,����96\��	��p6�;om�]@��K�Qq8� �{�)Z��r�5�S������kw >�P�֞���z��Qd�<^KQ���}�<1A܉����Z'y�I[�?ΓU�>�?R�շk��4�ޫE�$ӭN����ME[ C�#5`6�'��� CW�${��[��i=��x@E3��z;wn�%C�HJY�#�������{ �C�M5q��RԀ6B�`3�0	��"|��Q�_lYȊ��E4�]y'��K�H��k�����,����%n/�p��'��{kx|f��/�x�E)��F�cc��4�qȚ9��5��'����r��O*��]6,<<�6��?#���+a)((�,�ov�d�h\���3�N�I�!5�xA^ ��z���T��ϔ�bX���PHc�ue�u�gơ��=��>�а�m��Lb���7��7]�
{���L�����T(KO�t�s�^��N��?*���zR�,�]�������e�����w�N�N��n��-�Zq
�V%}��4_2z����7�B�-��2B1���m����A��N�y���W�μۇ�G[��㝆1�g�Nhph���g�l �㪮.EE37hntFxU���K���#��N�_!wm��WM�>�ƀ�CD/'}Y
���_���&
��|<���hQP�((Ko�!0��x�P���8�D�,���\|sR����L�a�m?�z6k�v(�H�!��=9�2�BJ��z�%�(�)'eG��nj��YA�F�u;����S�f�>Δ�7OQY98b7��Ob����<���1�y�_��?�u���?�%kV�L&���l��^�mM��Q �2Vh[�P�rn��,�T9-�B;i�W��	���Ѓ��[�	D�uԘ���Z�_��5%���"�� #���..bMH��)N6*i��5b��d�����긝-'\S�8��3�˼�BqȘoQܶ���
��?Ca)�ћɎi�wj���M~׏5+�M�꡷5ܞ6�|w3H�}��!�c7��aqR7��>�ٖ�_��7����C�_�+�4V[k1^����C�j&[�Y���#���ѸC�z�.L��<�����Y��h�a�a�����t�JI�su��u�������z~�H �@�ch�ݲ" �|�vI$ٍ���MzG�y����7W�aNb�+�j'1�^��S�Ĝ�r����9��o��VCs.���F2��+).3����g׵�9썌��^�@j�/���K�p�I2%����:�����|���8��,��AU�?m5�ȗ����@+*�)4��PMnk�E�c��5�ߛ��5bѤ���  j�Zc�۷4�#��ff�&Nnq��x�G�dN
c��@ �6�2���?�nf�N^��2�/�(���{�l�3OSsO�x|-����=gd����̐qss緼h�)@�.���5�	�kv����Wx���m���K�zMfVHF��$ŉ�]�_�n_�D�ʵ�=M�FE��r��;C`��ͥ�B��U�[�ʧ�����@i�O�gMY=��ݴ�/�ÁJ�q�I�}X���-��:�=׾}D2���h �D�A�N����m_~vxFWJ}ʓ~����b���!F0}Y��X$?�b�3UQ��?TP������]Bh���p���񓺤g\�c;��lH�-B6S[(�P�;��x<V ������Ps���p��e��뼗i�`��_mI�C�ZC絰�5x�[`W�M�볞��|�������j�<SOga	���Y�E�k��9�s'�"�=�|�#��V�yv��.Z<���A	3f�~�k���=��¡�xH��H�'I�e���;[2��;�m���$HcoG�խ�+��\�����T_9�ayl�X���? �H}>A󹵂��l%1W��(��Oj�,G=I�ZjÀ���]]��A�u��QݼLo��(��M�.y�^%a�?I�ۘKC�ܢ;gD\=X(Ш��Ο���b��{��'�o�Rҡ��-A������f#�;n^���<�~��Fm;*��&������ц!�{f�8��WL�C��3a�O����׸�T��)�վ�Z�%�N�M���i���D�9(�l��f��9v��������X�Ce3_��or�7�+�ʟC[��s���Ở�c�������f��T�	Qg�8-9ݡ��&:vf�k�&�Ɛ���`�E���V�le�e��k�bRgGѲ��B����Ј�ac�nx�^^�Vg�����`�_8��O�#�r�����;�1#��'�v���o�|�G+�&��F�Y�.,%,��������㤆�(\���)�o��$j^��W�7��I��4#Y�tBν��0�XKt�l���Խr<"]~w��^�3�u��<)Y��n�{��F��>����4�[��i��>
T`��8�>T��E���\T|od��I�����&|���Zφ,���;t&�"�uC�m+�ϭ9r���Oԍ���t��)me}�v_-O%���槩��\��R.6�B�j�F���"���rM��;�^� �
��[����jR�	r�zۈ���s�G�\L"�D#�;\�M�d[�n��.�D=	)��f�,�b�" �=�vFQ�IB�Ƞ
�ÿ$��c�~7O6!�&����褵Iڴ������!��p��O�~pív-Y/3��ea�N]��STn��-!A���h^{��h?�Q�R�d& �`Y�	�jk��������Wr��KU^%���n��b66m���5�4��t9.����g�C8�6���d�Nˤ0�R�g�N��b�
��C�(�\(�ޭ8���HG������B��}Y�6��H�ނ|�2<����)�m߁�ܾH��oF�t:]���E��7�]���
�\�rw�*P�$�4��[r9}X��7=���Ы�-��y����a��9�dt���D
 >�3�{����0�7_�@J��TN�-�6,��4�G֞]�	}g��p����Id~��q��&`O0�"Ae�!�|�#A�\p�hB��\~���H-��|*�Vf'Om�N��e��e�>�i?�9��ݳ6V<]�P�7�@�}��FQ��M�g��/�'Q�/r�}�����1 ��S����8�P�u�Ȕg�N�0e�5�? o���ҡA�o����,��<�!���'T�������8G+���V���=A�S1`�٨��ԩ�ʱd�\F��"#/���!�_ڰ8�Zz��3�s}�>|�y�F�f�r���c��gz��V�
~���OE  ����aRjK��7(H�ᔲ��s�H��q{C!,����I�������Z�x�¿�*h��r;@l譋�7�'G�D�{�2�fַ�ć���j���`fe�٨y�q�Ə(훖�t\U��vTR��P��?��s��1��r��U�HnN�
,�����{�uͰ������k�>�z�@e8�|2j��7M�����a4i_j?1^���HҠ\ҚB����[�#��0e ��55	����/���$^8�<��ҕA�t[�����_�[�MGF��v}6�B^Y��xq;�Q(�(lt�wb��#�
�J1�j�α@!,�)5�|�Px��'��\f�W��AE�P̑j�o����$7�D����V:v���h9iO��fA+D��p��f�r}"����,�0�����~=Q
yS�ST�M�V��/yf��"1>m���ѳ\G��H����F����1��/�N��{:������n�$�v��Rם~Y�i&��g��+�����(9��aq�4�?{����$��v*�����g���N���K/o���� �Zj]�8�(?@l���:��a�D�4]&>��sE��Ms�HZ;U�C'A�ژ&���(��J��t�M�CM���"�J�fI�����;�.����fS8^���H�<l{��<(V3�� �i�����-'>�E��P�kf��O*Z�@Mc�<s���L"E�+�K�h�[E�-���vCC*�hqi'�3��]Ɇ�8�p'~�U
�����ˋN�1���m�5E���7�/�%:V|��;8���J`�	ҕ��:��.w^T\T���:*Q�}���-�,����J)k@��H�IJ�x���D{K@�����"�\��{�`�����3B��?i�u"�^�:�+6q2�\�]��3g��%�K�i,�Q��ˎ	���GCi�����u��I'��v��Vhߤ鍅n��@f����F��m뷗B�Q"{�+�*���%���T>�L�ʘ#��~�u��u���B�G��}jG��Osp���nݶ.�aU@ZI�3ܝ2�c���}��&���U�G0�V!�����ħ��7�J�S�����]�"��r<�M�YI�p�:�E-n%V�ͯ�{���r<��g�M|��ԏ̓?���ǌ�2�������G��U`���Z�Z�l{�#�_~uF�{�����j~������N��;�"�����-u��!Of�Wy��3���V���=o!__�3�o��ف�?�+k�]��a822$<�J���6��c�e�K_����&1��_�3��,����1�	��C����Z��*;-�ËaJ�������@z��`G�H�@6�]�7ep8<v"ƈq�YD���X.�KW��$��9?1I�TCQ�e:v����惜���0�]��m�X�p��n m�dH�+��a6�/���>l{fQGC����$,��Z�K����bR��*��@�w'nF)$O�Ъc2�O���xS4ζ'tk���)_;{�÷�C�A����v�ga9�Qt�+�D��qw�
ы�awn�[�S����b2S=�gů�V�7q��o�6�]�,�O�BL�|%nZJYU����-i������/���g�Qԓ��y�::�ꮺj���>;���;g�V�p��G����`��2Zҫ���E�Ya���ƙ������؂%.=܂� dp=�A� i�^�E'� ߝ�Γ��i�Oߝ7t���A?���5��ѪǗ�OHnL���:���1�In`Qps��D/Ğ1߆����6�?��X慎�ݑ]�������.�����HU=���e-���}\ۀ�抗kX"��ԕ�0ֶ����$z5B�+�|o����-Y&aźԳ�� ���z�z2��uW��QHL��/_Z)]��@Nn��E�=up?ؽ��/����k�5Ř7�N�#7�L�f���`����x�:	�v��\]T���￷ P��ne}x�F������� ���>��;��2�_�9�Խ�S�����q��[�l�j�aҬ�:]�a�C���$���2��g�t�B&�5
�)魑-\���q z�X�fȿ��j���cwď�\W#�p��R���I!����|�8�˟�"�x���ˍ��>������S�T�MC�~��
���
.�E���](:�T������׳*�q΁k��N�&�p\�����%���<&�l�)5/-�V~�l��5��i|��\���zF+�C��d���ޮ��x���^��@��H|��X��#|@�d<�����u_~h�ʹ�_s8u��X�o�yu�[R���������֦u�M��v�`��f7�O![ݫ��m�����bk#��'h�C�����J����n92�l��N��#�4�[����_A�����ϙsʟ�8`��J\NuU�f']�&-}Ɂ��b:�����������zN���+�� f (�x�f��D�ןIX6@�mbܲ�� �X��hs�#���i� �(O��9�\�|,�W���
��db_Þz����.�u�G�Gu�����Xf��$f0`�2�^�dw�߁+zެ�� �����;^lܼi�/L����v����=*���P��-�>'�/�fy�3p�e��~hGQx�ǈ�����a*����Id�+J����GjN.Md6c��|SE#˜�	��>i|��V,����!0�������C�j�,���W�3��5y��4A�CA
��h�j\Bc�xB[+֑�\�s�t�Nz�BZ� ���c�V��]�ʿ%Y���V�!���(��8	j�^I��!���!f)���敘��H���%ob\��E�%��^_ڇ:���V��ˊ��C�X���w�v���(aG���N��-��A�+� �W������ϸ���r�MVZ]��G.�M�st�h8tx����%��&��Y(�0w�~����#74',G�����PT e�q�d�kt>�Z����;LKy$#�g���ؙ��yRL�p��zW)��":S��5�X�ل��Ӂo��~��ڠ�^��� �n�X����� R��Q}�� �&����	�k��ݕ��N�(�Iq�d'�C:���M�M�^o��b�L��S�B~��﮲�W	=5�܈07�������DFH����~1�kf�.bx����%r�L��������i$����l���`��������q�S�f�QȖάcB#�|,�.�auh��GmYf�'sƀ��̘޲��VϿu�+��������~	i�jm�,�]�
Ԗ�
��'�߁����٨S���t�j��|��]
֙$H�"�e�A"�.�g���*BGh"w�_�,��p���Q���o���R���A��"ۆ㶋�l`��gP������N܀��0�ҩƇCkE���X��e��?�^�0��s����8�8�T���O��jm���M��pW�����pf�t��r�.�k�%z�"2�C�?����d8J+(1�TQs�w�}�k�+t:�de� ��T\y9��bC����\f�Y�u8c�}t���y�p��IIL�+��^i�^��Q'��H�D{3�����+ɾ�i*z�;��ޜfMVCKO;�q�����_��S��%$
��
q�5T��q���3#H�0�z C�{'���0'b�AZ%��7��9���yVWP�تKhG��IL�`������v(]���qN�T�q����WuD�Gz�k���t�9q�/~B�����4��)E~���j����$��>_�:v�F[jSNj���%'s��}E8�1��0��p1�J(��Z��m���%�����Y��::�0x˭�n�0
�a��� i6F\e�G�U�0��;<��7?iꜬ�|�����Ȍ.��9.*_;g�#�ߓ�����ff����i�j��qcǊ�-(y����'��Q�3~I�S�5u7j�Se�a/����z��XO<Y�$gh#�X���h_4�^��܌�-2}D�jZ��tS��;�j@��&��2���&�7�V�x�Ҟ���DM�Z[��lh��|ۉ�� &ΔP �_p�v}Px��)?S�7z��Y��z	���P��aÊ���.֧-��X�ߑg0XS�~O��}ف����D���������E��Y��v�1��p�vql5��6�5�	Vp�##!!c��G�3�{��kIF:Ϣ�r�Fbd*�ur�{Q9�h�&�?��-g�{�{�ԁ\���'Ea�q"�	b�Eἱ�=�!2�>�B�X��;�B���ⅰ-��' ߝxg�|�����f��Â7��~��`�x���0E��W��4�?���6�8���Mq��ǯH���h�A����l׊�����V�Ƃa�W��k��P�b�M��5Ԗ�F\�鸁���N�(���vx\�V�?�&A�b��R�1k��e���oR�e&�3�m��,ؔ%���Vs̞�65z4�ۄ�ܮ}��<�j�ѯ�@�|���;��5�gϲd���f�6��3QU��9�ʰU��ģx21D����	T�xa��҇�)LhV~Ve��Q.��g�f��<�߹Q dӘ�K}���QiX��xH[=Yj�����?����到��-k�9ŖܪU�]ܚ�=�ϵr��5�j��|��2T1����Lʅ]��t���"U�U#���~�5E�;"��~�jܴ`^Ə����m�њ�-d�mUx�j����si��ف�5To�,��`���%`��Q�u�,���O���lV��1��|R%�t��T�W�/�V�I$��OJcڋLsv�x��D�#X����xK��	��&9Ari��5�[g�Z�ܪC�����+yYՄ����H8����M��p`7FGֶ�1��樨
��υ�YʾH��O2�Q�fY1��Y4�I�x2v��D2�vY�| �Y��5�k2�F��*(�" ��x;��j����>�ۃ���2k8�Ze�Ӱ��,�
����e3n��Q���[O��2��T���G8�������\�L�"������O����ս�^/I�y=�[˄�.��x,���B��C�41����iK/	����&�)^r�u��췥PN���:$p�y����$fGV�̛i����
Y�>\��ۺ|+�Y"����D�뿩�v�UVsȨ��#�ݬ87�Z\�����H�=4t������8l�����ֶ�0�cY~sB<�3����ı_d-���x�)ٯ�A�d�3���F�h�&�ɬ�*���z�F�����@�gl)�C����ܱT�֚��ϙ�c�G�4��V���O�d�+�~ &���/1Ü.������ʷ��x!0��3�L�E<�$�*�&5�=36���t�*d�+'�ٽw}=�8>v!����+Ƃ���g'Zg��1=��v�O��n!���C�� �-����,���o�ц�Չ�>�ptuO��yL
H����OMˋT��9�kd�� O.l�=dkHG{ jUզxt+i� r���Q��ҭ{m�{��������R��Ǿ\iLջb��^6��s�#��p|$p-O%��`��3�tɏ��C8�u�`���ل�uؐ�@s��Z���2z��9o�I6��!�:��X10@�P�'!���ÂN,�\cE�A�w!�k��A}���u)�i�b8[Q��X~���˲�u�	�y�^����g�d��Vws�U}��(����t��+:K�n��*�kXN>712v���:��l6k��u��Y~NK�B����v���T=-vf�p?�����������r�Zz�J�<���\V\�M#�m����Q��F:��V�_˃�=�>1gF��#%L�X^��s�n�@��~����4cs��R�H����h�C(_I�C��'C��m��ez.�XV�4����J�g�k�je��_�ׄ޾m!*"ҥ���t����HJJHF�D�.)���"ݝݱ�	l0���y~���kw\q����t��]N���oI�5fՑ�Y�ӹ^������_�����83<S2"�0�z��_ϣu�h��Ok��K�V��!Y/��gf �8���D"%O�5��k��%&cv�-�y�'E�)aF��b�8hZ�`/��+f��W:h,��#�8-i�����yF$,�C7F������/��;<�[l}]!��)��[5�$�y.�2�]u��{���^�h^�X��v"�+��ǧ�M�V�8�M?�h�b���'O�W,�,��ݷu������x��,!�_

	�~�i�qE[p�x��_N��=݉�I�S�����b�f��h��%�8 ]�z�L�/"^��*u8ZF����(x��囗wh��(��A��n�ܐ- ��I�Ӫ�n��M�?S/�?��c�y�s��Z:b�:�2��Z��3ّ�[��,6ﰖR�m��S�{5X|+��EF=��y_w*�}e�v���[Gc��XX�E�B��L�C���\ԡl����%��z�l���㤘�{����ZO��£ud:G�����'(لpΈW�N�e
 ��_��h�C�.��a���e��I�g��t��kW��g����o�@o�]�o{�M��R�_�x�=+T��'��&�ѼiFF���
_�b�e'���D专p����$�7�������e��.f3-�_$�l��6A>�hצ�����&z=�&|��Yw���9To߼;b�C��#��QM�H'Y�O_��J�<�����[��0
�G�|�������Ț0D/ô�d�~�/�5G�^3�z
R��1�
H����7N#od�Gy�y>U�@�|��"�i�5��yY�䇆qO��~�eQ8�;��r�	s�sR�y+��뽮r׶V����&�:m���I=l�'�-p�nUu,%��f�b	%�uI�/>)O>����{�j�9���a�����c�'�1�9o��H�t��Y��2�>qE+U9���z�r-����@M�O�q�ˎPB[�����l� ��Y#���iGk}�[=b���U��C~ARU�CZ=���&K�h���[����xE���r��$����1u�e �oك�(�j���'�����D6�c���J�l��1����irC8_�N �U-�4�;�f�	˒��p��m�c ����'boŘ�i�f�0O�B5تJ���Hb�aE�;�	z2�?O�5LC�6�:��ɣ�ɔ5]�>`��H�b��r@����O�m�ܳ��W�fW!z.�mx�����u
�C���Otx�����=��v�����l�Y^Ș�Bi��DR�/w�Fi)�$Do�����>tV�y'����590ç(��録����肜�Y/�卂���Y�];�V����O�G��V;�Hd����C)�4;�l	I%Z��Q�qUc�HLa���?�_�e�=Ah���)堋��HK���Ep]�K�5H�Pd<5�;�k�I�J	;;qT�V>�j!��;��}��!��o�c�.����w'C�Am;�h����c�$.����|��1�kxr�C�l~��w]�ֱDkV:��)��x��Z�����慪��m}�z4]������9�5�j�{���dmHOȄ�|$*����ތ�]9͸���"����d2�+ck�I/
xK��A�w�$t}l����f����������n���Cq�7n:	��g�O��=R;�؝�ʹ:Y��1v�|W�T����yx�Z^����xqs�d��-������]j�7#�������S�!��^z%N��j�ٔm���ڥ�H	����?"��G��j#jp跥��2�L�QM�r��Yy>Z����va��Eb�s��9�4��G2d���u��鏭�ą�n����\^�;;�F�}6�t+���E5Z?jTJ�x�`�K)�H:'�(O�.��7y14���Ι�*u�ԣ�W�JX+��L���k7�޿�JA�D�����@�d6��h�`�Wj��b8:Yݶ&/��4�$����gdWy��>��%pV�����\��BF�d	�d�j�r*ҁ��=9BM�s"y�+�L�Ҵ���p':�T�O��8Ɵٸ�)H{�=��=��E���Y��͓��Q��w쬼������4�"[�p �O�VoB���#V<9���rPf�����y�سT�|1?)׬���?��������[uCc|tc�t��K�ŢX����lX�Ω��P":�"���yHL����֍Dje?���0������$�Ug6ٰR�aR�|,�֯t,��ӧE�ku�-���������QN�7��3�����&b�o���x�����h�d� w �2Ր l"�/�H֏�׬܁�F����B���i4S��n���i���������\[�R�y:�H�)������B8�Btwf���>6�K&�譠�jF;l.�������֕�n{��fz+�3��*�����#�۩�\>
 P'��h�Ͻ�s�d<P��(����>6��y��<?��n���翰n/�˓
��ͣY�0��+�)I;ͽ��t�M�����*�J ����ũ!U&K{����
�E�/��K7��*e��e[GGqy�x�Yff�N����͇<z��XU�`�4 ���.�To��v�כ6��]��ZxJ�FK�Ve2��!�>KM���.��2@N2��J[�=�ސ54��r���!����1�
���dɝp���j�=�UH]ޙv''�<�e� �R�O֧��D���-m���v�|��Yg��qVTm�����롌-9�}�n�@����I�ò�7kVH��:����صr_�e|����~!�ו�-+wǄn�]-��3v��E���'_�Ew8����gA�'� ��~�h%�QdK�j7��e�dN�XV4�ޤ��O>8~qE��6I;1�m���5sz��k �.S��r��h���'6dZ�x52LO�Ȫ�K�[�X���3�'�����[}��B�;���x�>���ى,uhfQ?��u~ߏ�&q#���*��j#�;���<�l���7N+9����J�|뫄�bvt^j�Wd�H?
�h��
FF�c��n�<%۰��w#��F;׼s�q�Z���E�UL)Ѳ��ک��L��e+6����C�$�-M(���y��<%�7�����M�qK{V�DVY܈+jH��l�x�䅈���\��L�4�ܻ/x��^_o°o�?�;0�o��c<)�k�3ɑ	�^E�qme��$�k`�Ih:(�J#�V�l�M��7���L�ҩʻl�|fXd�;�Y�&��%�H�p2�a�M����=�|��6Uuϋ�P�����ҋ�s�+S��oE��@<v��\"Sb{q��OܿO�n�ݏ�r?��<�l,;��5'
�2�����6�*���䋌�2���CI���}.)f�9���x���M�`f�4���������2��P�5��������Z�x���"�^�08p�/r/d�E��Ґs1����bff�!I���=�ў��\+�S�g�T�*��˕6ʀG���^klE��.EܧL�(�R~NE�0#�ɕ�Q��A��k�w��V	�<�(j��[-���I7�ɲ��Nu��r����a˨�/b�q��l�/���)�!D<�[��=�Abk��ǜ}���I&iI�v�?�)�;'���s�Q�]6Mh��Tv��'�q�)�}*�T%~���EC,`t�f������&[�B�/�<a�;�;("6���n���!�?�oX<��
��أ��:���ph��c�3o<��_l��^	<�|�������^�5`ڣ�
cj�?��B��=���sG�0vz�q�����.fa�)�y�F��Ot� *��mU�ג�L3ʈW���n(�1y�S�;����7v2�f8�����B�Lbi��ؗ='��Zv+��U��Bz��}��H���o�P�Ҳ����=4͸?o�['�F�L@�J��2�mvh�j�fљ�����:����4q����]}��;&��� n� �k'w��iA7'��U	��`�θ՟���κØ�3�7��J+7�7�>sܸJk7�@-�v	��5k�2S�R6�{Z��{�_t��-�4lk�r��3�|��#r��(�V���E׻k�3�NO���z��I.�?U���嶦Z���zx��ޔ����~��bi}l!_t�Rg���t�c���uZD�Jt_j�dȮ��8�X��Q�m�k~��{e�3��w���:�2�]��Ӡ�쐌QL���Q��$J�v�P���\Nث�욒mP�S�ڏ�s"jN��Hb�LS�x�l;ZF.�I�y��4?3��A������g�9���~�}�w�E������?E����3��@�n9)�V������W��5P��0k�=M��Ԗ�J���}(��brЊ�t�g�A��<�)��;�A`���ؐ��"#¢��p!2�C%{�Ù��ڀ?zL�����2eP5s�y}g=��z�)�c�O�����?aR�"��	�/4�_��z��3�`k�0�;�@-Q��V���|5� ��xN�gG�H��ϙ��3��	�Kh�D�lZ�8G�Cp��`��t�\d<��trh��h���rr�[9C�$c�r�tJ`�6���hU�`�lU$����<���3�Μ_�z���p��Kt8H'�v�<8��6�[�I����֩�H��'K�PK#(�-��]��;bM�E��eg��hVF�G��S��g�MüQ2bIƐKR3j�]�¤O1^4�~���X�"4d:�W��9�r�/�d]�"���/���7�^�t�K�IOt�i!$�L��|.��C4����9�6��5�����]�?{�,r�D�!)��%��΀uǺ��D֬T?Ǚ�#ssc�'f�����M9iܢ1����]%�B�R�)~~�g��W +<��z6͖�JNԨ�ݙ��8�#���ӗ����`(�[��zqlEYk�	Gg��w��ky�wnn�V��?�����hf�pM��,�:��_ժ�4z,�$a�$��euqFH���~�RƯfĒ�������!/�$�LRy�)�p����-��7�k�Cm+?���ޚ����=�2��S�a�ޟcD(���m��z&�!k0�J�=;~l_V������ �|����U^�C�lȆ����@d��\f�Gi�iȋ�"���W��[ӎ9���M)����P݀c޳����>�{+�(V�iɨܰ��iF	��#�����@�d��}�ߒ�3���#s�Oɏ�� Ad8 ?sk����1���2#�-q۩�!����M�C��+��ă~�����%B���5Oh�j���Ƽω����<�z]m�U���e��,�L��8|�+h�9��/cB�/��M�%�Bw�W�=mY!'L,�c:��V�1�Y��i}�EF�5����wm[��ӻljT��!m��ӷf�e�Ǧ^cTLj�x�%�4A�>2�N�ܣN5����7�L$~���D��F��	J���7'�Rlށ�*pӺ}���}�(���`1�n�ɷ���/�	�یr&D~�S��
��[t�� ���6[b$�j�l��珞R��x��%3�k.�,�do�&���L|��g�>�6����z;6���4�~2q�#��>8����c�/�3 ��8�o(��Ȩ��!eu��J�o�w��]���ރ�}�߽�>�m*V�������MD,��%�3:7LX�� B��`�������Eѭ�c�y�ؕ[ѿ��V����C�����<�[��bxNdhOE8�8�׮V��Lg �AG宺�%��§�/C�,�e���M?c�hR�'>w���G��lwC%��;��<|�z4}P�<����*�]t��C�i��>����4O�V��ʤ��E�-��E�|����>ol�:C5��O�e�8j��J��HzlCS���ƿ��cA�/ �a:1#__+} �}&�X�S�D���	@�4�O�̽OL"�3]նb|DP� ��+�
�[�=]d��c>�?,��}<J1]~n���и�'d`�s����ō*J� �ou8]��1������b��m�U�_�8�x�u^OS�*uw��t���'}w�N���kڹ��|tx!����x7"EiF�bX�&��Y�������x߄,Cu#�:R7pHh��hv�� �r0�G����fx)�Y�}D�y�ǎ6rLҵo���Q3�ó���_���9sʨ-����7lV�"��?6S�}�i��	�Jӣ�m�$�:���������j���!�2%z��U��Òxu�˵x���Z}��߃���E�W!9��_�J>p�d<����<��֩^�Hj�j�@��@�@Y5%`��HG@��o$c�ِA���'��k[���;���$��!�h��'�s���a����$�p"<�D�@���X��-!ib8RX���������0��bE�BZVYH�D�mG���$�R7vѢ5;������x� �};f����}�W�Z�]��0G<]$̢C�������ރ������{�H��yP�-3����!D��w�1%S$>a���t�T��`)�� �U��˺Q�5�̯&a8�:��2�6���q���'���
]�i��o���V*��Ђ���E�.�[�@ٍ��-�o
�2�����]?p�(q����ߗ����5d��S����Si#o|�	Y}���y$��Z$q׃)�{�rkQ����۲�>s�%�?Q%�ė�
��@O�'E�kW�[v�@C
b`��]�Ƕ���w�:';k����IT��I� m�Ug'�hچ����5��3ߪ�|D�U�[A�������[���\�ڂn�綨�����k�0�A�}d�"C�}y����B�fvS��
�4~�lm�&$X�>aS�x�j��GKèoN�h�6M�\})B~ ���ƒ6Y�J�j�_`��1"F�7�	��Hn`	6F8�_Ԝ8��B}�ӧ�^�a���,��&�%�>��)L:�¤f7d'W��Ɍ��}!��o��	c����6K���M|d���S>B-���P0G�����2v�ҭ=�4jSi1�d���W,q�&�dV����q��S�Nvp�I6n��@Cr@�������<Y���"��c4�#FlG�^�A7}�)Y��1z~��ڹR�X�t�Ǣ�λc����ԝ=��W�Y�8�*e�e>~푌 z�R1	��׻)G�P2�ƨ�������N�#��!_�O�x�r�	D��]��Պ��N�%�[k0tAUo���� ��6`�{,���5����`�_�W��}CZ�prݴr��ݭ��q:]�
�� �u�"��S�;o�-X�����_��'B[:��\$9G��
���u�F�x%���Z�}8�-�]00�T�J7v��.FB;�A"=�������zc�����OŦ(��o!�z6.�0"���=py
�J�d���Кjj)�)l2Do����/��FC�HNa���vf*>�Sxe8 �U?��ס���/�#���%�'\П��e��u>Y���W~��I���,����'$��~���qu��O���RWw8c�sZj�^�Ԍw!#e���	�ת���u��՟��?s"�W�jciЭ���YP���[�-fO�й��|�61u���-vт<�B5'z}���t\�@�o�@��U�%��//�[so��+�����$��i���X㚠�C�U�x�U���#��c5цg��7e�ň��&�`U5�<�3��>�p�]("Q����c��Q�E����G�7���Y����Ao�@2�<al]�(���䒖�^1_��'eW��`{i7������|�i(if�MAl��<��˂SZ����(���}�K����bG\pJcG��E������6md�K�����&��uC�yR�B��UJ�#E���M|Z?y��� n��vM!i��3�"�!�}�#��[{��{���
��ە�� O��+����r���+JH	��GT�(Z��ؗ>�U�H���-J�3B29F��ȢyP(���l��L�.5(D�<��/�lT�_�D��įzs�_%!�VƝ����s����{�W�3�TmS�Vz��co���kɦG�խH:���	?'b��|}#��r�y�&�4��^7;p�,��m)8#t��l���kkl��r�ؘ? (�ǋ]��b~prrH������уw�k�Mk��ڻ\p���h��2������O��waG5�HJ�伪)�I<�p�p8���O@	��2��w�l���-�g� n��]��̄g!��&�7>L��fpM}D�4�6�.t�,��K0��-�+�ʼb^/?#>�ʛ)ؿʭ�<��gYx�g"ޫH���F�Z}e�� 6d�ƈӚ8VB��f���ҟ��F���-�h�VM_k9̿DH
��HM��O�i�:����3{$*��޶E�E�'`��9�����Q5h����5T6�AZ~��Z��Y�X8NJ��ѳ����ٮ��ʹ����B��g�o[�Q�#�GY�Q�a��(��u��O�L\�>r�����ٕ�8��"S���������L�_{�c��<�����A�=eb�^}�F'���D~>iM�N�CÉ;�-?$���Ђ,l��+�O|T�bdM ��ԕ������Z^F�(��鷥�$1t%�Ǯ�15�ěo��yoe�	!�j�f�	H�i�%�ڬ�+��yB����wOV���#�o?p씱�+�|ҒH-��G����a���5�w��[>������G�z"S��|߇�`ZYg4d��W�����i2�.��&O��oI�ZU�N����X�h6.Y����$��[�Wn����lKl�aΠi���.���S{�\�Ja_����$��	�ܕ��@��s�
[��o<���l@E���!�դvH��nɸ�>��[?����Kk8{�����lid�9�|a���{���t��c׾Ԧ;��,S�7�48�L� :,�#ټ��71�7��zG����}I~���?�]��ԋ �"t�W��� ������&��ETM�^~�D���c�o��B��3gp������SAh+8��'���wg���7�����B���Sm.�@���Ӣ�c���a��8#m/�-��\�aޫ���\Poy�jۗ2�D�L6��P���N��WW��y�WD���:&OQ�'�C͒%�r����s����۔�i���˯�tp��Ҿ&��>����R�}���p1��h�6���l8f�F�z�q�B�|[ܕ�mG-!����]w�K��G҇����}6���d���ګ=�]_���jN�;��@(�i�2�ۘ&�g<EH���w��2�ËKٕ��S~��Jw�ٕ�!�fE�����G�[H�oe�M'����d\N��q�S�ĵ6u�r-��=mo�V\�yџ�T�N����	;p��#}Hzī�V1��)^�&�� �uwl��0�5��1��VEF�w�l�7������&C�3;3�"$�]��^�&ď�ѮzF>�x#2_$9� �q�\5xWy�@,T|����y/���)����)�Uo�S���,����n?�B�Lu�n�����p�^{�ݰ�PEa�b�"Ta�<��8ʣN�v� ��PԮ�%~QEK;'�ٛ�N(�5�E�������H%>t��c���
�-"*�\%;lONҮ�T�d�΁ O���HM%�IMZ�>�&D��w;Xn�M7�Lт1�v�*��Z���G�K_�N��w1ۋ7�C���2�$Ք�g�0�ͯ����O?��b�kK��-�EO�VJ���̖[ٟ:�F��������#(n���,�� 9|��E]�O�Y4»�89ޙ��Ĵ$b�P� up�E�^��r/ ��|ڶ�%Hp�?�(a-3�֋�3x(Y�Ox��vX�Jg�gN-�R�I$uYצ���t����M-��(k5�����oǖ��6̃��#�?� 6�Ix=�`pI�zUZ~�����~\�6D�l�3��)c�J�Νi\"�t�L^a�M��2Z袰?3���ѩ�<ґ�ƽ$y�0��/9S�M��z�+��J�)o|`�Q��m��I������٘����T��<_��;�u!��g�ɠW�t�[N.��x)�qnn�\�=ZD�_`��}��f��V���s��Wt����yf��(1�-�wu�⫽d���##d�ᠠb4ͲI,-�UmJ̩�>a�lsy!��I��ֻ4��S̭�FD����V��%���4�,�ر��(�j�j����0��R�Z�A����]p���s�#�!՜�:�:�d�[��{͖�g�V&7�P2q��a�L��}���ax�Ǵ#hA@h+D :QL[�"Q���D�Hh��!ar����BOO ��R�B�Mu\I9��N2<���?t~�9��˫��v(��J�gp)0��ٔ{,��~H��o寋.o��^�o@"�����p6��v|�.+I�n�w�jn ت�_��󻰷�u_T
oX#�U�-�R�Q�-VX�)�V�g��xYGxN}�o�����$�?���y� (�f<�0�0�~g7l�Q�2�D{���8<@�P�:]/�a&g}�I+/7��Jy�us7ǣΧL�j��~޼��A��dzҩ�OK�F�HYٽ|�9��Fr!1���m#�W���C�i�5ByY��L3}���}���+c��ǲ��l��
{���/�X�WS���&<��2�Ԏ�|C(���SP#��s1�J���_p��O�׶�l]��g������%G<xE��΂�m�'5k�/,�����NSx��B�͞)�=���5� #sƪɓD���\�
{��l�ոBӂ}(�M�St/�7$V���	����hK�͡�Ac��hM��3���:C�%�@���%O���O.Z@]�/��=�}LZ�Q�n�ٯˑ���V�t���[���9�g�̀5���.)���Q���6�ޫ��`�P����!�9i/+N�~�HX�ٍ��>�¨9��[z �R�]���4O)� I�a�,��o &B���H���ϓ��{��g*�����W䑁b���8/���� bӛ3~
�i�,	`|�s$�2�<��`r.�'u�8��Xw��|	#��lOG�fV��/�Ѡ�� L~I��%ԾOy�!�
S���*i65u�c�l���}��J�LmO.��������)����$g5Kd��$7������""��������i�#�7��?���e|�ʌ�V��@�,��uEU�$�qHo�;��������z�`f7�����@���-�M�a@%�ތ}	��j�CC��7Ov�h��l�l�r���n����LS��(Ω��I9Mѥ02��r}J�[�϶��"�ʍ�d.�D�Ɉ��;�b�������^���]WU=C�EL/��g�w�]yi�:,w�������ژ�`<�����>BN��TL���ʏ�9�%!#q�:�z�py+���4��|�u�/�]�$"\�����.��4S�߾k� Θ�^��p+�r������X�t�5*Ư�r�gDx{P���:l7��%���[���2��6{�Z�3.g.�%VQ{�>��[���s\ж�0A�E��{�vj��i����s��\����/�?���d�o���ߎ3	S�-%���j;%,݇�Ps�O�6Q�l/���>��[�D�ڮ��������;��z���˵�����:Nč�h_�Ќ���#t��$�^��4�s�y��w��]��@9���8�ȜW�[�0U�˝GH��f�|b�}��=V��� �t
�G2]�F�%�#ĈV�yd��E�Q��T�a�E:��J�|���f����N.y��8�J���Q6<?�U�C�>�,"��^KX�m��f4��_��*�N�s��˹J*z�6�D1>d�AzƆ�$��oB}CcNtv)�?(�W��3(�_i�NZ�'��Y�� m��ۉ>��e_b�dh�MLܜ(��n'9y�'qǈ� )@�΄��J�.��`a�q���f	��Z �$}�nxC�yБ<O�.i�N�O��fT*y>:��[�x�.��3x������i�������M�Y�=S;)�	��Sǥ��H]�߸�PR+�êll��������[,��jwrSI���^����B��,���rE������K~`_�=�>g4t0��i��M�~'.T6 ))P��]�Ĵ>���\"��ЉX��.ic'\s�32���>i�� �If?����T���_����0���^����� *�~��[N>�<�Ih���p��I��i�f�6ŋ��;J�$*�O���k�@>%���O��<�q��p��-i����+�CQ����ᙈ�!�����<��-G�F��]���=��{׸�2~�-�vs��;���A'|amLmD�
(����"P�}���dx=h���Ȩ�ԯ�xq%���ή�о�N&]�rC����JM;���-��B�	J>2�!">�˛)�M]��iD;2�krt��޵�.No���a_欄nk������6�Ȃߚ-�^��W �a3���*xR��0���ڬ�����@���&�d�&Ո�p|�׊zc�1�VB�0�S���Y8��k�[��=��'���W ��\�!�'�՗I�,ZW�87���;��8�/%�f�>���N7�)"���|[�����FvJ��̩�s��t�\M"a� F��-�+t�~�:����ǨY|�Ⱦ����p����^��Bh���b�ӕwT��d��}Wo�n���aJ4Yds��u��pv�o�;6�c|�o=�|W_�{k��^��X�C_��8�5��ߝs�w~3Dߣ�I�K%U����k�������d�H单Oc�l&b����_Gn���W~�ƪJǧ��p��φ�v��'P��R㊧�E���q}Z�O��oj)��Ie/tO���X:3
�]��D�MZ�b��i���>E�v�4y5YX���<��}{Y�� ~��
�ӯ�N����[��#xݨ�O��f	͓�7]�	Z�0��>�� �Jr�^�\��٘�c1Q'j��=	�����=&����Ϣl�.��'n���q�s�bf(�,��ud�����/>e�%ŗq���s����{�wϠ��Q�z<�6��1�>KW�q׌D(�X?�ht'sGHz_jK��5v �JQN��P彰�,�OҰ�TQ���$����z�tr���jR�B��TY���&]�A�Tj�g� � +&.�.E���<��?�8��3SΑ�l#	\V�g���-��-���!nO�f��	�W��n%����vĽ�}�G@;�V�}v�d�]�Iֺ��6�G��Y�눕��;ܾ�	��6�XV�����ԭtY��ݷ�ӷ�o[�U_�pFK,�w�7���,.��c��-�rK��;����f�Y�K��B���	̓8��{Gg�@�. v״�?�����������t�W��R� �������C��#�XZ4@ԥH"���>��䤹��:QP8�����}\���5f盒7�BF����;��і��V΂s�#�í��tf�ι�ocu������,�zkH������l�$z�q�~C�/�a��̝�i!�Q����Y+[��7��<V�P����!��؇�m���X-��I�)���I�"ƺ$9�F4,���xhX@��q�l�~�;��K��N�� �bP�
ѳ�up�%Ҳ��Z�͗�X���!�P=� �O��Ƞ��>�U۸���ѡ��l>ϑIX�e��bج$��#�<���c��$��n�M)� 8��5��0Ψ�*E*�N�DQ��.>��tzO�G?!?���	�V�;xk`}:��S`u�p���β�*�R���O��i��
�ycTs|Q04�V�yT���	���3h-A �(��.<�+�f��Y���b57N��h�G��kNX�hxJ�\E"jHZaP���k/#)��*$��#�>����D������qq�t$�S�8�}4h?�\�< 2ڂ�se�(�����U{u����LsLn�@�<YJ|`�B=�Yq2z��y�h�`R�C"�/���|���q�
�[3�1�˧�����E� 	�l3���{,*p�DP��u��h�Aws��49+,�D�_o�~M��=�PX֫�	��4;݉�ޥZN5zڞ93�̯*�fВTI�|��I{!R���$�m�R(�~�I]~�(;�-$���'UK7�$��V�0�xe'���ծ��h��H��_*~9$����6Staz�h3���8|�?�Z\"�~t:�#�%�L�~pGZ jؼ�Ι"9��w����R��P8�W#i4��c8&���@�a����u3C�/��D��2Lm̜�΃�,�Jk�#܋�z�&�ȼ6��H҅U���vV�SQD���O��ψM�]U2`�H���p�?ɾ�v�s:C��'1v�.(�q�42��
X��t~U/}�3�9�sB���VƉ�߾a��xE�|��L�g|�)V�����>��R�E�����7F�ZA�8� �V�w�{��MG~��J��F�5������2VG7#�Ѓ�q��I�Kۗ7�+�Df1��Y)Қ��Ph�$��	Ԫ�kB����2��� ep|'l����n��l�B��Oo��h�6qM��[���yI�pv�v{�gk��Gl�K@�Qy3��O�4��9pG�|�c5����Pu���iP��_��ٓ�,��թ��U:�R�������$G3{�b�k.��x{~�P:7\:n���?Ž�(�d�m
��綟�Mi.+�E��?�gb�G���/��*KI话òZ���#���,��%ބM�Smڊ�3�^�9
���v��R飹����=2��Ŗvs'�(��I��gF������g~d��%�a*p�Ӑ�^�;�bh��%��L��$�4骄�+�|����[�*9�v�>�y��dJg�)��堑�t/�(14��a7M\� zԲ%j��8��4p�0���ͼu^=>�i�4��c���[~�)m�q���KF/־��U[�g���c��b�B�@p��$� �وw��:�V�1 �b/��oM��h>���vp����NS��И�#"Pm�S��^�	
�",�g��2x�p�A%<��s�/e�O��yW�Hw�/��w�?OoA���u���|��=��[ �o��.~	�����x%[O�c���*B�ښ$�MW�ı�5��X7��1����Hl��ݤm{����
;�kf1��s2��&�#�������-N�+s�����37�����O�5m
q��ڨ=SL�*I�I�jp�k(�K�1vA~�$�3�]��������Lb{��eF�����)�y�����G�� n�w��j)Et���= �r�ƛ���/na~p�L5���.����8���~�5��75�?�y�4�x4�������u���T��n��y�7v�̴^�B�Ғ�BDJ-��~m�cL/�˕U.�y����mب.Y*�r�/.<�����G�fM;��p;��
���ƥMX���Hbo��4K�͍�j�q(��)�Ia���E�*��6
�%��\����IC%���6;i��W������w���r2�|��->�n(pα]��+|$�KB�*.��HcߵJ[��ޡ��jw���*���'gk�K?�8��#h��ߪ?��9c��P�$��bL��fw@H�b�{�gi&���<�k��YD���Ž$Q�g�d2���$P1��,IIgW���ܴ.�5��;aq��ݶ����	9��@O*L��ΏD���L�t	LJ���n�ȯ!��%xCQ���Ѭ�.]�β�#+^h����d}M]�� ?R�ĆQ�t0�~��b�a3u�r�U�e	Z������e�]zX��n����b=i9�^�ްe��L�E�I���tяʬ�!&ю<�
&Eqo���?�| c�(�îA�o��7�^>���b)�i ��<�X�I8_~�[�.�J���|��ʠɜ6<��|>�Y���7V�+��َ|T�iV�=z�S�F�����j�T�崛��b+7��~z�F}ىwº$O ,�By��3sj�#V�no/��2��j@�o��fM�S�
�gy^����[�TD�/v�!=���
$أ[�\�H��~uhm>0�N���sj7W��0aH1�	a� 7=4-�;������r^>�����ghx6��Y��k��`A���<R��J=�A}��r�ѳ���!�%�ˏ9�9^�:
���	Na,�Z���J߃^��h_vU���#
}��u�.� b��m�>���4/ v\�d���@ +�%��4B���CK�e>?�����zV֤arQ�����}8����X��،�*��_��)���m���,b� �ȟ�9b^��'cu��E>(�?�ӓ���P1��4�,��yG�շB���y,Hj`��)'�֪��l���Z�e����<��	�ޤ[��a-ӊ&ߵ�w.�$�b�j�Us��Z����@�o��R�����ҵJ>vx��/H9������_̇�5��4i]���u	 =r3���O!Гv�zs���H��~a�r�H�ָ����_hU�bF�Q��f9��,i��,Vi1s��g/B�|��_�6�q�wk�'9�xy�g�\��q�bMq2NuO�ɩ�q��Q���`eT,l@�R���u3-��6<ٓ �\��T\�#����m�RU�RiըZU�v[�vmJ�-Fm"�^EQ�.�{o�7�C{�H�������~�{��=�9�s����}�[y/�����M�%���'���t��'�k-��	��Ա=a7��k�kT}�ۛ~��8�Ƭ�����2v���z�k��eMf��To�f�[m3>,k�c��x��&}��-�0q1ٍVk����Iqo"�CÆ��κET���F��;?���:5(a���������~[6h/��!�Tx���#"Jbt� 3TG|�����0|/�0�SRw<i�<�5�L�uTC��_� �L�̔A����y^%\㝙��ݻ[������Q��������յ�;dSs#�k�J%��q�:\���)·J
���W�AE��|��g�w�4M?�Nm�L�찥��T�9��\���Br��w��/@9���uQq�xV q�Ǽ3ܗK�� ���$�et5�vM#����]�
��oT �4�@6ng���l4c��*z(���W���/+�k��gؓ�]~!��1���'z��8��I�\)xEo��6�w@Q����ގ�}/���)!���8��dP
��H}��~�l�����N#�jT����P���hU��0����V��B���{���aB6t�;���#�D���u�]e@���]�(f[pq�^���4=����&@X\mj����u���S%�*{��{o�Bָ`Gna�ȴw%�ؑ�P��G�6'�mZ5~U!����h�6BdǢKzP��տ�XK 8�{�~�5�����OP�r�������wYq��	�N��k�����zJ�9H7
 qaWZ{|vXs�#tď�F�h��B���֓��A=�����P���]������Y�V����K�M3	��)��Ry�)���J.:���2~Xb!�wk
kE��~�c��_.%QƊ��I1@m�TG-��j�nR`����o3KA�K=}?�z�E�|�Pua��!|%o6Q�U��tUi�G��a�:��I�Gɣ��yU�'?�e�*(��+�f���]��܆'����͓�z�y7��
�,�%z��Isr�Kq�s��(Բ��f�N�����ҷ������I�5g�Q�{]��Y����e��ғp�V�P������ѧjlxe��&����:����"ę��ffODF*|Y�X��`��d"�z|�}�=Ƈ���c lv��՝��G���z9�/|�����4r�w���f�
�L���f6�lLA�X�ڤ1��3R�aٻ�d�ڍ��.�{������C��n�&5ayY/o��� !B�{22��g3D�"���s�Xc�}�$>�@��� ��s{t�������A���&��c"aD�Ҵ�(�HʌM�C����]V���4��w�����Fu����}�؆k��l;>��T�,�S�e�bպ}"08���K��38�{S SB�/_��֬�����E�W�h�#�� �������Y����˴�֊�:�o�w|�5O+��*��~��JU�=<��#��*����)=޹: 8��ý}�4.�q�s왮�?��!��jy�G�"*U��-3�9�Cz��3d��
Z65v��"d򳰫T�͟��	�<���=l#N>�Kz��,�>'1�'���I��aU���g�%"�o�#Q:�#�"5��#�=嘼�9z��qNd��Di������_D�]UCw TS(X]N=E�>.Z}����+��֗��p���a �Z�5��q�t�b��CM1����q&�=�^9�dD�쟂m�|1C�Ǯ�J�a��e-ǫ-�̞������'|9��s�ΰ2�F2������P���mS1;�N��ȕ<���!VU��c�������[~��I����_q��Q[�8�@:#h�:G����������|��C����^C2��iV��<qW�MP��I�붸»M�L�9�ބ��f���]���>�(��e�S�6�d���z��-��c��B�"-�n�3z)�֗Sg���;�d�[�/>'~8{4&@�[��>�[�ҽ�q�pt��I'�N�'�pV��-͚�VT&4F_8*ݱ�à�'KODh��s�70~����j���/Iј6�����g%�&���0�fi��7A<���jZ����<���W��ȭ2�L8S������A�%b�g�'qTH�]V�i&h϶S���/|T(m�����>���ϵ�C4*N٤����u[�y_G�[���l��߻P}�ԅ)Bꌱ�U)z2 ���*V/�f6�����_�&h"�+<�!�Tԏ�j9�3zf���el֜���E�[��ǪՋ��2��t��ج��+W)4��$����<��z�ؚk��rX� �bOO�+'��鏻�O9B�P_rB���Q�-��[L��K�K�����k��4`M���2��嘢aMo�q h��c�l�D������lO�طQ��	z^�xR�ݚ|C��(X!a[��������(
M�(.��.a�Ǆ��Z��5��_!siq��@�x?&��;ɉ�p���L�R�{-�q���|oA��KǤ��Z4\��=Jq���~�G-:�f���G���@얱���q� {��K,^�s��?m��ө��r���X��4�J`�-+^�PT��;������M��O�}�}���!�Ƒb�;���K)���p5�y���3�7���p5��f�K�dKM��k�Z��H�^�rL�շi�v��Z.�bq�w��&GGz[���&O4m�WURyB?�UYi�R�(��m��������x+l�Y��5$ ����ûX.7�������Gtew���&�-#�=�<��#�H�cL���S?����(J�)��j�z翆s��Z��5��)ɧ�n͟��&�Sr�cy�*UW���*�L��p�����e�5��"8�{��I�ޝ9��<�N{��e���S'�}���|�W���^�0�*)ʨZ�̉%ؾ�U�c�{$�xU�BX�z�1��޾t��=+��E=��"���?t�L�8|���=�~�3��i�����L|<sO)��_4��,z�cQ7%?�W�#ł@m�v*(�� J�u�_B��n�E��a;�w�H�:�&	[T�T���z6<J}�8������BSG��<Oi��E�:b��T�z��{�r�@ˡE%\W1{d�9�@���(A>6_�ӆS�������Pg(yi�Oʡ�2S�v�DT^`�%j�ۢ�h�Qg�U�W=_�>��۞�z��6|c4�HZbY|�t88K���.�nEⱗ꺲b�Tͧ������(,�3��Ju��푲�vկ���i����w���	g�d'�����`#2�����m�u�K� �������p9�q<4���Ra��) ����O|�2�ձp����J���ns�*���<�7f=y��e�܈�h���g\4�H�e�--�6`�����ᨴ���ٞ?�Z�V�V\L���QTM_D�M�0����@����H��kigIh�A���!vP����ME��fYb��'`�˟"��ֵЖ���:��rً�ߴ6�V�>40�����]RZ�p�a��;�jZD��t���ӲO۶����vjޤ?���L�-$�H��Iĸd�NJ������Owf��C���f
^�'v��_�+���b�^��p<b����1�{Ty��������'�΢$Q�����E=Z;��]�g�v���/?@�#��w��J�.`U���� ��o~��j՝�kx��*í�fw	�>��x���y��ꤥ��)'V��hy�sHe{/�rb����/�R�4_�K��ՅZ�]0}eH��ep�9JBזϫ�=t�P�r����b�B��v����1�7ǏQ>��J�,S�C0�K?�4b���s��K('�"Q�X抌p�jO�8�#�/a�ގ���&d��Q;���R{K��(�$;q&���$�57�Z�'N}ܳ"0�ּ����E�i���܀�ͼKҶT��|�P?9d�'��ER�EDm��N�;c��O}�No�m')���ި�{��魥�l�YiA������36����wN1��0��P��iv�A�\lf�Ǟ�[�J���ؔ/G�.����'���Ӊ�S�2S��uG���?�6�u�Fmy�	����a�� Gd��q)�ձE
c�"�_/���m\߇��������o?'�܄y� ���s�pi�z��,�u���&�	G�<��k�=�ۤf��])c>���u��/q�/��f�
��<����@��/��q� o1r	gD|�d��X����dm��~Q��&Yu��DZ�t{���ֻ2�8P��V�XW$���\�w��cG@���n�^ր��tC��ܕ���E�^#'�w�Ty�n�g;�h�9�0�2S��8Ʈ�Dv҉r}�\�D��-�6s�_Dv<￷��C*~#�� ��4��x�<ظ�[w�J���Y�� �V�9����I�b�X3�K;s�K]Pp})~K?^w"�����~cA�S���t�0+�,X�sd��-8Gm�v�/� ��-	\���%�g�̤+�6Ʒ+ w7���D(v�1t?���1a�[��Q"F����"��-2c&�̻V�߿�>3�a}-ЛBm���ۭ���"��!g�]�E��f��d�eYMo��H��E����E����9�YU����P1�Xׯ�s2����K�
���{h�J)k���t��>�P��X��G�<'83;<��u��y/��<�$|��	��K����MV.���q���j��k~�>��C�]#T��~֎%hkR����$��s�p_&K��PW 5��"a���i���F��b?^����?0�,e����Dq�J��he���ʾH�
.��])EE�mA�S|e��e�T&V�[G��)�~���@Sו.S�ٲ��>b�Al4�7��+���e��L�n��NO�ڭ�G��Sa�$sL=xfi�C��o������0~��i��9:0�ծ�t?�9:�z�z�����=��HF�0�9{��y���x������w��iH�3o�C��w��K(���[��|ۄL��M��w a����ЂR�j�F��^��k����Iť�L���e�&�Vf�uI܁-��_ƞ��N���qKĊ�#^�_fM>����y�c�©ڧ�?	�Q�HFn��x� jF���wA,~����l�Y+ݴ��%4�B���TY�w�RH��_�I�ʚ]q�4bP�A�P�QL�z�w�! ��V����3י�����߉����uWhN�c��\PZ��^�;g���\Qd��Β��
���-H�eYJD���vwQ��t����Q�.6���O��q�[�mC��r}�r���kd,�f��\Ѽ�Wひ��f�|��6��8~^����R_7�!���ґ-=���p>��uA�����Q�7�T���;Ӭh��#aQ�r k:�E�r���\!����F�-�ܞ5���:��I���m+̈N�*��'���>/?�L!)��r�Iˡ5�a��8�=4<gP�tʮMܝ��+q#��7�T�d �(M�z:�4�����H�*c4f����t��
�Nݟ�#I8ˡ"s9ۀPyE`�Le�d{=���ʁ5ړ:�w��\���>.�0fq�Z8�BFm����#����92j�d�����IL�B ݁�����߻�� L��U��#��l�Ǿ �1��]��̧��)���'.��{�O�]?p��;�}<u7I�+w��8m��.U����}�{TG���ϻ��J�*�9�,�t�qy�ZxN,%���9�҄¤���>G�����%=g3\��pyT�@��B�lyZ���'U����D��w)7Z����������VRė�{@��k�����f��O8�
 exM���RSR�i�۸�1!���^�)���?I�w��o�JM��*��/�]�/����(��RѦ����Jz<��`u��X ��&O�h`6GT���.�d��ޱ�3��Ui�K����V��Ӈy b���ŤV*�FH�Y�q�sP�j�co�ؼ��l���?��\z�&KiP��M�j�b�)vyO9�Ͼ�̑��ɖ3?���
_����ңBO����ߺRm*� �>HQk�-���tEg)_�M��8��!k�=��2�@�l$J�z�vھ�P�=t\AD<	c=zb�?��~Dtbd�)�3�L�O�9y>}���-g*��ï8ӂj@d�H�A�ص }_��x�FoU�����ͅӫhp�Ur�g���N�2���%tTS�LitAj�<v<"e]ms��M�������TFH�#Y��;R�����>xP@�Y��c�;��0N�zdm�ڶR���s-��כ��y�8��%�,�ڕ���r�u/��T�wJ%U�_�B��+0�p�!9|���繀䟴��bvg ͑<�5'�"��?Ns���y!���:�]%�ty�$\�����>��; �Ψ�3�u��s�O&�#&����-�`��os�R���ߒfukS�#n��5E�X��-�^i�/�T͢�����=�E�Y��t]���Ol�Or@��=���k~1E(�/��ׯ�F#7^f'��B�^��� �_${bt�8�i���5�����U��xtJ�1[����A�DNG���f,s+����z���|�MtN��d�E%�E�ʙ���
lcX[�Sir��\�@��΄v]���J��Z�.Uf�]���(�\�X�vL��QrY������{�<�@w��tʔķ���O2��"�Z��&�7Ѭ�l1��F��S�ib�8�	���,��ȧ�)m�d:�)��ֿю���mr�ԪJ�5D�����hA���;�p���(�*J�?O
[�>��)pAˑ5-!dУ�ԛ�E2�|'�f��PD^cqNC���YX`�g�����<K^� Ak�iOߧ�v��*9Ĥ1Nl��lmb΋3%�C��1kzV�F�ӎ�^��ؙ��@�3�����}�6�4ԋD��c�Dce�Y�Q�@�G��R�{�/�t	�5�5[d���߼�^)�q �TX�kŀ�w;�[���7ʯs�,⃶�e�N�v#�pe��	��P�� 3�@{MQ���N��ƌNuo����fP�9�"/꣑���~f�Nr뽉\K�Z�{%���f�b
=2>�V�|b)��q�;��9����?��"Z<�D����[�h�~��J���ݍD��Au��]�2AÃZ�B�o�7��������c���n{9�l3��937�j��.[�N�_�U��v�?Y.˖>�Q����+��|k�����V��bO����>Qқ;�I|�S�@cS��tq������AS<v]N-�E��+�5��q�<���nq�sDk�4Jg�ц��f^�Y�����`��#|K�K�Yj���\�?5�M����q��+;Y~{�۔��$h���� >����E�9�eK�QI�Y7�.���H�ܓ���}�@��Il��e���hH���2�98-vƴߟ�mc��,��}˥r�O�4���o>��I�э2A�鈅ң�
< �G����k�_�q,������ې�[��7ۯ��u]�~���.A�s_GKW�:�W&їƄ��OZܺ.�Wv�X�~���uߍ�H�����/�Ե$��yI�{���@�����|�5��h�"K��K�E�5���z�����i;�Ӕ���#�q�{G��Y����HR�1�-�
3Q1�kB͏��Ț�2���Ws	��G�o�"R���k��1|��j�P!&��:�l�b�)�����^���［��-�gQ�dx�h���ې�����fb�c6:�.ܵ���,�T��.�y�2��!��A���GC�m����R�l��a��<TS�G
�Ym��[��A������["I�~�i׊!E�|�Ğy���U�.��K�۱�p�I�Z��ol�:�4�+7�r$|E6�����o�*�y�!��'����6������o>�I%[_���rׅ��7�q1|v20g����)���ŷ����D��>b�T[�1ϑ�����m�˸_J��b��9k�n	�&0����g�����J�Y�#����ڃ��;�\�Ol��^�a�*� w-3fi�^�4@�5����:�?�"}����+��h�[�Ը��)�(8�VH�cI�8�εѹ߯M��R��)q�v@,yn��|�@��5�h?g2��8?�}��T��2�tU���n�C��Д�!N�4����y�冥k1@�F�;5�٤ZzfG��wJ��o�Ҵ��
���z�gw�U
��Ql�/�5��[jՎ��(L������ޙ����7����ˠ�v��wA�	����fZI�]]O�M� ��v�ڣ[��"���� ���yJ�����NV�X?��?0<F�@�ko�z[z��|p������=Լ�Ϥ'�N�o���7Bc�:��?N1[�{e��k�t���/�Q9�q���Yg����2̰�$��l��pt����ُ��j��+k��e�z�ϗ'����¤GYj|�x~!fl�#��_�j7=�����O|�.'.|}"jZg	�X�O��%�F*YM��@�"���z:e�<x��!�����OZ�<|�����J\���'�jnnP���(��� ������3�sƹ
p�R6UI̹���+?�\�6�B0�v4���d�䪇���͜��%��z�^����4��`��@���ܩ���1���F�\Ub��D�&�Γ��׏�'�O;��f�'�cn��[�����I9����߉L��P9̩�]W"|��1|�Rt��׷��r���[����k�]�����9��wT��_�Hn�w�XW0(l:^�k"#ׯ^��:������G�b�YZWY�j_Y���$��բl���QV+�T �q��;$/_������;n�
�#�_�Q�dW�.��z�Ɛ�Y�H����<��$��-Ƙ�"�K�Q���B���d��/y��04���ؒ��ez��0������xG<��4�F���hՅ'�[uAb��Y�]n����=�]��s����'ډ�0@�'�		;o��<�v��}ql�ߟL�?�8��yOsE/����wVW�/�Ƣ���
�re����y>Y'S��Gz���x��|�$5z��+Ћa,��-sqھ<^���T�aQ�NlNR��?��p�M�����i���4�JU%C��x2�����}��C�׾`�����D3�3l{� "��Ѻ�Ȣ�U��q�o�Gy�F��'.��'�+
)�D�A���ɧ�׬��b��t�jD�v�	U�*�,��ïyM�B,8��F������ ~���	=бO#�2O1�)�����/�:�6���kà{9ZB�~I1j�<�ȕS����̻[w�U�:!ɬ9����Q9_R;�)rR(`-���0�o�R҅\��P�փc�QQ[ʤ��m�E���w��b~�.`�a�d�Tj[qZ�ڧΒ�>�w&j����L��M�d#K��X̍�M\�{�V½oYSL���5�|j��.JW��ݠ�A�F�^f`�?�1Պ�M�]��X-]t�#���9V3ȋB�@'u�i�]�j����'#S��`�Y��ɩq>t���hn����;��g�W��6>P�ͫ�\�� Da�L��d�

LE��MM'��px��:�ŎP�R�VB�}|f�qk�U#U�K"�O�W�{n��I�>�}�Wmay�/� 
�ଝY�(��y�L�.�R�'���_#�.}�Ѓ¢�]�x�����0d^y�4��������\�����AM�/�ԛ���}�m��X�Y���i�T+���EL����Ҝ|��9g%�n����xh��ݓ�t��}�{��%��67����k��嵋z6x���\���˱��r�{Ue�7�L����*��xZ�>dͻ�ޖ3��P.q��Uԗ�X.�F'%g�8��|VB�ؑ,x���b�k��.��}����3�^�d��Q�b� �.� �EOW��zZ[�����JG�8j&6�5�L�C�iU��k�j�Bo#p�m~K�����!�/�ʑ��a����;�MK�`g�Gi�qX�$���oV�����}�_�>�1�3m~���Q�Q���p�7/�����L�Y�.�.E�B��W	g�W^���o8��2������$�.ȭY�˜W�^Jޠ���K#Sr�$ݵ�vuvd�F��hߕޔ>кnt��p��q����= HKZƟ�v��I���>�f��Ag�-��R:�Fų��&_B?Y��@�O�}'22F��kB�b����<SmT���K��bi��5l����/�W-��ɒ,r�p�'��934%�S��#-�<�Pbg��vLo~�l}���K�M|���Y5�Wg����[ 'ªoD����^�k�!��`Ա�uY��!�S�a�E A����/��ބ�\���C���ѕ�ZU�륻��uU�Ni.��e���گ[mu��gߑk��r�	��Do�dF�5���/Δ}$�T�T*��!}&�q���?;a����)~�k�8���aX�v'��C���6:	1|�˺��~��8�vV9%��I��.��L&�h<��^sĆ9��],�D鿠ڣ��z�xf��� ��;,3s��`V�D��G4/6��n��>cD�s��?u��:I5AR=��_�Kz-Q����B�>H6/,�~ȴ��Bn�/7R�k�K��N_�Y.���φ�"�<eeN���	܀9�:�n��
F�̫�������q���n���i����}�lc����j.�M(x����tP�;}e�e��e�=a@� �q]v�u������.a�i�"��_96�HQ�!�c0�=������˾0��$pMa��[���������?ƄW�~Y�w�=�uߧz1�-q�k����e}����R�Z��-�n�EH����t<i�y���5s�lӑ0H�� �+ ��}��WBDj�'f�˩���0���W�0��f��¸H����%1�_,�'�|?�B4�x3pK��!E��kn�s#��?"����z ��6�l�mX�E�����z�E��>F�����ho,޾���K~���Cs��bff��+��abwZ�����v�����(4ʼ�59t�����Mّ���j������Ldh~wV�P>�|��zJ�F��X�`LX4�������c� �}��8�������0'��+�Ed����I��Qb_��]�D^j>
���f������d����w��M��)b�)2<j�_m>0��h��bZ�^�'�(�lۺ`� (�5�K���d�7IQ�(�ʖַp�Y��)T��e���_�^�3�j�Хuҕ����ݞ֜Y-�Y�qk��k&����LK���o񠘫^U�����Xi4�f<U�ɢJ��=�]Ў���wȪ:C�ߝfy�BY��/T(1L��Gw�#�s��V�Ì���N�kId����_�������s֓���9[x��U�S�?��P�G���0ٕ ����C�$$o��@Yz><U�qa(�gq�	a�J�yg���/X�ś�F���	N1
���D�P��N1���>⡐��[Ϟ6?|��q-��A��c$������sԸy�)�6Xt��s�O�P��kAf����p�� Ѕ1�=����ܱE��MD����O�T�>�M7Js]�Zf�t:����*s�"�s+�]$��+ᛃ�׾�
K4}�����
?������e=�7����\�\fhP��E^k�~��ɋ����U���:��!��T7��ioO+M+�L��K�*s��^�bF\���I�y��TF_l.��V1f�����e97�O�	�m�[��q^01�V�ڴ/�ɴ5_��M����r�3��iU��F���V��Y�`B�S~�z,���p�&�[��و_�70�I���' �gvi���w�O�5�=�>���u;�Z�䷻ц�U�WY��ؗO*����M�>}��e�9�����x�+���
a�d*��G��ƌW��L���O�F��X�
�R������]�>j�Ew�������.�*i	a%��bq��;�0TᩋS(놀)=���iSx�J��v)�4�K���f�<p6-w,u�Eq{V���5D�O�r�k�x��%Z����Ù��ž=��v<o���M��©C��{�#{�b���`/�⍰/��Y� �YIo`(*�K���`��;)~$ϥ,�2��vذf��L[s�ǹ��Q��ڀ�\������>��3����p����?���B�H�F��)�M��7 �rwD}'n} 6�����o��fx!┕�E�n��mj_�*�W<Z�\-����D|�¡��e�j���\�.��>�Ȇ���%���ev�LL<W���b�1|�}�zux�,���c!ۤ����(MͲ�Db�W�OZ?@y�����y����35�նx6A���l��SO3�V�+��!2�a��_C�U@d,'Qy}�l^z~�	�ݫ�`�ѳ *5��eL"[=�����5I��C<I-�ħc�Y��z��SY<��[��!�;��[�?�K�ў���k����ص(ܠ&^��a�D�}�.�)xs&Ct칅ʄl���"֙�'�Ѿ�FJعdAz�Z���V�����<G�Ή2!���0�ｲ����&/Bƾ�\�b�/����6�dC�����_���lk7���>�m�ak�G{tJ��Fwn_s�bܼ.�`b�S�;���q~2���G.2a9>�&�x#����&ƣ�Sȁl4��z2�_麏j	⯎WCI�9�._��I��r =L��En�f�p,;��H	h�����>�zBP���K0PK'��P�Ưt�����^&��h
�S3����S[�Rj/�]��8��F؏7�p�r�����4�IV�Gޅ^������v�r�^��|g~���������NS�G{#��О��)�h���y�v�C��ê:��}��[h�5���G��y�=`�x�J�pv�ژp�N�s�`>S.�l���\�n�nS���Z�Utza2&�7W�}^<g�|����XL��*�-�}9��ȀhX`��y,}d��;����/��]3g�������'S�y�g������>�<u!|�������<����
���qБ�@e$�/n�B.w��~А��u^^^�w}j�[b!����$E�޶�sO�f墩o;n�]��l9��K�J�k)7��B)��� ]�EUӦ����5���>(,�EO8x(,Y�,z]5�x����e{�0�|j��>�'�T��(9缨�R�����~��/��f��Ҽ�Mg-Me�S�l��k�;p#@m�����ZR�R8!�n������>���}x�>�R�1�c+�^�Q�=3q�{���C�H��kR��g�� tK@�L���f����:V+�4��U������D�m��r	k�3��W	���ʎm��-�B���ʴ��|x�|�-�e��7ϑ�.�#.~j7xmo���k�Iw���Е⚇ ����yyƹ��ڭ*O�}Y/J��l��gI�.���/�"���q��i"�Үsg���q�N���V!�f6Ưm&��؉^$�օ7�MRf��$$�@���m���M�O-��Q���r�y��)]F�ׅe���,���
mF�#�7������T_7����I�Vq���Y�fUQ���$3z�!��[]EJ����0&�a�`4�El�*פF�iϚp��1�|V.��,�Z�~��⛴C������P�7��G�������ϣ�u�Ā�F+%)�Z[N~���>DOG`�OƜr�0j��ߓ��'�LNg�����K�g�={�73���� )��[���5>'1��="�> a������_^����D�a��I�BXQ�	U]�P%�Nm祤���$0�Q� �t�%�a�Bz��N4�����ܿ�tK�T^� ��q��Y{��>���g���l�[B؄pvK��7�����o~��E�Y��K�>�6ƣ�|@������O8�H��2��ѽ�:�&�W` ~��O@R�WP��W�o
/�-��`������������vƍ��4��cӻ�'���:�;�0W�g��~��ܾ�U����&���b��+�e�n����[�_���]�2B��W���uX-�uz(���!��I�Zlf����u_'�4�e�ٚ�6�b�%�������t׊c�
��1#� �P$�5�j
��L�e�U��7c�QiUOAj�w��3��x�\-/�f|{M,ǧy�*)�_"�܌��P�e���O�%��.ɶ.���<�T�4B���c#�Aމ����R�&B�p�n����W�_.v�_L��k���R�t�����<��8����(�u���捖��<׎�\y�9)������ʷ� B�Q3�����|�_��8>t�A </.�u���|&�5����*G7&��-��h��Za��J�\@v&��m��6�"F��weNH���Ρ~��4��e_�&���w�������}~�3��=#���ކ'o�z;�R�b'�~p�d�~�&���L�F�[��E�g��M;>��4ɴ�Tng�O��ܛC��n�i�[u١ ە��Px͆�H��k���6���^0��~�O3ӏ��|"Q/�t�� ���,V��%�y�,6�z2p^5���I���5�#O�4���������%g#$Ez�3[������f��m�7�nPj���=���jb��w��Tr�I�ݽ�P����,��ۨ,���C�E|���H��D��kF��[�EB�|�v"�Q�+�6*�-z|�?��O)��2��Yg��Cv�~?>&��Q>)�Խ��N�rӶ�7d>�j��H�f�y�T���ix�ZQ��>Uw������UW&(ǜ��(4��x��nqo�܀Oh�
�@0����Ne���?05)�pҞI^��;y�|t��<�N��Om�.���Dd�9�]���
�}�5�繱?�7&��bBP!AF�Q뻵�ܘ�B>�A"�m�)v�ͨ�-��:X�Z��=���H�QhVo�Ĳ�W/$9�LQA+���	��JeI�N��׏<1�8���l�˞H���#a+�s�i�EI_�/�a_wxl�^4zxz�!ܐx^@�ߥ�U����T*�%�:�{S%8U����	)s���e�������~�� 9������F����Є����jw�FP�)�,�O4�<q�z��.��#��������o����Q�=�P�7;PI��<��uqK˨���Ø&񜉄��с��� ͦb?\)k[o�U�1�y�OI�i6f�|����1����@�mLD�y@������f!ԭ9w	�,�}�B��j����=[���/:97
c��(\������ī�i����3#���୯�?�����]5ᡆ�WV�kP[$pdy"����N����v==Cր�]�٭QMpiL����ha���-�,ZzUE6����0K{N~�F�S\�"n����S���t�%�����A��,[L@Ԗ�ov�-�p"2�S��H�>7y��������QJ.�O��8�ꋇ��6�(�&���;���j��RP��zO2DFB_�w���8ɳa�X�Y�n*唤�c��.����S=�7����^�T��Do�k�����"�S�Ś>#h���Zק>���8�A4]EvWx���Hr0�>A��bᄫ���N���uo���a<��{�?�_(�L��T�;*]��I��/���J�M�JO6x��e���11<���"q�'�}4����ͻ�;�M���$q�8�6������Z��R�L��#�hኩ�GyZ%����w��3���_�w����Ǩ��_K��y+ �Ә���~��z��7�U��5 ���G�M���U�D_��~�Gak{Ä	&�Z:<��	A�R���'�?�I�7ij�(�|��)�D�6˸Dw,�ʹ�I��6߃܍�f�M�Ԯ_���}C���8],Z5r�^'�̒����$��	�e�-b1���������H1���υAc�l�BW	5��v��z��*�2�F/���ư��H[�����9t'�/�8���u��.1��Y\FH�;��Ct��g�l�D�ϴE��;y�<k#ˠU�������};ɰ)Pܷ+#3��8��zvQ��oT�$q3�{��Ω�C��g�(8�0f陌d-Xfj� H͸5�W˭���v\�}����a��O� l��6m@��O��/�"�6�_K��w���ơ�v�{[̕R��d�X��ݏ�$��VT�jS�Ϧ�Xɨ�+Kg��������,�>���lc��]�~�Dnf^�9g�@(e1t���-�{���#Y�����3��3vƧ�.���9�'��Z�:�M�H%��(�vJu���ʯ�,��_��]bU
��׍������uk�$z��c� ���S����g�4�;c��Gow(�	�j�@峺ؓ&�2Y���U���m��;����Zkc��Ԅ6F��Ww%����]:ݼEo�mJ���h�=�/�֨�ʻ�~w�㰞�ڣ����Bw ��C��Ǧ���y��	�z`��V��w���(u-�Boy���E�i�̓��s{�;�Ñw��Y����mh(uQ�������e�P޲��ğb�C�i[�]���K�2ӄ I���Q� ^� ,_���QU^����S��B�^���3��^M�ˎ��Ro���2�������d�����ZmU��բ5�Z���ڵkV�Z	� FUQ�R����N"�S�V+Hb�"����_�����r���{�s��s�+Dq�<�]��&=���ˤͻ+&O�u�fߎ��t��<~Z�l2J�<��Ws���_j/$!��G���ޏ�$;�z2�C)�>%�C��O6�Ylwwl�����E���z�N�1V�[E̞�iYi�]`�IИh��f�������/)��%�=뺨r��(�=��ؾm�_ڨc>@etz�y*<B�&A$�=�h;�P{G)�d]�����3\}Z�P�}4��)U �^��+G/{���c�[�6-���c����k�����霼���\FZE(�⏍�Y�QZ[�. �H�k<�W�͸�]IS�!"W�R��uq�����9:�P$�e~��|9)Ǐ4��\C�"6�vI�u��|���p=[���p	(CN����"�v�Q�T�T)�����|�#����F> ʙB
\���tfI����ޟ;�T~�z�)�������lݏeA �/�ڵ�Il��p�RP�[��N~n�U��=u|c�+��M���*��`+���%3�U��`���!��3и����'�%����<m�X��L��YZ�\ ���ʇ��5���9A�9���#���`�Ѹ=��E���@v�KЈO�H(i[j���=�8�3w�h��R�����t�H2����gh���GN�d�y>݀cD\��߬�������M~�Ï��	�e3�	MQ#� �I�2�<�(��1 �n�rUsW��^�4�/�rh�2�v�$"^I��,�Q���މ��؎]�I5���O��D��w�����9�$d�̎Ӱ�DX`>���u��XŖ�˲�
�]~�d� {�t�N������n�����v?�`���N{㟿2]��[�u����n�C�E8�NA�p��јO��kևujq�����w�H�b4ؾ2Ρ:8�n�p�۬2����A��ߪ����,���~���;�f]�{{��؅Q��ѠK_>۰����U^`����6z4����/�<��r�Ń���ScSk�G�Mv�ɣp���KW�~�_ȿHzx��,
�JH�A�@����5�S��$\�rUW�J��X����[%�e���p������".@��}0mh�q��'�WNo�el�r6�Ut)�l�|7�Q�Qy>U��:U�P;�����Y�_U)�$v��*���+��� �@�� b}"�Z�T6�?z�;0w�LS [��?U�f���X	�y������q%�"�_�����jQ��W	m�kk�P'�:��=��eg[������5��%���]~˽��QF0��[���gE+�?�΅9B��C��3|�J�-�J{r�=1�b/ǜF��K2'zl��g�[�����zU�������x��NX	���O�;Q����/��F�U����{|��j�X8�kq�P3��bq���RY�h��i�Y��;H�;�)�f��j�ɒ</��=�Ĳ%�j|��$<p�p�� �o?��T�~'�Þ2^��l��@�@f_����Lץx���l
Ʋ���7��+���1=��]<��TX��q��ĵ�7�߷/uc*�[27�8��{�;���S�B\
d_�_�\�<��=mXk�1=7FV��즒O���L�2��[y.p��=ގN�ܕͿP 7�M���
�Vlie�D�2�W,�V�m� ��TrBŦ��N���S�'ܲ/@�z{B����-��П�+�H;�c�eG�����bf�%T�����t~zwӰѢ���Nf��wㄗ��v����|V�x��[�a@CXIOT��~�K;���;��ˤ��4.r	�+:Z![}I�����']�&�}7�k}�I�3�K���B9����]����+v�
^�K���,�M�jR��/���
��/��4b�����D��Ѵ��~���?�K�$Ī����A�V=��cb�ۧ���\l!pd����L��48��~X�"�>��a%���n�+�c*x�r�>������*���߅>�c�8�6k93ih��V�e{r�^�W�Ґ�*m��[�?Mr�����i�K���K}</��1z�}��}뼬���];�u$����W K�ru3�������b�cs݊�)7kP��*�e� ����!d��0��M�����+�wD�B��E����R�:�a��n�a���<��)Fլ����!Ƕ�R�zL���ɀN�@w���d-��1Á�uM6\o�,Lվ ß;=�����I~��˻n���K>3��G%�z&w��߼���Op�nO>�8}%��+j��W���t�ZSo����+����"�#�o������_�Oʼ�T�����sv/�
��0�M:���v59;d�R` ,]����}�A0��V6t?g�H��.?
b�^!�z�t'�n�����xt1*�@�l���Բ�����Ti���ۣF�7��%����2ʿu�β#��.zgO|qw*�3	���pX��w�ع�|.��|�{�ԗ|�����]A�L!�
�7%j{(rTh>1t��[�)�t��C� �����g��U�1+hw~�:m�� isb�]��z����������9Vwn_i˯<����4��I�%D���`�&�������S�UgoR ����>�_#>vr/6���\x1�yh4�_��5հ�]��0.�#�����_׉�H���mۗ���6�	̇���&{@��Q�O$]��z�Uh�|�Kt����[֭�j�UO:�-���C�e�d����'��6n���Y9�������+T!�o���h�����)ִ�y��/ar�hT�tFf��'M����.n"Zu����������j�����1%��0n(�KE����[��ш:/���Z�5�Z��B����J	r;�~����V1wZ�?��!����!��3s��z�l^��YA���K|P��:O��j=��Տ,YF�ypr�(6�b;�z��Hw�5�.�|�'hR�Z0$!�ʣ�{�~����~M�N��2WY��ڸN�d�T�Y�GN�Z6���Nu�����ˎ�ɲ��W�T�p#���9=�ڤkH	�p���nu�WRr�QS���w��b��5��@=`�_�DFF��?s��=�4:���F�8�A!�e�߹���o*�
���\�h,�&��q��"&$��Ȩ&�jW����"�r�f"����ME����o�VT7M�6X.�ny5?��/��M��)E)��
���0��?V��}M�>�ۼ6b�v;�8I̙%���[�U�s4Ռ��7Ҕ��F��|�n�UF�]E ��]���鍥1��ӄ���(O�����鲵�����y�G�P�%�r���2�Sӧ��ɝ{ʾc�>(���� l&`�̥3&˗��#t����nH+���ef�"̣�؇%�c�ء�=Q����}i^���~��n�b�ڿ�>ק&�C��biP��ָc����a�ޞ�;&���Xp�I���^t�n��S
Jb(l<OE�^�_m�_&e��5p����Q��\��L���c��gָ��i7u'-�$��Ն�"/�W�6d��!Z�D"��Շ��?��4��f�>��,�f^ �H��T��������٨���w�M��e��x�I�<W��n�h���#�tMm�9�}�5�K3k��6����2c���q�*e/8���h��^�(�|C[V�)W<�����f%QK|�Q2(�^��d.k�ػ�MIf�:�Nn�;T1�O\*�����B���v��,Q[�@�}e�Ax�>�=�t��cV�x��R�D������=�W�������`=� �!�܍8�'�@l�D2�J:���Վ+���G�؞G���R�-�g�R�8�o'��V�Rt��Ͻ��Q�H�UޕCU�P �^�v�$-�;�:��&;��=|�D^�8� -F�����n9�W�(POd��udy��N���l�w�`���/p����̸P�\�8��a������2�W�8������{6�~��(� ��\�L_~ҡd�5|@*�	�*b����ԯޫv�۰�ꮗ������0N�p:HͤWI8�� ڥp�Y�Yn#��i0l�
�l��{�WN�l���.��/sl�{_V'}��3#�+%�NT� ���R���Ŕ�$��%h�V��&��@�4_|��~w3A�K�`0~:�;1�wd��d�9n�1Ujy����W�T����*�_���t���	���%ձ0�9����_��u�݇��ۧV�PW��&7���'���}���7�R�n��N�)���Qd��s�;��?��w0�ܳ9�k�*�QEX�����.X\�'�H��[��č�'�K>l["�z
�����L�E3�=�+:�"��
�N5�Jӣ�̤jS�X��z�fvjE��_t����9�m!�^�\����d���A !CmygO?���v��	����b_RY@�&@��mng5��^�ۺ� 	��=�#F^�̚!J"lo�yp�Қ^�� �n�9:/���췦#0��}�_C(l49�7z4�7k���SGG 7�Df�I)���A����M�����"�;S��S�O���Q֖л�l:�����PL
�}|��DUs?�����uy�OeD/��kOf�ˬ�r-����F�6ۘ1]&�z���e<��{Օ&������ܪ�[�+5K�}>�c*@�I\�Ito���<K����^��_p-.�~�"m�t���Ö�a�s5u��j�6R#�u� �5��:ӳFWA^��~slZ�{'%��x�D4�����4o�׏�7�ґ,�Yd�̥� �|?˪omؑ�x�+u>�%}`4�����6*�E=�~�F����r���r{>�O�ɸ��p�/S�M
ݰ��"�V�&���e�h�XH��$�CJp�3��@�	�ec����_���`�'�a��9�'��~ߩ �(���.w�W��+�\�
�a����N��mU�xד��U�`|�2���&�u	�G?,���Wԅ'4lz���4.��V!�������UA
נ���U�f�BzL�4����������=E��޳]R2�!T�mk(,�Y�y� ��4_�������u@D!�4�"~,T�x���@�a�R�<I �����kZQB=��LG�T@�dڼ��M����y�
�UNT~�@r��˥�W�z��嗣`HrK_~�!�<�UpZm�]���0�(�5_��dD0j��f��qeO�Wq�S�-cZ�������2S=J[H5I�wg�{����݇�t4��_��'��F�C����q���{��!��78.����QlJ��I���O�Q>7��3I-8��6�+\�0X�ީ� 7�����.�⥺�N����Թ��� ��F�g���S[xq��;��3]��`����8_��� ��Ȧ�
�kΡk�K^�|�TNQ#i��]f�7��hh��Y��;�>��X�sC��7�~��:����㡼wt�.w�G=6���δ����̶�'v|q<�������)4�)�1&sU>��V6��;��z�;���ut�`fSBF]+��ⴀ��>,ό�)�r|-q[��ӗ���
d�Z/��5X����*���1ZΠV��f��5�R�*�f�MS*�˱չضQ2��@~��=�[��nv��܆�b��n��<�/���9Gq0�+1�n�X��aAh,�ڄ?C��v�)��N4{�e��?�Q�[��+��n��D�v����k�?k~ࠎ��2�=��A�w@Ew ������<��J��o�ןQ�]�7dg-^o�t}]&���������+R�󩕖
�yk�y����4=!<��ia�F�1���n�i]��a� ���7L�)�Y�b�V��n5�D���w74O�7�y�m�D��ˇu��/���?Ny(�����V�m��Q]�U�i��߹Q�?���|)i�-G�1�"�*�žSux���Ygab�[��]�	��@����c)\F��u�'z�Rq~O���4��Z��r����t2]�dI���f�'�����Y�_Rc��qߤ��,�w�1Ήk;k�3�"���J]�WOM�\\����FNߛxk3��;f�ϊ��Y����D��Ԕ���Z��PklOw��[��c��P�ά4�+�F�=�R���F[@�����\[�?k1AD���4عh#a�|�K!K>4��5ZT>.�\l���8�a?�`H6�NA�1�����P�����	Hsn����i�L.�W��9���	i$O�5C,i�'=Uf��ަ��p�x��\GW��l�q8����u����/B;�Ӭ�Y��	�6�0ЀY	�H���������1��e,�KNs��lw���X`r��ՅH�6鈆�n�Uf�A}��$7@���O\:z��+<0H�+]��J�h��U�"�ɶ�� �����9G�yF������90U��!���<I���\z@>������ ��;cZxN���,2o5aJN�p�yp5s}ǉ:���MA��:�C�eb\�
~�&h(%-��e-�"R
il���ղ� |a���|�G�tw�<�1����@�r�}�$�Oԃ�[̰��Wi63! �-�6�<����#��:�%��a5r.�9����R�hn4^O޺8E;��R�%�Q2_�ҧ�����_$�$(Gq�p�'C�ni�wO�2Ms]�ΈK2}�o'�_�����@�k�G~�W>��c�s�7�K���� d;���w�s4쫵v�b�b�4�,C����0����P}�*@f\��vUO����^�Mَ�hpy���[vwm�ӫ�X+$��'9n��a�c���u���D6D;o�~�"Ky5�;�#���n�D1��|q���C�?�N˦�6������I*՝��7{��������:Q2�^;���SB֪H��(ݞ���|(��y6aa:�����`sO\
����K�� ��o�Xz�Y{��O�or3����|}��Z!�����?Gz4�V �V��c�O.�ȥVcll\�шa�j�7'������|<�W�Ƅ���O�J��L��;���>x����4Oo���*�Wt�Ҏ��?Kڢ���D�&rS����iņ�:��H��	i�O�)U8��\�6����������[�Z��tڜ[J"��vjE5����iMf���XJ�{�����TT����l(���b\�"4^f�a<�n�S�òXA�6W�����u(����=(7Q�z�̋�<C�dU~)�/�e}�_'ц�=cxE��3�&IPh�R�_Yi�}��Ӥ@����+Ѹ-��E�DtrV�"�bA�(c�M
��iu�oP��Y�zE�#�I�?ɧ臺���EYM��ǏP�kS^%w[E'���h͖t���2�>���Q�F�χ�r��I�'�J	z�(���ׇS=(�m֗�IPw˺�ݘ�O�e�!ɫ Al�I���v��N�s�`0�<�@�u�e��1��}�gyr�w@:��Q��3pe���^{�Z�9���������-���P;��pL����NƎj���wN!9��w�#(lɌu>o�>,L�G�����_H&�����������R�߮�1ߨ
I���f���D}=��n�V&�#��c��n�9�"K�(����b� $�`z�b���կVf9�tr����;ƒ����LM����GP.U�=7�$Z�WWv�F�т��L�d~�hn��7�l��%��w,���u�%�����'����lX!�#_s���nn�EB�mxngHlu+ڔKu�\,yN7��BH7�E��S��4���<Wʲ[+l(����.i���gڭ�� ��&�}��Գ�Sudb��ͽ8[�r" H]5�h�=�$ lXߑ�N����'ms����¶O p�| c���h5~Rv� V-G_�9J���/��Tђ�6wo�u�vn�3���(� ����k���ad����}6��*.�-��-���?�/Q�1��(�Ŵ�=�طH��,�1�~k�����J�Y� F�M��L[a��+-|�+g	��X������k%��5��Յۮ��{�)~?6�����Yk��9?�B����{4h�q�Ğ���������`B�rO�(Їn�@Η�d'��x����b�D����*0j�yy��ԣ���[S�k(�ڪ�_�
R�r�蕣q=~Z��r-�ͣ�rZ�����8C,��׾�����Tk��
��w�|�	!��T����Y�(�c�fH��ʕ�8r����K��5{U��(�m��w�3B L�pkm���妶�Q�ۮ$��i=�n6��CP����:4�F�U�����CCm�ʨ6���;m!�6c�=��v�b�-���_ݟ7d���'M'�6�U��ԙ$��f#j3�:7�H�7�v�2��=��?ޤ{N/j���xk���0K��������,d@��sbh��F>�����n����ʢK�\������77�{B�J�/����_�%�����Aa �ғ|�S�$��E��vH�
�.Ǟ୅#27'E���ބ�����27�)Z���&�@��d��`8�e8�'��x�5z�n�JX`��S�b�-���VXt 3r�5�"���p�"&2�~��E�d�<�^~�9��kv��f�23�m2\�:�%�~୅�� ��$���qO�}�jK6!�.0�(ό4��Mr(��A� ������&��`���`�ds;!*��eM[�5�,8�7�_j�Z;g��ܜ��f���"���@s��<|�����%;�0-�k�mY�P�4.Px�+��1(��FyE[���ԉ7�f��ѫ �_짱���sn;q�/k���y�	�#�h�z���uIQ��D�]�ji/�"Ѹ�xT{�[f%2d�6+�Z%zs�퍑ai�HI��*��2Y��}�n�^T��A�#nRm.��0yV� ���X��p�X?���:Y�*�8�/$�;}i[�$��}i�O��G��.q̀E?!��v������X�q�%���/<!�����yAĢז���=Fy��ڏ9 @��F9�jF��'�(���ԁ����{\5^t���E�刄�opk��Yz��;GEir�m�I	�<M�K��7P���1�T}�{��%��p�䭻Cw�;�?���劸vw��'���X��ۿ,��1�"�o�ǋ��l=��r�,�?�Mǉ_��Exĝ�+K���; N%kf�{���[E��t�b|���B��2���	BA)lza ��w`�����<�����X������v8��i��A���;�4��/3�
l��Lz36|#C:*�xIJ�,$�����c�H/A(x<�`��\j���b���󚜱,�6i?Z���Wq^��c�I�5E�̐�E�Y�U��Wvz�b'	{<��y��UKO;�%��]iH���slR�N���jY}�
��[Qhqz���p��E"�����CRkKw��\C�)K`�2��n����/S=����x���Hi0,�����N�����/�<�P�ke� �2���^K�-2n�	��SLg���sWfJ ��G���CA�+�x�A�0��pqu�U��^�P"��f��j��LK�r�'2��1���F����5� k��Ý
a4�5u�$�Z���'Ĺ|��^4�a��!S���I������ꅗ�xV�kz仝H	�8�7E��g�/WV�ퟒ��ў�̗���"@Tm/C>�-c��~H�;��
=��"q��so��P�-�+}L�r� W*��A�����g�{M�A8|`�b]���A��R�,=�|��6w�����_�.A#Xؠ�_T����YHQlD���j�h|�ty����x�mZ�D�W���'��S��C>O��&��"�#��҃۞$5��&�?��l`A5�g�7pm)�ό���6y���]�fN�#T�1p�%3�(,9����zp���Ox���>gRxX��x��06�T����s���w�s-�UF��a0�y���&�vbD�u\�?��`�#uB�iCQ��8.%I\�jS�}E�����z;[ž��%�w-��xa;k�!\�TJ`��$3NbJVN�WZ� <B ]`/����AI���>�^x矾-�z�T�?5�{�<>;��k x���e�����AĨ��*)�s^C��10mP����������%�U�_�ݽ��x�N�_�Ұ_1��G���`�����@���O�I��&��͊��+� �,�VR_y���
2��R���h�j�.c�a�b���7l?��ʗ5��R~;��]�wz^���G��L~Bv�f{g	e����w�����*���2E|��S�dR�18��(��=��n���L6BQf�R�TJ�>�`�M�i����|��!	�P���/�0�B\C�B+-jӌ#�G�`��r9�J]�p�ڞ����[-'M=�"���#̸��U=!x����9�ap�x�������J9�@=��b�+fd����#"�z��̙����2�gD�5f�\�}צv��X�����U;UF���.�07��Wί,���<[]'4���yT\$y�r�G1���h!a�ݝ�?�>���7ގ��1?D��Xj�QS�I��/혚��i�����8�|��L>���-��t�Q�r-��}��qXCQ�ˋ( O�Z5nb��狠��;��O�X�f������tS�y��V���"�������pH�~Wm� ~.�c(��- �ȯHa:�����f��fÆ�J,֭�ԯ<�I�eε��sۼ*�e�k&��d�ں�B��'d�Y����"!+dy\疃6#u��
��5���L��#�Z���A�L��+����v�,�8�]�3�,z-��|]�OF�i(B�u)b��tu}��O7�u��؇� ֬�#��]o� 3�%��;�@̄ol4/.���G5���(7��4mc��HW�FI�8K��=���_#͞���E�]׎!�)��,ZJTZKT��Ϻ�>���Ce*~�fQ�2m��/u2m���aԉ�}w�H������AR�>��M���� �iL�*�iWS��>Ų�{��|
r�������������Du �7[Ļ�Ŀ7"@��,�|�i�9��u���� 
7p]�̫0��B.i�z��[��ޱ���Yկ����0��D�>?����]��*��#�p:x�WUS}��|V!��N��8�l\�q���&�$i���c������-��}�"��P�_��g+D���Vw���^Lj�s��,FM�_�F�<����'��7H��M}j|�K3�����DI�[���eї��oc�;=��#B��yj�1�hW �<�4�c)`	�Ӹ﬽���ܖS��ӷ/=�_�*A���th�"/���_)kn@]���Ρ�j�� ޢv������{<��+��9�??P�=8���8�~y����VG���n�^ش]����7���qw�6|'�f���H	�7v�fl�m����1��+�ƴ��%�\(G�d[@�_�7]$I���Iй��$�*�?7��?)d�K��������(&&���+���q���r�`9�M��0�geHԿ��H���98�(q�ةX���Nۛ��p�c-m�	�aE�m����%L��7��j���g�J�H?�,;�1�DѻU~}׏��f�RQb.� ���|���u��o�n�����3�a�"OO���j7����%����c�ҧ����-p�今^|�N�������2���r�4�3��{��׎<<��=��o:bŞ�׊�*�~��p�)�K�~�It�W�D��;�l{�!��=��i3��Y�p���E(�	�U�Ӈ$FM�ۮ�F�q<�`	-`9��u��{"��a��m<l!����;+)�:�QIDCL�#�D뷳O���UŞ�W�n<7rO8�c�
�}eߟ���1(��ښ{�i�����.�_���p��%-Ѷ���s��Ie�D:Ŏ����++�y�9]��W� SQ��~M"I�>��Ŀ�8�Z�I�AW����>��ܦ;�)TW1XE�Hl�X{vtd56إlo4�V���/Gܞ��6�&9��yӴ�g>��r�+�b.h�$��t�/�ݥ}i�
F��9�?�G�##-}���5C�E�Îvb�t-�N���/џ�|��ʑ�:�)RL�1xzkT��ĝơ%0']H~��v ����_�ؿr͂D�U1��D�S?�`�t�9��t�cK�N a������ �N�"�Q^�3����|�g�ԇh�}n�y�ˑ1V������ٜ�d�q��V,.C�lt�4@�������;b��oSi?�8��\��Άx��-_@>5K���U���f��v�����MW�D�� ����Ӎ�hz�x>'+�%Jm�su*~h.aG����2������_����0�=s�>8!9^|D� �V�6����l|�9c��+_�}�a���Tͫ����&��֑���ˌާ��w�Mz���j!r���"�3]�[>&�?^�ʧ��hن�pY�ͯË�=5`��$���K(��!�WH���9�OT�t��ь�*O"�f�`7��;�;�T�#N����T� ^�{j�?���%�hX<��;�%{���A��:�Tmk ߴw��^��e� >�?��&;g��� ���U
\��P�C�!�:��c����5�P�8��cڲ����h�Ӈ�`+��y���]W";��n�����Ԙ�F�����J�PY�
��|vvg���b"/N�ӧ�B�k�����2	ߨ7O����>�N�7��W�tnQ#���p��:��C��Q��Ϣ�Nw�C��X�'�ֵ�\d�Y�{�$�w���}*c���_m�N̓�"0~��1�sX�Q�^$f��L���\��dk��Q�<������$gd����޳���I�]}�=��S���f���k;��5����"c([2���y��"ޘe[Ti�n ǚ<�ä�����ݟ-u�Z'����ٝ�Χ���*ߖ��,T����Ut��w�v�9�-�w��z^�2-��g3�;�c>�ߛ[$�-��Κ.�tۮ0^��^=O2L�Ů۹Л���A�d.:i����[@�����L=�8��Y����1 �Z�X�8�M���F�����E�rRa$�k��r�;/@�C�&���>,W[���i�l��e�=��?�b��(��Ұn6��-5B"��\0���e�z�L, ���A���|8��y|�:�G�E�Kn^x�U�(��5�d�Z��C���ߋ������6�1����������.W�0�d2[��<�E`���Hn�y`~����yBvw'��P
&mwP^�3T2d�w.���Y��f��zE�E�r��yf#	��.�A|�SG�\������n=�C'�m�ç��+��>��25�����'v��������z"�i2���b.X83`�����v�nKFd>�9�X�%^�Q2� �ᷗǯ�
�{-f� dԯ�X�sKv�G^&�6�����2!�U!�3(��A��Y���g!!O�΂b��qeqK��?��1�2?�-ɢM��1kKc���r����8Il��N�A��_��<�w�L��Z�΍)��M��VߤEw�#x�ou��[b���#���h��?����76/`�g.�Qo�k��"���������g:Gbko��}Њ�y��3v�6�g�5�iwC�ycu��ĵ�ya�_N	�%�nX��U��Ix�Ѥ���c�K��HLA�1m�4���Dl=��i�Z��S��yq���[xa!��h�&~�����&07���g�;�eL�7$AFt����w�Tp�6�S����x�7`W,hk��P�P6d�eg�c�wƜX����{�������j��#�g�.�N*��y�#�_�r8�� Ҳkq������y~��jcWu������B��[�R����wty�`���!K\�
��`UNo���{�,А"'�o�]/_C���
����lR�U}d?�;�?���941�G(\���4|�������n�B���g��y;�Lrٌek��e7�Jts'�9ρ�a��>K 
ʙ���L�M�m���Wz����~yO�� ���31f� .��yg���	��HO��s�Y	�U��x�_E���7Q*���ݪ�66��{Hd]����_PI�*y�%L�r'���8.S��AYa��䣩޾�7��� C��"���M�����I�濸����3�v�C5��(g�Q�����4��gȕ�����������`&��VZ��r��'P��ښN>c	e���Ƶ�188K�����=�(Z� c����3eA���g���w&�|�50���Y� %h.14��F���~?�TM�x��{�ݳ�&��v���@ؐic2��Co��4-@k�y2m�77�IJ�hm�0c�Z綖�xB �xB(�;<��6ٚ\���
�K�B��fq�N̩���"��f�ij��;n!��
�y�d��W�ɸ�&����$c�)~�5�\lS��9��~��k�;#Ա��!p�,�ߗ?��}wBy5�`nā���
���"�V4:��E�kZЉ$����H���ѭC������ɹ;�Te�4/C��;ML�T]�����q�1f�'�omP�=�%X\Y�n��C��cV�!�Y���8qG���@:�,�,)4�\i�2�~��0|�~z�B�3�=maX��^�R؏1�I�����1,�-�Y`�e�;�-K��6��,�4у�̸_��ְ\H�����73�wj�b6�t.Qx�v��1���|{�K�m5�q4p�~HH��歋�0D�'�z0�����s�]h�Ȓ���E�� ��:(�ܧ4��]�,���J�)�d����<�AQ�j|�0���VJ�=duX�����I�}xI(x���`?8+,�s��*�?#�q��G�:�dwԻc:R a�K6���zy�D���9;����^0�3���,�����W�������{u� ��/n��.3aO�\�"R�R������*�����;jj��q�����z�'���~�Zn9Yg�`by���H�ױ���H��^�1����q���3�tyt���ܤpz�$��GI���殧;b��y�^5>�h�+P#b<cW�?h�?ք0~ 7�i!?��s��h+_fNw��H�4�r�j���qAD�/�O][W����F�����+~�tYp�9�xp��׶H�|=M����tQ����JMAF\[�K�\����%�(2�Q=��jm�8�e	��T�Q�έr�7�w�4�,#��c�J>4�*�'M
_����h��+�j|^}3E����­Ք�2j���Qk�W�9RJvz�y1�v*�	�`��{�#����s�Z��d�Ə�l�����-�²�q��ۭ>�$K�����&/s~��ϸ-�T7��a�"��rU��G�o�����_#H��1�/6}�vA��w�/ߞ9��ví�n|�%v�Dp�OO�XͲf�s�f�@�@�x�n�Y ��3Άo.I�q�%?s��U�=V��пw��5��V�,�]�q��VK�I�0t� �N��TԼj#�z��ۛg��$
h�4
 .>��V��glt��K`EMj��'��W{� �%��x�� ��R��r��13Jv�+�z�fe"���G>qy�?�T���4���X/�.+��ױl��*���h@�_�=������x]�R�P���cTs1�F�ɲ�k�z.@�B���`9:3���
#��u�[c�l!k�}��ZJ�6����!pC�c����7��EQCdX��lj[6�K������lY<��9'���fV>�i���o�)G��D�5�C;�o�����G��>^$�i�����Ûy��?mB��%�7��eh�|�Go�TI,��׫óc 0�f��������Y������=�&3�YF��D,dQ�W����n�U{W`<����CT>��R��)&/�ۤ-�t�h��]V�g㊍0���vg�x���H�I��W�_�aH(`?}+�g�ӥ�{qj�<EE�D��Z�e��goٺ[ş�a&Ӕ��,e�۞>�;�Q+/�Ν�U�G��ܲ5#�����M��e ��������n*mgؠ�T39�%�C� ���> u��N���N���x��Bp�q/4�ú{�����P|�M��b����yr�����v>r�j���^�t��*Y,�u�d$�a(A�Z�X9�s�<Xt8F�������<���(,pH�k�z<���L=�e1z�HVa�$'(�Y�N]�5��@4������ˤI�rX�:�w$.72$�-4�h|�s�Tk�N=�wOL;h��N�&��N�=\\�,���:Y6�j���ɥBY���ٺ� �׿}\�Wi��%Ϩi�i�*ü��'�ú�k�ǌ��mT�B�/�I�1�ύ5���=�7Pw�v��'���֮�w�Yp��8�3K���9V�Km�S7q�A-�+c���)R�����dٵ��g��Vg�8��q/@Փ�ZE��2Τm��ٔ��X}�kL�a_��i,���o��B�md?ѣl%�j	�� C~o@N��P�Nj�k��gn��������a7�[p>�\ �d��X��`u�,�����f���J��O�6��s5��s#��h����:���x����7��.�0>
����z���]���D��u/�]D��䓲��v�c� �����>g�'.������_מ�:���}�'z�ω���$�M�����T�d�=�'j�q'�:�?���|Y��,�*;l�}M�V1�@���`�e��2�+�"+L[OO�����~��8b�� �U��������J�:B��B�!�J9�"1�!1g��9���C�P9��36�D�q�4��|�m�3~���|���}_�u=�}?���:���r.��h�H���u�?([��:�i|皚_��̙�5Jo�,V]�O�Ԟ���G5P����,����q�V�����������=!��N~��L�O�ǖh8J��n��)��_O�~ù3�!JГ�wy�v��ST�mͳ*�S�̀�:��3*F�G��E�D�)�Dw���N��]�|�����̯w,fqQ��mw��
�Z&��sw������>G������n���^����*C��b0?��S�x(K�tZ*y(�X�ɍ�'�vKN�t=�N����|ju�4�v�J�׼�]��Y��_2�)>}�u�칦��̪Cq^Ý�5]����~&� �nz궤��Դ0�p#��ZѮ�6\�OOĞxv��Z�q�z��%��K��t�28Xt�W�pJ��锳簿�����R�/�Tl�:��s��|�n�~�[�-����[�ŝD��~0������l���w�; B��j�g-iA\>[�z�H����|G �5��q��^6�ƛq��q�)$2��5�r+KG��c�+*Ed�2=��fI^����~��%8�RR�/!��xb;���0���V5~p|�^��,���89	�����]�p�Oy�lפ7����@���8 ��cf^N��oYI\���4��tkޡ�w/�
گ��S�>}��Yġ�j�����K�g��/�gx�uD>0G���Jͷ�WF�2*��"M���B����v�L,���bs�)��?F�ڭ�kf����yH�����L7���C���R_�yg����?���TJ��&i��Z�|D�|��E���:��Hv�¤��0�v_��|�N�^ԩKTQ���%OK�H�x��$���[SUx"�zZ�ܿ�N
竒�u���0��| ��9t#�����2D��YMl\�"&#\��/v�ԕ�3w>�x��.����ԍD����.����w3R[�,i�CjW� ��[yT��jD�,[�H����;d�EPc�L7�ז0�
�Vdl�s �K3�.�dձDX���X?�H�]�N�,t�Cd�[�����"���W�;P��/��(��.�Q՘�ؖ ����*������w�*�^���}��hޅ��>���G���w�C����]4���+kz	��R�pvn�9��XH��~�\zwSC��pT�ş8S;$�V��zc�@t������?8���{�4�v2c�[.V�aI0��\h��~l�DDخ�T�%1��ދ�&�Ş�v3j�JJ�R�<v�;�׏�)7؁\�1O\sa��T������_�:�U(@��<+�,j����sȌ��/L+]�sxO]T`
���P�:�����;�7(�p���X�fI�Ox੠��fs�CTpz�j8uE�]��(��)�9�P�rlzИ*�ܪ4
TИ�}�˨������*$A>�@eˮӡ��ڝ��_�?���ԥ#V,�ވCLZ�$'�#�r��u��1�DJ���T��m�e�8_8��;粞{�0&����{�m�Gӭ�ouVv�OR�����2YUN
�Q��0Y�Ip�B9���I�D�>�>�S_y��xܿ��$HqӚF��!��2��W,5m�G��,hWk��`�+K����f���)�p�y]����QZx;�����w)��)�}Bs�5 ��|�2��V���< �����"_έ�����ⷔ�ďE�=��>}5��%;͗�����K{����/��Z�����z'
���]jǠ���T������O��t_*;]Ӌs�+��Y����N
��!@u�%*p�{��	(?dh
+�G���i�I���'6�ey��,�/���/�����Pp4wƾ�8-�����
I��S����i_�KQD[Y���V�������'�L���;��dq�㵋M~yXiz�0v_���|���a�[);,�Q�9�7ȣx�Uf�ԛ.�3>�W-�U�w�<.܁�*�Q~�?���#+U��� bm}����h'4Ya��es�5*1�!"�ϗ�&&��x��������;�dg�%��!l����.6�����<k����!�^y=����u�Z��Ɨ�����[�]z�?����v^:Up����{��$�5���?�Yǲ�:6<Z�#M���!��o�_іbz��9����d��.�x��kZE:��9"�A�r>��[�2�E/D��Fe�}�st"�Ъ�x������f�/E������a
��)첀=���#�T���c��h��f���j���!A>��� �EP�`k� q�6|8%�wc�t��w���;��Т�Kj#��ճ�7�j��1-��8�jm
Ms����%Rx�����ݼm��{�����o[;���/R��	��+3�}�^����eR�]��tZ���Հ� W���~� ]�F�c������X�������SO�"��Se����C�^	7��W�Ao�_x����N��d��<����p����(!Z$"[��q_J6�/��[P�<q)|����[)���>�&+��C��~)�`���Oz��HC#/��	�s�;�Y�q��3�q���#��d�ߣ����u� ?�=��.��2T���"eq?��@��U8�S�q	�xT��`�ZƖK�YO�Q=G�a�^�[O����=J:�tZ&N��{}|)H$Be�0x��Y���5�$��+��P4�ks� ���2i��n�������@Ϣ����I�}����b�X�B�`>_>�4�3�[��\�q��j �GG���:�󟈔bL��$�~��]��7L�Z߻d��y�j��UR�J>��ּ���4������4b{*��EB�E����&rR���9����u��w��Υ�U
�u��^k*�*U�t��:��C�d�%w��ݫ-�N5��O)�����\��W���2�݌!9U
#}�nM�W�#~���j~�ųKѐ.�nr2j�h�A�F�0��&���w2���o����x������3
�]~(�0/:+1��l�?)L�I��'�h��渆����0�)��#�KT�uh��^�;d{b�Y��$�dg1/�ϰ]�[�xU��NV �|Jk=Uч�q}�a@����$cKh%�Mt�[��駁��<����T��CM�x#ޟH�U�n���A�G=a�9���+�l�<Z�ٹ��4D��{J�*N0`��'��мٴ)^�Ϣ)���;��%gl�We���Q+�
w&�w|i�'���A!)��XZ��A�E��k����� �RaN����J�4�9JV�Mú��)D������i;�|����g8֯�u���9�{L7[@(2[D�%�T�SbL%���=$�h�N�c�8��6��8����E��&mɯ�E+(�m�,;f},�{��:��LuȄI]���6<�9��B��E�C�{�6����á;�)�C��0����;[�5��a�ȯ�//�Z�)��5S��t��K����GB_C�YS9:��;�mcB�b�tڽz�*��@M����%�8� w����C�cQW*�3�^�.����ap:l��������K�`���ü��҇�o�SWF������8�f�l9Sqs��M���1Q�3(���G��UV��!�	�j0�������{`ܽ�"���#;�pnb����PV��\+T%�N��w�az�Q-Iwz?��m(s���<�O�j�D����}��y�N8TE��	���)˗�G��JJ�3-��	�[�:'G�t.�]��j�楤����}�N��݌��ej�cq�(n8�K����ۥݲ�w�֍��O�����N,�R�F�!6,u�C���f�V���w���v���i[���8����,d�3f�RM>u%��uDPo
��l�6
�|Ta�����:�7,wk7�Q'�T�jg�.�"[al�T�_���d/斘�����7��#��A�e�lu�!�+��Ot^<��C����GJ�����4\���*�hξ��|ŝ����WP���*z�L)�1KXeH!��~|������qu/M���c��ſ,�e���v�+����\ K�'94h����-�Op��dȈ��Y��ۣ? 4.�]��k������6���g-P�9�a�����4vtF��5Ĉ�H�/k�(��*�ΰ����׽��)�G]i}M$�a��Ҽ�"Ĭ
~{���K�ym����CJ�;/�ܨlÍ���x5߳6+C���7h�P�?�6��"�B2����YP��[!�9����'�#x��ͻx
>��(�[I��9Z��R�(��)w�?����-c}�#�~	�Ǘ`�ϵ��P�8P$5<w��>�{���'Z�P�e7of�xE+c�f�9��?���F ��>��>�<-Z�Q�Q���K?*
[_��u�!B�xɩ�Q�
��)�� ���1��O�f��ͺ�휗����gPg�H?;i?OqӁO�^_~�2�r7�O��Y�Ȑ� A�o��ȭ%�r���a����H\�?�;��U��][࿗�	{�����5D��`�u���������$$.���5��� �s��J����i�����噍���i��^�-.{M�LX�a�m�Gy�(��W6`��.N;��aQn.��-�D���{Y2o���D�\��j�a�)�k�w�fO����ػۢ�.v�,�ީ�Yi�������Vu��YFâ�?��5.��S���^��_5��F�g�6[!���u�ܬ�4��v:M�J�}5��4�T]x�~�#s���vl��awH83k ���[��J.�y������x�5+��4�AR�I�v�m���\��SNJ!��0���C�~-j"���F6��ID���5E|(�z�E?J�SN��p�B.34�������o�FwL�R��Z�i��g66Մ7⛺��hH\����=;Z�x��MI� m��<?���i&���gֈ��i[���� �Gk�,-l�V\!����ͪ���;��{0�+���1��t[��<T+��{.��>!�T���u�9� Eh>Ye�7ཀ�ڡ�8@5ir��
vjg4�����S'��S�J ?���$!J6�=z��~�PGe��?���5��ZV�;�k@�"��:=Kׁ��-�^�L���9��*�۽��z���������:����f��HB^�oтO�)m�m�!$J\�]�f�#Z�̨��2��t�Ԧ��Py�۴�ڈ�*���ԕ��J%(@lv8S�&��
j�`PS����Z����a��.�>�0�� L�w�VŻ���o����d�Qd��k �Y���<�K�a-H�΍^	m2�(`oNxQ�^Ӳ���N�"�^g\��IQ���$��/�]�8��4���B�Qn����o1����Pf�E�>�X#��)���n.�>>g>5��G�%j8�5+_�ӟ�L����u������i����6vX5,���鮶V�9$��N�Yi엽_MUm�5��A� �1��Sݣ�n|Ѭ����w�jA�+���#qx�9�C���!]�C������8�8ST�:���BSC�N��[:1Vj�#�`��w��<��k^�c����2�: %(^�l�C�U8�2��	x=v�T�7�g���KlV�K�juN=��g :[�"��nOa	s��7�?-u����Y��g*���ΰ1��I���L���1Qe(�c��w�%h�"e��ʦr|ù��*�A:1����lv�'|��2�	
���l~V�=?+�#�g��"b^sg'���M16�[����a؞�*�Tb�LD�-��(3lm5C	Y�ۛ�_�.���mQ��"���Ӣn�.�>
+��������\̴t'��D�=��G�-�?��������*�:t��+aX���N�N���H����ۮM"D����%�a����C��U��=Yݼ����'�[Y~�F�3}U�^��E�w$jҕն���U?J���i�<>�������1tY-���l` u�4q�7v]�ޏwHs�nV�\� y:
U#R��M��`�W|�wkMg;���K�rn���6ˤ�M����>P����ǧ���Uu`����v�w����|���\W��c�n(���F?�p�^AHB3<��wzV��ޟV��˦�&�\Q��`ҳ:��l�NT&�6��M#R�@��KI{+2��+�qvL��Т�ֶ�fa0MG� ����9U�W������A�'
eq?J�lVH����`�����SOy��pZ˅���cט�B�x�Chk��`pp�hqR '���ǎ��YH�q���v��r�L���T�C��֢���לӉ4%����/��	B[+'�K�dx�/��g���S-s��F��3���_�/>��15�d��t,�O]�h�wG��&	��	)/��E2��R(��Ru%��s�dgԿ�?|$[��g�278����8�z��Qi�_kܤq��,���#wz�	X�J-�p���!P�ӷ�3	q�PDY�_� ��+Na��.�K�m�)�?��u�=�0W��к���s����k@-������YZ٫n�Ӳ�rj�ۑty�B�ma�X�W�XA���}۹B�>�4���F�	u��*�x"|��)�G�wS��.P�]����ԕ�������ym;)>�3�[���$>R�31*џ|;׻���CYĳ��H�H��>#y%�C��=���mP^ �ҫ�K�.n������_5�z
�Z�F[��c��"�Q�_c��)?�F;Wn(���<�./�g�YfIDߒ'��7x=�SO
">^]j�)n�����e۸}�3�%ܙ$�����Hz�1�K���T<P�� ��B�T�d��L/5�d��e���a.���Ċy�o�T��S(���#��Ƅ�O���!�~��A��c�}�"D�z��@�Y ��l`2@�|��I�j�Ә��zͬ�H��
���4�u&2���/(��nW&�YZJ����q�1�m9�~��>����	��5��(%�R�ysRǲ9wvv�`��;��ц��5�,�HD�Lx�n�B	/���!x�þ7�۽�|c0��UxJ3�.i�O5e���:XܾM�fa�<S�ƴ�2�l�������7!��/���%����o���g���p|d�S�u��c�%�gb�Qp/u�~�\��y�M�g�o"�F)��.ۨ��8�3zp�MoV�JRĳ�eѹ�A�*3����`�� 3�~Ŗ����C|����t�Nv�i�tV+ix)ᵵ�2CV��e��օ�né���u]G~��o��u�Yǒ3�fF�8������=���:���������4���_D�K�	�Tl:r��ĺ}RԻ�oC��h����3������p�%�,�L0����E�D�0���-�HX��pN I`6���*�{�y���w����3QUƔ��S�p�`+�O��m��Y�'��p)^|�G��p_**��d0r���P��N�2��ɡ�S``�ela�G�n���#���R��`����@z��;ӛO=7�1��~����r���>!��&����W�f5'İ
	�q��VE_T�{� ��4���S�A�����;ęp��c"������K��Fe�=�+�� �$����^�v�W�`�>������潊���%K�02�Tu�|�p�Qu�|*�c�3�& F���Ža��m`��`��L�I�qS���`m�iy�*�g�оU��| SP�.*��%�ӳ{9{��1�;��s�j��{�V&�Z+���?k�������A���m��	s)	H
��"j�*QIȿ��;��#�[�Y�4��{�ѧ�W$R@x+We��i4$sn��viD&��v��E~�/�y�$2�~~����|�R�A�_���� |�*���eg�՚��n�,��| ��6*m%�MR���
��$�%q����d�Q(_��⠗�׉Z��۩$&���z+x��N�}���+5rU���u�w�_~�����/Th�*n�9���'�Y���i$w�>�����΃�o�J=����E@��4�wi�?�7�)Z�M�eq�� ��	�!���x`�ax�j�EG��u .�oڒ�˪\�yv�F���N� 	�[`~����E�Қ���1��Y@v�d1�����%�/i�k��?�{�T��kK�mv3֙���F�����7J� s��l���;HGj�7�K��������tʈ�sO�D;�窙8Q�����?�e��D�
�͐7�k:Z�0���|��-G��������@f�~3zA)�O�4a�;Ƕ��!�\�UW.��ej�����9�YǊs|�9��;'U�M������1X	�M/L�]߰�[���o��>������4�)��3��~�O��������HB�5M���,`���bF��H��5����;���IW����=��;:#�>��Q��I��<g��[oP��a�֤4c$�q/��ZS�%-Oe�Z�ƿ�8}��g�t}E�a9,@����M���?�H�Getǎ�{�q��@�ُ{��f����m�wM�6����'� uȚ��"Р����i���w3�7%R͒�[��+��O:7��q�'>#��=��:�d_,4y��J�
�6_�R�I²��T�l��pAʗd�S��.+�}=�)6��7�Y�0h����>��1�&<n�B��qw�iK
<z�&`�v�񔳧�#1lȳ�0yZ\�l�;sI)��.�2BS狽X$r��u��B��a|C����/�����y�[�**ym�����E3�L����h�i�|{�|0��F)Ü��r�P� O��;[�M�흲�i.���*N�qA�L��MHN���|���0n�p��k2+�=��RR�p��v���&s�
FyIq�$�i�Oj�PJ>��Ny�����_�v�2��ۚ��3�>��o 	!�;���*mֽU���
Q�Va���E\[sF�˨�����ub%g�.�����i)<�g2;k��A�������R'����*�m�l	���'PR�jND;<�&�f���󴻧���ʷ��)���Y���񌏹z���٠����#K�mȝvg%�j3MAr�+TW]�CE�B\:�N�}ՀLq��پ#O�{d��k�܏
Pvm�\�f���nn�]ôB�.��g�YƤ"�����K^22�KR���e�8��a�_�w�`N]*�x��j�����D���w7�{`��ʼ�yO��������!���z2����F� ��}�E�Zː���t���Ӱ=�i�n.��2`Y]
r,�6��I����ˠ�d�ѪtuH�.�å����X����;r��d�T�7�wV�{�ӑӻw3����7L��O[�a�'�^��\�s���k��Z>y���mɊ��P�8�+ܷP��� ��6��l���`30`d�5��ߓ�� �#������� ќ�1p��D�_���Nj�\|:��Yz��k_�~���1)���6�������'ꤑU�)�3(�aD��q�g�:X�`�_��u,�-l�� ��iM-�<g:�|�WRp���Eˈ)3�v�`��\l�I'9EM��yM��[^Q;�ha��F<h�G.$U�G���.���8_�ž+��Snj��]=�V����>G|=G��N�k�_��nuT�;k�_j]z��dy�V)^u*Tu�۰�����,_7�a��N#��<عf<�r��� ?�=�Я��_�V�bV�:�u�ir����ä���E�u��� ��Z��?��@ΨP3��0h'@xd�d����l�U������������{ ��ߓ;�s;%�꼢5
}MN�?��=����P[ּ�`tG��/!����}%w��$�N����DO�2ËgD�3z@_[�4���y���jw�Lu�x�ܠ��0�[�8G�$�i�|���=r��爰f��h���vs�hD���.�xWo�Z��#��A���j��{��t�W���U�
�W}!krc6Z��3�ji7���&�V'Fķ[:
8;t���(���x*�:p�J:��V%Y���Q�y�yJ�"���R[f)��U����ј\g1v9r�k��TNQC�hH �v@t�l\�� F6��������I��;n%�n|tT���8�aZc|׎G��Vw�9���c�:Sb�u�KPA�<���d_�f�%�*�a5�����j��k<��������b4���_�΂l��أ�$­�u���3W��5G켊��ރ7�u�/��Q5!1 K˶kj��q�s�G�_���]�����3�e�Pg�A�'T��0��W�
R�W@x_��d�W�*J.T�P��{f`4�2e&����'Y� "��������՟�����t�s�C��������0�Hi_��(��{(A��2�V^Mȿ{��Z��!��޷����A�����g6]�CAJp;5�w��������<Eԃi�b��z� �Jr.jec٥��q�KDbקB����n:"��_������LZ'���v�w����z)�bd{�)�5���N�jg���_p�n��A���x�r<��RE�x��$���z��=��yQMk�����w���@NCi㎮��[:�Os��
�������2�`꫄QF�	=����IC�����s'���j�� |2�ɺ؛�$"D%�E}�ll.����¼0�w�<���6XO��(�-rDQ�=h�s�-v�W_�c�T9�jQT�5�l����O�2�B!v}���Xk��Զ��c�q���_9�+%Y�\t�9P�˪�m�lTI��&�qGL���j���6��¦tDP����ڽ�?��<L:�I�Է�j��oBu���@ ע���?��`�7���k�91@�3Q�Q��y���7�ئ�����+��#�D��4��ƺS�x�A/�@��+c�3���K�F�&��-���O|�(�Ձ�Ҡ��V��"�o1�T$o�jM���E����7�T��Q�c��#���w +T�?`�[���y�C�Z�����Sz��^R҉��?l��	�/I1A?7��Qt��i5��U����%`��㻌��V���q�΄/¦�}}V����{��;�C��J$�������(�e��"e����q�V��d����D��J!�HO�N�'Ա,�̺,ٵ�f14op����*�!�pcF���ŃkyO��UQy��ͮ�F��.��BK��Dl<���>j�cd9+gW5m�"��fl�wK��=��m����Y�ʶ"�
L��\S��I_��rh-�/�b�Fm�S��/.��Wld�{˹�i�~�	��V���=ۺ�X?�Æ����:�L�!3�wj�����*�BK�֬�hRs����e(i���W]Ew@\��������v�|��nZqS�985����1���[�K\(Qĩ�����)�֗�W�X��=��7��m�ˏ�Nq��t�i��k��0eƺ3�&��5��Z���Mf	e#(^�3�H�Z'yk������3��|��bDo�EE��6Ç>=������&��*h ��/�V�`1>ۀرk+�נh4jT�> v�)�b����[�[s���Y!����ogk���ߖ��`�}�z�-~y߫�Ϡ�U��)~��֗4�}��_lYZ�vo��k_3��	^��Ăٳ�N�w�r�t�o"}�-o�d}Ŧ$0�9�0�IMx�9a���䙡�Z��!P� y�+d��4rS$��it�h�Z��7 �,w�Bh��º��w�-�'ڕ��1��:�@�������"���[�5�����9��Z���8��8~ߘ`E�"WV�Sy�����_9�c`W���'����7�S� {�*2��N3�\���֬�SNR܅�������Py���G³<����|e���3!�]��C�
�u�@}_~V��ʯ����KVV|�{sGɈ�?ø7��K���0r��n�Uc��!�1q9GU��35�ӡ��%��#/��>�:}��ْ�.�%7��F:B�ʻi �Mn0Fy#�����ɳ:�sM{�0���������c1��]���GBb�ƨ�[�ϻm1䱔[1�����	<�8�~���on+�E�MU3.����zڮ�8n�3�N5�>n�1�N�Ɓ2#H	����������Cp����i�붥�V�]T���m\*�/����;K��k�u�LV�o��ԜMU'�D�݇5����L�iM��xp� o{Y2jqK�D��X�p���&��(�����?���"�X�,K� QvB��B̖�Y���3j˅+�B�'�TP�+�B�Z�O�C"�L�H�>�` :�U���{�TX��o�H�3_}	�|�nE1���Y�JU���_�`~��w��2{
c7V�`v<��ּ�J����l�(9]�o:1�0��\q��v�_Y�������d޻��J=����s��QW�d�j�k��6�V�e�s�F"��z��/'�ɝ����ŕ�&ↂ.�0֏}���ܴz�r���3�8^�����=�����H�=B�/��@n�9ޘ>�!�e�ޏBG��S'x`Uj�=,��AZ��%E�W:.߫4�et�V���3���)��xW�J%�r��M�P��Z YV��Y-��y�S��	�&.��p�?M�Q��P|i�B�T�/tf�k��>�[.7XG�1y�9�����}���i=��#+u���Z:ߕm/�xZ�D=X��4�v6��i�NU�e���` �b��G��T��ӊ��{W�XQ|^�p:���O�ҹ�-�e�~sҪ�鯸����銱)�Wc.�����X�G$��(�ιCqs��I�<Įj^jd���b�x���wC+�'A������(`����um�o��h�iSՑ�cO�PYt��SdM��>�*:��E��O�f1�s��1�7�^���l�dU���,�\.��G��d3p�f�jڌ�x*[`uJ�S�v��]PM]����L?a������F毠�e�JGU��X����Y����z�mB��zKsӐ�ܸ���JN��!���Q	��'4�[w3��[���e��޽��'�[�_Yj���Xf��7�F���R�(p�q��I���z�����
�v7�i]_7Ae��4�!|f	L�����1Q�}��Y�I�#?O� ���q��׫G��)���i87�0��$W�_;#��R�
z��]�\� �}���ZP�4�������nf��XV�w��)����F>kX��s=�,�9�(�o:{�ӗx����}����"���e�ڇ���C�Όu�S�^r���+O� �~�c��0b1�v@���*�I��7�.6�)c,�S��gR���E��/$D҄ޕi��ێ����3L�߼�wz���E���&jT�f��z���k���KH-6J����W#�S��)(o�$[̚7X
oL|,�s5�Y\O��ܳ�
M�\���b�ύ�a߃�#E=��!���=�)2[����^/9���S���\�c��UF��4�B�'������@u������t&g]rH�I?첤/dG�THm��c'�fԧ�FA���Yd'��-�8��J�2�h�$��h� �#c�Ym#�"B���K=���Ry�"��s�+��p��/�p���b鍄�k�,.��׬����q�g �w)�ї��!Tp�9�t�T���%���^[3'�Wg[�?pAˤ�-���V:Y�b�_�9�lZ��3-�u�M�l"�a��ֽ"��LG�+���͌��?��C��#*��Q��'���w(�P�vܑ���%�U�Z���]M�{�e��[���8�9�7n�����yrW��;���A~���oB�0`A�I��a#��3e�;8Ů�|�t�m�}�	P��>��4����
��J���]�V�R��حѬ+8� n�2�lv��%��oY��y_uY�b�'�;*�"k{E���A�G���������m?/9~�`��J}1�͎$Yv�r(̞�Ң�����f�Y������߉�<C7�@�Q�Xi��,�y9�n��S��p۰���,��f��t*CFS�xK{P�l�#f�>1�2|�鬂�|�A%�)ǂM�S��b�� ��ڂ�
�|�ģ�!���茄�3F�����Ґ#+?���F�u�1Rd�Z;�������;i�Sc�S�.�7�M�r�����g)������O�M�l�oƂB�[�'G�2L;�U0k��5��`��L-m��#X/�2����n�q�����s � �Yh��0�֧8��M���%��`@[+ڽ���j)�K)�g"�2�TܛQ'�Q�8�vz�SR�QdMM���Hu��;۪.K3�����{J%���	��9/���.��ԅ�P�����0�J̲�Kؕ)Dx���萑�Ƙ8�E�'�.��{�H�(����k�x�x�g�����;�s��
ͥ�]��t�f[#�:�]"����6"3��b?"�λ��� 2�)��m��+�F~>K�F�3v0o2�]R�����L�B�ЉɁ�����&
����ܭ���i
����]5\�R���9�0�����KfH��Ս@����u�vP�!	NPU����-�\Z��G� ��:�J���q��
�){r�Q����{p��&�N|�%������m���������;CP		5�gM�U|�O)���<2���4�V<ߟ��W��+�F�t��ޛ�+W�1�!��irNܢ<2�_��+����4�����Q�z�6��d�#��(�S��`2[<D���/��>��|5"9'�M�3������,���f�כuG����:�W�z���Cj�����kb�ɰ����w��۹z��{��ٌ�k�՘�D2�^��"���\[����eL�>���rl�	F�f<kD�m�I������ߞ�oZV�'�f�y��s@�T�mW���@ J�_d��q��i&����sh<�f �u�t�cK�S��i������|z	�� �;簃as�����\R�ztì��Y�t[$G0��.y���YUd+If߉��U�^Jѹ�-�����0���l^�JX�@\�Ǝ�烴��ͳB���a��F���Y��4@��].߼�e2�rdja���Q�3���kr�O?ra�W�9!�V��������\0К�ш�p��d�HGP���JRO|fi��\��4d���b�&2��:�F�	>����U�l�lf�Ȧ߮:�Ca'&7L3]��2�\��E��YQ���NW� zr]4����5 K
Rp�N�/��@�v/��q̸�.�����Z�Gc�<W���?��eJ_�/��ܰ^�ǰM����{:x[�����~�N��X�\	
��ݔ�:�!j�ƕ�^Z9|��1l �� &G�*�6Dt�$��p��@Y��-*0�犲�HSg�&���7~������	��/���!��s��PuHu��ϙ�й��B�+���|�!Í��C��T۲l�z~���f Mcz�<} �ݿ�+��>�#�+��q&,�)������R�R�4�9�ݽ�jV"�{'̆����m7�'����){�O�.7�;�-�J�܆��y/�+���L�aE1f%O�[7�d������!9e�O����/�E���W��F�ީFT�`O]��^�S�]�TA�*+��N#hD��]��"�!�e�9�.�l�Fy��n,_��!������əOi�W���M�u[Q\���K��n]ۚͰ�s��S�gEev�#������졚���Y��BW>L���o���9\У�-�>A�Z9�=h�ͪa%�����Lg����F앥�0ٳ�^���9]�5�~�TV�x�4`�!>�se5�0�|-�nσ�����2-gX��%H�dܖ�TەZl�tY�-��D��v���қz œ��`�/
 ��J+(�I��Gx2)5�4�8~��n�!�����5�"����<���}cFWܧ:�1:N~����=cqfo����0� ��z�S1+q�Y�H�ל�{\�i5'��;Af���������I��&�n�V$SRh���)�tV�qtr3�j]�tuN�*vyy�Zf��� ��.;X�Q~��E��5~������yp�J��J������c���2�z&�E$�7G0��[j �g�#��N�vҾ�ϊg�t%V��oZI]I�UK�Y4oL���N���I8\<~1����?�"3%�˦l�)f��?���D����ȄO�/z���KD	�6� kf��8o/�`�0~�$m���V�׷�Hm��Ծ�Z�����׏:�,�/k��������y�v��%.���	j���c��XhE��o��I���+�����M�?,۲g֙�w�e�Y`S[J����?�N��|):Y>�����|S��m"�!��7g�V��m U件�����?���LGP&��STۙ�ڵq�\F�k�>��?��"Zt��ѶE,\�~�*�u�h��'k�!�p6��sݒtX��޴��(9�8M�WB<�5���d��s�Mkr���Sm�/�f���nv��8��Cp6��,�N�����Kk�Bs�W�F�L��"il���1C@b��ŵ��8
� g�����i��� �ٍU��)����bb�H���Xuxn��H��>�w٣lo9r�� Qz��sl��PX$�`�MMӊqu��Z�3)5�К����= �I�H����-F%@+��7�pp����O�n�}�h"���{�<B$���<x�z=�u�1�/��呩���thu�W�8A0;��~�>�e�х^��j�����X�y|7c��e��@�K��F飯������J$��x�}�[o�������E,�AQQ�nP)��&!#�:d�ҝ#6%��5Bb�6r�����}���8��s��y��޻��L�po��#�M��"��#_BR��_u�kϫ�Ϸ7J�(ǽu4�^�y_�.�2|Oe�ǵ��/��E�W�`͇hlW�Ȉ�M��~XJ����1Wb*��qR�}�\��@\���\����Z퍆��nj�ԉڥ+U��Nu�c���Ch����!极�8�bƘ�����8 ��fζɃ�����ʋ���Ƀ�G�ubU+�G�8r�H���QS�����h�{k�k�O�?�?ZX��H%�����|Z��H�k�	�d)dF���SI��2$����!	� +�ke�����V�7|���	>ȍ}BL���%��o�{�6q:C���A����5��<H��c��rȜ`v����琯�̠��9�~y)���?��q4h�ˆ�I�/ӽ�J��z�Ǭ��7�4^6`Yf�n����(�[s��<�k��Ik��!쐶ͣ*u|�N�ڝ)2�r�"�N�����;W��tl?�;�6۩�SⅬK�vNC���=Q0�J�q�K-6�q�`:��W�����~�@��sJ$n��话�9`��4�C`c�J�QC�6գdo8�%���D᯻����[�3�J���Ux���G/�̚�8��In!J�D��s�y:E�?��>�I�_����v��tx�z�S���lu�Y��S@�4��Z�%�B����:�����mt�ʧ"l�X�����N��,39�S��L��� �%���=�@�+W�)&��rD�ڸ�9}ϦR������?R�H��u� �i>x;�)�'MB�zB�E�..�.���;ƚK���[�SG?ɼe�46թ��� y�G�ߖ�˳N�ћ���<�~ƉC\4k�1�Q%���! ���^��$����ɆL0�
*M"#�8����gG�-�:d�j�����������Ⱥ�����M_7���냷:R����5w>7J��%3	[�.fL�?Ѳ�I?�YJӈ�
ήb���S��[�5l���2�}<f0� �ͯ����B�Yr���p�]�S�74�٫BB�E�Yū�M]=a8#`�ekv�|�&�'d��9�P�1�BN�n����@�V�ѩΓ����V�i$Ef���;7�w�_��W������ T	b
�1�ݚ�|��	�J��eUi��Bi����B��N�|�(���->���ŕ_�+��c�w��fE�+�S,�'xLڮ\�����r�/S��n�|t��im'���;d��R?K9��N��W�-	ׁS�6�P�n�y/�ʗ��Zc�Y�=1 �Dt�Ovs"U�̃����6�궗��	�,�\&�r�o퇯 �uF�9��H��pM��)8�j3�ԇ��]��z�Ss;��X4J�HM�sQ�S�bcC� FՉ��-�R��ᨄ%��!�T�S�?�>�Qmb���F�5+�Ӟ�T��<
�c��B��\�jH�|4�k���o��館?;�ψ��0["7O�y"7��/�@3�7Ȧ�rb8U/�.�{y�z϶lENI�R��g��~Q���v(B���Y�m��m���,�D
r\∯����'�z.����;}�5�lQ��L�����s����!j����\�9�t�\	3�ie����������j����5�5Ե��F���Yc���d��*�t;Ƣ�Y]�?���*n:�����p����%�)��'!F���U��p�/3%F�o������.��c�N`gZX�nR�lfvnU$pYD0/�V\??�;���S��p+ؾpaJ�j9@�>jes���6�A�d��Юu�iHG����OD�T#��[bCg4F�&͘�U�G�2�5�L��-�"��*��m���Ut�틫�����Ix�se�SD�*�N1�8�i�:��R�]�Q�3� 1\Nb�bc+{�WX1�"g_�~&]?<ܚΔT��B!FS��*.�y<t�.�~ޟФSj���Cs���p�祝�QApNJf1 ��Xm!%#Ο&R������8M��kdDF�qT|��f���ŋ�����\�@@������h��*Y�9�G�8ŷ&�y� �+'n����L�J/�X~y{5�Q����"wD�u���tJ��I�pg� pD*�!�G�{d��d��Lв���"rI�����wg�K-� ��o���f$� 9NDo4�p���%������H�G���_�/"Rv�-HY��v�÷P�aX�Uv$��&�@�>��79�_5��B#3����Ő�/}�FQ���"�e��><�T�e�v�|�r��L�J�C��(ֿ���(��~�����,j���Ҫd? 7�w�0�:l�R��WrO�̢jw2�;�U��\���G2�z�&C_Ԗ;�d�d�q�a���w�a{P*�~�t��:=�	~ �o���zTN��~��w9�@v���Y&Tυ�ߚ����Z����~"Z)��\�	B�6����r{T���O�Җ~)9p"��@@z�$��U��@oURH���~��N������^?��y�F��Χ�'��=���*{���/k@�s�h�{3u�E.R\�����}Y��n����0A2"�p�f�w��R��[Y�*��r�s*�^Q������hO�K��J!x�r�@pc?S!f�^-�4dD�+�GDD���K��(~�:p�W_�#H�s�0ǡs�i�g�؁��o[��+�u��C�h��:���\&�[����kY�ҿ�18*����[bp+�+����vq�|�:���8b�)����M	�DQ���A˒�s��J�j���˄�w�����;#�Uդ�ճ�G�}�aY��C��H8��9���и�_M9~is5p��@OAE(�+����rMZ�CZ�����g��?ǯ�|���rCM��^WPA`���7�`�!��{.��,I����L�L�L^J~�L\_Q�MnMʙ�������ĺ��Wz�򉇔�#ǝ��,c���o�Cv�s_������k{�MK��P�>�����h�h�	G�:�+9�~5l�#_���}�~H+n��7i`V�mm�ep#گ�L�(	H��J���ɟ[pt-u���� �!qY�z���lU��]܋w6u}��e�>>��������l�$��ex���?�o)WO�S�<��HF��t�۱�$�旡��m�R��׍F�Z���~�x�7�?�@&%��r4���V��iur\���PF��u�x�P�����{�F'������JI�3�G`:�w�f3=�@�E��%M�j��UՌ��������9� 3����haTNڏF��9�<�RS�3������%^w���/���Ì��x���X}��ʬBS�*,�(,����̔�$�
�7���ϴ�n�V3��|�G�\)ܓ%l�h���O��D�9�?���Q��8J���-@<���7`�7�b`��`ݰ���F?4-Tn�g����(}4����� ����7�ʂ9�{\��<������	y���m\�ۥ1�F\��W������z�2+\MPe�����--�f�U�X����J�W��,���U���w~.B����~_���V�;o̾��d����xC��3/����r���4�h�k-O5��&��5���h�I7��J���n�����!��mkv["���^��|j�"�GC �w��Y�u���I����T��C9��l;�k��{K�<�[>���|��R3~�Z��=�j)�c���_���G����2Q������?���MF&���'iH�m҇k��݄�c.϶���-��/�k�-���v�\y&�y�� ��~�1ۚ��
ƟB����>��� �!o#DH�-=��>|�V��#��8��i���G��o8�O)��J�v��{��R�[�%�y�:/gWX� {.��p,���Y��z�4u�ca"���]C�Vwed���Le�#U�Y�G.u1o��|���1���ˠD�� J�*�?�eM�_��	�o�U=��,A�:�c�O���l)�����<E��HW����\�O`.,r�Y����ϵ �C'35a%��/��I$���/����꟮����n	���u�Nc�,���"ot|#6��&�7�W��W�s�âT����DH�}$vM^&X���P���)h��IO�o�l���4�ܰ�&BP\��uw�u(؁��LknBZ���Hqd����Jx#|�8�;�KIB�HX�wܜh�{!�,�	���ԣ�v�x����U&�(���t<H.C|^�	�������^S��tޟ������F-b�'��m��N����Ph$�K'�̿0��1�/HS3]�t$U�/�]��|
��7�e��ل�®�T��,��U�ڳ0�G�N�92��'�M�' 0��Lk�T�4�]��j���&�߼�W���B��o�k���.��!��Z�#���Р���/�Hp��m�����'/�}E~����t�ooBʈ����3�&���X�Uv~�8�h��T�t��e%���؀�����A��	�٪]�y95��g&W��U�j���0��@��şjTe��cìG���o�7)Q-�ؗL2?��}�=�PxF�&2ٲ�q
u9��m2�^��+2����k�ը�����^�P�������^�otޱ�� ��|:�]�4f�$ nrg�3F�)�*
�b^Ec��s�Yf+�
�Lε�����T�8w���+�P=���	����K6`U��׉Y�-��7k��=�����~nq�z1�K�����4�N�c��o�3�JC2_��ϔ����"FF�ƶ-E%����ְ:�����Δ��= c�1۲�8vJ⛥ii0>v���&�7��7����;�e���O��v�a�r+�B��\��Si�������R�������:YB9 @F�B� ���%y3���C��Nx<�x�Op�~ �9��{o2��R�kf�V��B�۵� ��,�8E`v4r���f����qX��)���Q�%Wa�����ŚF�pRR�X4@�t�ԅ�7�Dn9-�E8�n*g���v���Vw-������V�̢�̋;��4��"x���aY�6��L>���t���[En>�oPv{v��Qnv̠�q���,�\vC��^d��ZtJ&ǝ�w��]xgC���ٷ��?6*�vs����j��6���q������:�5��F��D�Y�0��ʭ�`B7횄���-�G���d����]����p���,a��8�����/4�!��2��Z�����!w�$�O�����M�)�4]��{� ����ɔʉM������'z\@�t��M��=�],���h��Gr�s%ݜLvu<"Z�(^c�3[��i^f��px���U惀�O��+`8ʗul,�y7�6� "�C�r����cN#�b(ZJ���$����[�l���;7��v!��/��y�n��ն�K.1_���Qʃy�Rw�����R�J�\�����O:��iI��[(@Ë���0��ĂNk=M��Ѵ�Y<���Ľ��9m��b>��L�{���U�!��)����$�������T�J(�u`y��Xm�(���v�6f}N���4?@�Z�=j��B?��ضB�����A��X��v��+���}?��H�"�P�#sI�/rS���F9Ъ�}#��LhM�hs�)>���f^~�(�T#[��#�}C�=��~&|_�:>Zjkp����H�/|l�}�U:K�bd��9Qu?�0��5r�;�P�H��"�USR���}���
���<�LE!�79�#��15��`\dq3�����"T�%��4�����I���<���J�Y�^}��#����0�%Y���Pf��@�2��GtA&f��M69-�}���}h��P�+e5���6�e�Y�#�lj�J�RS�e�d(�Vd��ϢH�d�8[6zp��w4&���1�_��?n��_?�4�9"ZA���B�������p��F��-��UR��(�̦�0��ڪ��y�F9�+w���= ���yy��I:�֬4��dqR���!gwu����6ã� x����l��2x}8��ܷJ��m��[����"W5��F<r�#��0i��FN�l��+G��7V�m��va�)¯�T�N;�fz�-�_�VK���ʵ��V�r+�F1�GC �b�	�4���D���Pt.aC���b�Ǡ� 9d��È�n�_��Z�������6�=*9;��	��o�2Ί ��i�9Id]S�6��\T?���ea��Zh�e�m��9�W-��t�L���o4����B]f�B���eQ�[�M2"�'�R�Rqgל���%�����j%򵴎�6Wov� Nx��q�"�f�:�v�ʭ:�u�Xi�K����a�C5�):��T��O������]-)F�"9I�'���2�b�;ƄL����ߡ�^��I��V;��5�BEf��%;.����TNT�n{Q;V ������@�e�#M����N��(;b���eU��7�49wr��#XAs����nٓ󺎗���R����pKAR�Y�i��[�K�K�! �����Čs	A��������p��r�\pS�~�����j�����N��X��ȪN�����ڳ)�_�
A�c� VE��fY=��iE�O�59�C^�0?��'�S�r�6o�d�?�G:�H�)5i�W�����[^&�89����x]�/[0�<�S̒�߸-+OU��\^wh����Z�{�}8y�����y�K�]���m��:�J�URB"Ap�^]l7�3ߗ/��l��P���3'\�������7��\۬�v�~���2��g��`c9̷�]i�J�>k�&�Se���+�*=��KN�8��hZ3.�6��&�n�]��b��J���z�c��/��N����?F��C�ٺ���1�|y�_ܜ�|64}
����r���>(�E���	+��o�V�v�Dqo���28����?��{�у�\�׹TM�Γ��}z��>V�i�aX~�$��w����Ss�^��L�߭u����!-���߆iDvj�W�M�W�ǁ2�S����Ž_�I���
®�5�O~z��_9X� �O�n4�կ� X�\� �EnoU��K���3���m ɴ���xǁ��=��:�ʶ�2 '���S��!y��,��N�a�maU�1JO5�f�Pؙ�p�\�-�ֆ��mH���kͱ�>C����yռz��V�z{�sd�{��49�iL��? �Ku �i�|��9���r����|���@$W4)<�ݴ;f6�:�����|��e�=;�ȥ���[��E#.��lo�{H��WO!�[eJ���-�e:2"ͬu<5��Ǜ���Y�\��>i?~?���po�n���Ї��C>�%�_���h��{�󝍮�Kb���/� JAs����G@��0!�k���Jnf۸����{o���ع!l��V�{���}4���H����*N����΀L)0���c�7/�<��2��(eR���UWb��O�h��{3�a��[+�l����6�N�5cShX�d2؎���ZQM58���]�}�D~���%����S��ɛ­�pe;�W��9��6�������_ɒ�0I�K���V�h\T:j �E6o�i 9=I|�.0h.ۺ�^c��`tf#�bBI�x=��������a�P�y��lM�s<����E���{&r\��=��*��9�N����N�y�o��ZVd[3�[[m�:��p����N/(�c�Z��p	�d�|U��:�:"�I~�J��Ǩ��3����/=F��JV^�>M�����IPq^���6�5C0q����&t����T�_�����5�1�O`���kwz_�2Ɖ�_�F��Jn���L�����M�L�s��݊�#XcAo��h�j��/0�(A|�_�j^�:{Lʚd�z�r�,�(}��bo~���ね�Ge�o��r�{4����k-�jqs4���T8j�g�;�=im[��t��}��d���v�p����zu����8ҰMҢ���Hz�߷�%眳��Q���/�<n/��Ҁ9	�M_��}˯>C����M��t���W��<�^���Pu&(��7��p#;�{�唦^R~/g-�l��^� ȯ�N��927g=���F�N�ӳ��R���[@o��ª���K��B��:*;��u��<2��1VG�(��Ŭ_�5,C��T���~6Ee2�����p8����ٺT��^.������K;`$j9!h�ѐ%������\@���P�,"��VW���۸�B�th�}��H' �K�;����N��:o�'��?w<X}�t_�a��]����u_�P����*bL�E��2�Z\�N?Z�8����/Ff+����
$�O�"����Z�IE��zi�P�z�z�6��O0��'��/H�k[<�x��Ŗ)�1	G`���^��qd&0��72I(���X���h 0�6	'�|����F�oB8~VDJ[�#�p��6z�3�h���O��O J1��'h�*��@f�x�u;��@�I�|[�C\?�/Cձ"Ԥ�Hͫ/7����k��"FK�n��W�J�C=
�3gTTj,fNM*������8Ko����gW^<g�Nݹaxj�"-�j���
O�x�5^��|o
'h�G��^4ى��L%t�_���%"��hSȑ�ϔ��������T`���.U���0�"I~�Hܵd�z����1l&��j���W�[��{��-I5.b�l.����j�֯>V~"���3�8�ȏ�✥}լ.�3aP-ˈS�|��y���T�Lo2���t��@ܼp�a��2+�1�L���З������0}>��(�M�3ɩJ�����A��78~�A._0*�t9�#*`�S����N�/V���#��d-W`7,^��2���}�c~>C���T�}{���>7`���� ����=�s��BI*QNa��l3/��jN���@Ff7�ٷ銭�w���_F3��D!IE�E�.��>a�g��) �e�2���[���R�wӽ��>�fY���<g��z���߼V�Ni!*l�6�t,AƪeͲSc�C��~��f���պ�����6*<�6�'ɨZ�r���Ő�]@�Y֎	g�Q숰{ �V*,V�3x���`#Z���wyN��m��>P�[@#��Zŭ�[��R�f�+L�;�Ti�:2|��� M��/�|�!U�g�M��_�-�\����I������i�?1u�ʢ>͍l �r⨾־��%�S�^[���_4G����Zz�y�;��ka���3}����Ȭbh$hQ�Yq��L��ei B�sK9������E�=�V{��o>-�
� ���F�l_v�o���ž�m�A�c�k�\�%�.c.�m�X"�� �>��A%��H�	�;sb7�^`y�I�jyZg��2���(xΝ����Y�p\H@9��=٧L�xϗٞ�3�_V̩��ه���%���|z\1Y��s�<��x��g��_��}�}���t� ������ߔl�671��P�� �����v��xO���D�5��r�;Ǆ~!rc�8߻=!��U���H8��̝����ͱ�Ά���te�7�F,�,������}���o�V�]��s�-��;pc�n)ŬH��*�����xX@�wn߸��*��=`���%��C)b���32�x��}�����y�{���<\�2-Y@�R�`����i�V��5ĉ��=��ޓ�Ϥ�SF��l{\��G����o0�*�����Vƚ��&f�R��t��P��1��D��������;�(�+�+n�)aYf$����wn�l�tރz*��(��	����_]a�a��H�9��-{l�Ȕ�'�:�>T~� a٪H�.������&w���12%x���m�����ÔA�,ȨZ���&b��_Dr�=���MD�� ޫ�+ºp�����0�m��ul*��ꚹhhPP�Il��EN>���a�Vg>��쪌�?��������I��5�A}��f�Pv��m�i�uwܡB_��I�C9�5`�*ﯡ)�m���ŀ��Ï�������x�N���KL������%\z��qF#���N=S�6��z����s��r��d,�H,m8s���I|z���$��|���޹]��q�+A�����5�i�:x:2"F����P�l5�I�ǵ@^���З\0ۜ�p�,}J٩�qM�K�
P`ԃ߲4%]�Ox���繉��%N����ҏtm��<��+��[ps{�ȷ,� I�Gx��3(%�%`��
=�c��4# �!�e�������6_c!�=�y�Se�$r�k�'oO"���
�+Q&D�^Q����xM�7�Ĵc����ODc�a���D�������b�H���;�8�!���@�H�6�]?do��g� ʌ_���pih�$`����:!=���A~�o�	)��QET�7�v���<��E��U ��V��_���{؍M��5-̅c�ܑ:�� qώɠ87`棙�WD؅�Ua�U���R8F%��w՛��q%\����++j��]��
l�R��N��ӗ<�W���]TsK� ���?ʎ��=�X�l�&U�]/�MjH�'�
�"&F9@�p�����8°)�h�P��J~Q�L^�7����6o�/�r\-a��(0D���� l���۞���ݕ�wk�H6�!��3�=����D�V���c��p���ᕈ��G�L�����ŃrmJ:�>��/��N��X{9W�.4]O���2S��t��6<��t��qNF͞[Q#��-���ޕsD��D��U�Z�d4W��_s�W]�N�|��)� |�8���u[Y=
���S(&���Ig\��F9�:��G�SՂ�Q�(�K���5=��k����z_�E_�����&�#��C��XT1[��/c�*n�������7J{I��n�ulP�,��F,��OJ��݆;��[��x/y���E�J�_)�{���+ �al�=ʱ�O��(i�_�����S�bi�q�Y��[������g�We�Wn�������`��.
����`�P�M�h�o�,�'��w�Wl��NS�� �]�|dp?]�����H���;�k�$���i��D9�yĚ������/����c��5Ҧ���F�C$�k�zѧ��#�5Sݪa;-��TK�WW�BmNt��e`�?����}����#e��5�p/Xsh���O��V�[���s���Pcp�7��8��A���J��R�9�#���0�ۣ��s=��b�,��UTZ����@6|"_ ��'6$�mv�8��e�i�w5K��*B�f;�]��Y���@��[{�d�	B�V�%ڠ�U����m���^o-TNl���	@����p�V!̘W��5�i��d�?��A���}F)?2�bJ�:��[�2!\X�Nr��劉�n�`VO�*��/�U=Q,�C�J-č4����0|�OH�v{M��jh򆇎3�]�����ӻŇ��x0�pW!q�u|[w�a=X���+vS[9�Wž�xcjF���	�������а�Z�y�nEe�Mۙ���฾�O	q�ps��x�I�i�#�v^����M��U�E|��j�x�Q�����1���MI^K;;����z���4�Cr��މ��:��<qx��|�^(�Z�,;h�jĀ:u2���s8M��"s&L$r?KZ��:�Zak�ZQ�<~���s#S����'�"d��ޅ\î�;�!�롂��0Rf�x�Bf��_�c��D�vMFM����ťQ_����m*�7@9G��=��[
++:�v$�~�)�D�~�zim-�����M�Կ�yH�d���6���2S���uC"��5���*vξ=��G�N���&��T�\~��mI%���''gǭ�o�:ȳ"�ȷa�~���Ο-,�ޚ��pJG7��3���|Eo��6��g�<���2�M\^}�mx���<���<��ہ#0"W��v���{�Բ�V?��X#z?����Q<�*�C�^�}��͆(U:�k"�;Q��8g�>���Bo5<ΖL|3)j�r8���k���L�Sp��u���4�U?���. ���$�p�'��\��M_o�[G�ס~�F�!�8�o����{AX��b�|0�)�+PLq̘�ۄ� ��W�JC���P�.Nw��cÕ�[)R������#j3;��|�jHǪ��#}��_����_���p��� g���|�n_��q����X#1�U������;���u3$		��&u��.x�G���uQ���Q�M�j����D[X�����K�l��(�;�F�&)ɫCU�i���˫�6��j)Ш7��$Ie-fQ�<&��;�6n��佪�zM�Z��?4h�fB�{��z%f�Y���~�F[$���R^g�<>����|���-?�t�2�J���mJ����h�K&��J�|�0��b��7�y��k�`}1�f��N�6\��!,Ck��ŭ�H�t�T��<���=m���:;�>Q�D~9�]�0&+���3������;�ڷ��փ޲�İc�G�)�WA�����+c3��p��2�GnoJu/�>�s
x�ђ��iwἰRV��D���p�p���D�/�\��:�&y}�y�c �1�c��%s�uثХj� �E�E\2k��]qܓ;�TU��/������;��i��E�6�/�-y��ɵn�B��wy��?��� ,�He�ٝw\�ϩ���z�g9X�&���\��uKUYb�ǯ|v��1�57�o�;2r���M��t��ޑ���K�nN,n���~Jva�ټ'~��C���(J�H`�L�}�tL�:��!�k|I�Oj�j-a���`Õ9����4^��3|3&��j���0='�ѥ-�y��(��ZH
���4��?=�g�ũ�/�.a���5.�@,I�"q��((#^W݃��y�/�4�@|0��(t�m����{f��e�%6``؀k��u�R3�N5`x��\|d�8�]�C"�K�u��؉T���ݎ��{aϘ6`r��W��$�F�Ϋ����'i0K=��A8e�^J�H""V��1��2�/R H�Q�YWO<>Z�d7`��_�
�yƃʗ�DV~
-W+9r�C�0=��[����tf�>j���q:A�]r��{���������3�����Ȓ0���j<~�v=O�z�3{��x�����{�`I���M�Zu�+"7_�����>9��~�`s�d���_�������죝�D�qII�]
�?Q�n��,��KG����.[����?�i��oT�:�+��-w؟��"�ȡ�{?�]������v}��zDҡ������~t�'g�P�k{m���#'M���k���4$
��å�>)���q2`g�/	��o!�.���Ve��0���Ua�`�	�Q�IC��s��)�UĐx��"y�Q�(O3!h���ȿ%Oh×�?�����T8�����'�-�$������9��V'Hr��������[�ј�j���� jj�#V������<)ZP��m3��9���8����qi�)��1�����s���w�X�͆�[α|���N��>0�+����m^���cՐ�"rg�;��6�'�~�P<�����O�.Ь�Cӹ�"��^f�>J6����;�É!'o��~OdaU�@n�����(GXq��Me��&x|9��Xw��N�~���?�G.�,�z�et����*��sP��tk�W�xǠ���s��ږ�8�ZE�&�s-�3�up�Y�?��63�p�ٞA{K_�_�@�w�lNMi���=y|�]��=q���W���{�E|/������j\�+�͏�l��׍j�&;�/�)�ڪ��'��,z>H,V����Ik�����-��OWp=�36%T"�[V�h*�l��8�D�R{��ÜM�@mTc|�c�D��{8�w���t3G�
�f�A}��?�<\���$��������]��i�P�c�$��_��O����j8٪1�^|o���)� U���^��7.R��>4������f�X�������T�-��Z�'�&1��;���ɘSN�x�W]���>��;��z�a�_6.8���>�:���a����d��OW�6=��3��
e�D�K]��������98 m@hb �x��Ѻ�u3l�ְk�/# % ��U������Ӓj�Ǽ�4"w��@�N�����XuU��a���F�:�#�au#���Ou��K<Y�?���5�|H5ݰo��N}wK�U��L����B�t��Ɂ����j�����p�P��A���P)���'eB�[����O>5���QI��>���5�o��x_+C�pB[y��/��Oϰ�52�,�7E㼞��%�����^��;iݕ�(�+�H�w�T���K6m����UTlyM'�p	�+$3ݘQ�}���\���ږn.��y�ʈ���g�w�f�N: 9p%�f�3�,>�~���y�1�Ș��D4�'�ߴ����_��-�`�8���p����:�H��gI	��GO��H%
 Qw������n|�ӹ׊���L��Wr'���<�J"�d/`1�+a{�]/���B�)b���>#�k#�*Š36O���8T�n����e�����έ�(�W�S��5�mR��7t��x�� ���J�v��m҃�u�8U���wIGG�!��g�_Rx"�Oc�\X!�BE�f������F'��˩ec�@���a�ZL`����,���;��c�R9Y6j�ʾ޷����mR�������2�����RGL~�:������)ͤ��\5E��p!fR�I%�sNAv���Á�c�|#>��y��K%@T�!�\��>p?�\3���f���[,��������=�r�dn7�R��R(�O��EOl|X��ez|��Фwt��Q��ɽ@��8_l�u?�Bp�?+g����"7G  ���޹+4B�9��N�J0�j��W<�t"5�Zճ?F)ޏ�z��{���~����A)����J������b��\̈́	�4>�Ne�����	��|p�k��{'8ݵJ;^���j�:~�ȃ�23پ� �>����Z���-~>=Y܆����H;�����V[Y磌�iu����IIo>���=~E��(M���"���[�j$TkD�:lݠ��2��5s��X����苯(dz�OSYl��S�xV&��n�������;Ɣ5qh���<�nXײ��e}�pƉ�埔�c,Xv���ԗ~�%���)A)��U]�;)�5��σ�9e�[�T;�V��,
�A�nqi��CW^� �`vy���U���kw=�e=�m��G�lִ�B��n]�[G������{�aV�FM'���r�WWQ(���_m�����lPk����!���+����,����<��Uc�L`�1�����[��u�q"���_�ƈ��>�!鋆�+S}�=�"n��H��F��1�[��t�?p�Aٞ��Q���s��9�v�aR�6`.NY��Z�S^��U�8���hLby����d��bjQ�O>���45H��]O1(�mаZ!E�:t�18\��ؚ/��Qے�P�KEF�e{��}y�?�ȹ�su:7�>~�7�%���K�W��L��Ν��9>�8{gYe��ǔ�ؼ���W�۪!4�^�Eu�1�P�a�T�2�N7'���D{�S�J%߱�����P��6����\�(�+ݍ�S��7,�-�L�{�@Y��i��nk,��b�j&V�����[�V�{���|���[�����5w���=�
�` �h�(M����Q;Fu9�$!�҇�f)/�T�@�o��doǲ�8� XO4߇`H,l�a#}ױq�"e[�4�^"��b��]��a��M����)�T��iT�dK��?�;���8��};|HD=Y
HM�1=�7���f�b#%���i
�";�)+"�p�%� �gt�|2���Pdh^��ԁ��q�x�����,o�cm��S�XPc��F�}�~��/S�wҘ2��:�#�Mz���`�(�������,�q�������|����%Z�9��)��vq�K�����\/O����O}�_���M	$*���[����������?<���6�bŘ�A�eo�1"�+��Ēj��#��[�GQE�ͺ=�-@��o����~���;�LO�J�V����)wL�r�K`0�,rR�7s�ȳ;y�@G#!�l&��?�_B�1	-����-�q;�,��P��)�ii)E�-ڱT �p�O��o�U�Y�G��j�!��ڥ�;���Mzz�-��)�����*����|F�@g�����������RqR��ޤ����*���1�pE����9�� h��!x�G���K�p���}�|8�ۋ#䐦��G{����Y&�a<C�U�|�ð��b@��'�<�8�鲈e�v�VI��)��?�}�ks��m��bU���z�=Wm�Cj��u�5"�}�'�y�%��*	�'��p"O���}S�u?��Dƞ��d�3�H)%��B�Y)-�~�߻�/����W������_d���o\wptX�7�r���q73܂�h�};2�$eK|	��UuY��.�y���:������,�iqWxg�I��+V�����m�#1�x'���7�#�(�
j"q��V��нx÷�P��
��i���ix	�70:���'2�{�2h�&1�c�[�0�E`N&�6ְ�?j�앉��hxǈw�J$£���c'�m�>0iTgQ��%�Z�z7��T=:I?�����{uO�X�0za9��:�凿%��p�Ja>�#�I����8��n�6"n�����	vl���K5�*5ty/�-yrA�ܪ�Tc�[�#ñ�5��q��q��N��3��P �Y�F��+�z�Κg����3ˣ����K+&����S�s��ḣ��2�V%�IV|e� �l�s�ܻ�06y,�[��U0����Ыe��yE���Q�nJ�!��30x��u��.�����ީ��_�Z|���P�QQ��� � �R"�-�4J(J!�0tI*%%H���0�ЍHI�C��}~�^_���s���=j�5(��.������(\c5^SF&&w�*��"�/#�6�o����(��f�^�Չ�00v�lОE�}��a����������S���L��5zX��Г�^=�F�|l��+�#j�����$!b:2gџ;��P+�1�4{�%�mkrk�WF�iT�N�*��Nb�ٶs]�s�����cBX��_�}�xv��9�W8��Z\|��Ml8h��qϭ��{�l�팪2w�#�&�|񿞺�z؅�2�:|�?= >�D	uĠ:�8|t���7Ζ��Z2�ٶ���W�3 �۴V,HN�bw�����Z�P���	u;:�l�я/�7��!�h�a'u�'^#m��Gr����=Wj�.��s$3���L���eb����\���Se�h��Y�cO�1tl&�Yqr��^he���s!b�A /�N�)��e�5�>mk��$a�P}�ֲ��/drO�"T:�"����<c]4�?K99#ј�z�)c��hi,�ơ��-JN���R����q����(�1�8}�;Ъ3�O��\	Z#��1d�	e�s�ݪL��mݬ�m��^�	�#�,��1���+ ��!�5\n>곑��S�34i�.}�%�����콱w'8%W$łe�v�&t���7�3\��5�}aL�Ò�@I�!?�Yt(N�p޺,Wq�?���a�{Il�Q�]L�����>-���f�T�/;��u$3�)����~�k�=��pV�7Z9	�d�u���s�#[>!���P[�m=�r��F����T�S��ӶMW_ϙ��I��a|q��o�'�̹ٵ�I��4Q�;cJ��7k��u�B$�M*yV���U��U#�P�ϧ���L��.��pIi��C:��[~��9 ڇ��[���,��V�s����}��l��r�v����;�F�L�Ui���9L�Ϲ5#� ��8���~�����y�Sѿ$V߅��	�l�Mg��{`/š�A�rX�㮳��tx_�Z���R��'�~��l�S���TCk�_�)v����sĬ���E1��M��u��}������A�� ?����[Φ��Vͣ�oF��^����{�,5/;���x´f����O����o�X��*�O��g"QL�������gK����1<�ױ����s��I#�r���NOڈ�4��*�;1���@������l�%�{cm�4�<�<�}F�~}�� t�qQ�B���&&u5
1Û�X���ف���Q��PW��B��T�����#>��(�P["^:���1+�G�4�F�������&P�zQ/�p�=����M��;3���Vûi��:/�;���v����A�h��VKC�%�9J�C�V�����+sg��c;�/��#��{�A�Śih�]��-��o\C�����KN��'��F���?�����2�ly9\�������w�'���3�$o�f;@˭Em\>�]V=�﹵����A�;�b㓸m��ڲ�\d׆�S(��l^�yfo��7n	�8� ���
`ڗ��R����[Ӏ��*��ο	y(�ld�������N�Փ�/����{�>�8��^|8}$=�v�'�"�Mj�@��b,�EL�nI�Pi����x��On*fM~���(���Z����K�qv7��~ǹ;��gn|krU,�<�/�[�5o��;�O��}M"�Q���nw�a">���l��t�x�>�bC��G��Z�U�\��s�����k�����͜?��~�!��i��g>��K�r���:F&^�[B�2�7��54
�	�i����J	8�݆���d���*i'j$ĵeZO�Zj~	�{z6���a�	n�w���u��$��l����iJm���j�
��J�!ވ��i�I.�W�xw��`�{h��?4��v���YFz�M�W�F#�<�&�[�;,S�h�q���]�,s}��4����ߩ~M������'��7l~I{�3�
7ȭ�|�y'�7>a�n�fw���z�L8utB;c��C�$y��5����_����Ts�ZzcY�4{��L{�֘x�&Y�y&h�y���SO���GxV��MXp�B_޻^���C��r}.A&�#��|��Ŝ����rň#T����1��vP�By��$�O揠_�)��������M�_�?����1Y�Y��k����?r^����wOk�^���L�l񷩕r��9v_���`�&��a��`�e�x1#�Pt��ʽa�����8��.�x�����)�G�֣Tԡ-�� $듕Au|�� $^~��ȓ$����?������|/�Zb��(�-��"��9�&�	��'�c�_�h�	�f?�$)j@�pWV(B��F���
�Ю���x��n+GTRx6�5Ο2���3��~����}8T��2�u� "��}�}*A�A��,�}����g6#?��ha�{A�6�a��`5D��Zcy�?�M�f8}��4�ƴ�!a�EУ�2�,��s}�
Z#�`_��s`���w� �N��נs�vAZ~78_WE
�ˇ���_LF���A��cd_"��d���i���ﯳs��A�ɬˤ��=��#m�-vi�掎ͬ��a�ۭ��;����ļ_Cz���������V��7<���E��>����x_�ul�S���LR�K�ɶ!ݼ��㦲������̄��SÖ6>��9���T���[�gd��x�8�&�{��1<۹.y���RB6��c��$���y�p{�c�� B���S����a��UZ"�UdhەK{(yO��%�T/�^�b��v��{4����՞����+�t}^��
��K��oqlS7+7��"+b#*G.Xb�N����ݗ0�:(ט�P����{���6o���>lY�j�5iP��[�	���7��jܛu9kk�P#����z2"�l���������P���Q	yt:�����z-���	{T�-R���?�}��������'�YW���In,�`�z�����l~����������a6m/�����K�."�~�0.코d*�7�{�!ҷ8sL3���BD�&q42WR����
s��{�Y�~��ȲD),O���on��=vXeb���kI��|��e���D��ew�+���#�87"iz��l��\��K��SM��Dl��y�xySMT�uE�4�.�Ӭ�{Գi�ګ��Ɨ�Y��z^���j���y��� ���bs�0�"'-�S��3��ƨ�,��z���s������(�������Wҹ���5){O{����e��-�<���b�,��#���:�����.`y�����!�Ћ3U��z���(�Ь1ص�h%#`��d֍:�x�T�Q�T�����X�����[�I��B��.�f"͂g�FnL�D�m^D��wQ����+�d��-�hک�� �NK|�I~��p��:}W�$�nL �lY�.�i�lBL�<��a������Y��H�P����׾H��7I�塥��>홰��,z�W�hv�-����q-���8��g�9G��<�Jnu��s�t0�>S�"���f�R����3��8^���g��^���`e��p�#�L�Z�p�	��h��O�EW���^K9�R%�YUb�"�j���i�k})���x�2�>6Λ}y�� f]�y���	j��H��\��[�ְ��3�O��IδDc_��D��⾠�q����α ���\�����?"�a|B�Cl���Nv#�磣���k
��ѽq`����ƃ ���H��2ׇwpg(���_;������~K�nوt[}|+U	~r�b��SgfW[%��k�,�X0��gS�)����s�p�m�7�ĎBB"�z̭&��o,�x��pr��8���V��b�:R�N7>~5QjPv�p�j4d'�����F��&�뵦R��jBa4w�O����_R|�t��@P	M�0��>}]�E�up���м+k�3F�x@�>�:��w�*c��kQ��^�HX���rf�_D.D����c�t�%�c_I��!	:�Kd��R0̹+���\n�D�H�3�/�y9��%�軍�nw���l<�=��K����9R��G�s'o�M�zv��܅P��>�� ��a��_;9��[�5�����P����͞��Z
�M5`3��C ␻�͡�-5lK�ȋ�����ʼV���ȬT�/�q	m�0g~��g�z��&��=�E0�;G�^TM�y��!j�����+��u�f�n� �5M�F�N�.t-IC�̌�5ń)w��4o8�J�%$BiY�&��U�L6�N
�Xu2[�oB$�&GF������|[��a�/Q:��=� 
�`^G����0;���#]O9I
��Zԗ���P�?�U��7����w���0&''Q�v����\�0�v�H�a���wL\&�m(�K�5��ڹg��q��)��6���e%�B{���c2�[::���R�2�)8�f�>�a�_j���c��ٛ��l�[	1�?�,'�^�:�'�;��nR���ެo`���U�2���;z�]����=و[��R�P���m����(u��2���^�K�!D�6���Ez�����K�� A���QW���Nu�{�d��c�a�1}T���1��n�ʸ�E�D��l��w@�����0^T��/>�+�تƍ�aj7�r.!o��ۣ n���#�4��[�&b���gё�'��w�ܴ"�2�qk����	FH��wS \XRoo���ۍ��kq�'�>�e��G�o<�T ��,����vYa滋>�ׯy����h�&
@���$�����t=�a��JSB-��,�y�~@�_�ەD��|Az��x�e�nP#!�x���ԍ��O�ufA�Ɩ��p�*	�&畜6�N��i�Kj+���X�4���]�/>��o�M�xw���c痩&hX�����D�N7�l�G~f���2RFդ\�������:�ZY"
[KNҭ���§)o���"��M�/���@�Q0q��*��j�@x#�:F���B���X�t�H���_�W7-��HDF�10@� � �^%�=���'w%�D��\E�H=�`S��Y��~u1�;ܳ��t�	g��/E,n\�'
�^�6�Ab��`9V��&z���T]���v�Z.�g��G�|��q���Ty�:�i��*�-��f�G	����z��]|��8�
�w�M~چ��ۢ�S��ax~o�s ��#�)1
%��W��yu���vF�"k���b��F&��i������VmV����&��Q*�γ?g\�����y"���iˍ�l 鰰��<I #1� F�\�r7[:��+=5��%�E�)>������M�ZK�>��v��W�̼b�`jc�X�Q2�iߋQE��S�H�߾�a�3������z���՗f�_]g-Q�n �7f�ū�� ��M��DT� � <;��i&�
\��}ԭX7A3_��G��?ۀ+¹$�EHQk�%��L�kT��nB��9`A��c��'��7��Qؿhc����!�r�t
�8��Īy�� ��@8��<~�����/捒�j�#��6f��@�G�Y�%��4l0a�%�E@=+M����s#gI�B�[I�w�&�)�+�������[9�G!�-YU:_ŚwdP��C��T�
����y��'�z�>�Dě=���3S������C+���N0X+�Re��5yM8�d����+�4]]���z�f=0���x��̽���ϊ�~c�ӷt1o8��3�J�7�`iz]6K�C(��RjB�u��\@kߩp�<�"A�$��p�_VSBlX;E����a���o���� ��8�e;����ݕ��a��s'�B"�]�f�F��a��ܝZ�g�r���]�2"�.�RK�ɘ���&� r﷢�$\n\���p׷|KN����c#���%FY|���g|��@����#S]X���H�9븪��a�"��	�3�1��4��ɀ��z{��޷%Z���4���b:�PEϵ���aAy�X�w}K<$��A������R�;;sVXd�9�����>����8J]@�#9�-�^�Hr4|>���s�-�G�.>؊Dܳ����̱�z4��=P�Ǭ���q8s�Z��@�^���	j�F��~8d�4v��T���(ʯ��')�҂�~O�� 0���Yhw��/�Y�o�M��޴�Ąs�&X�ljF͎;�jvm�h�Gr�*:�o����E!�Q�ِn}:���%��O;wW��%�Q�
iי�c�&�s`Ȯ�n�����̫�&Ő��f�cii�A]e �v���nQj/_�6�2b���'�a�Sצ<�H��Q<C���;O:���p�mh���v���T���|M�����N쫞�}޸F�!��� D0�Y���7�ﭫgVU��ܥ�4��"j���,hj2sc�"���1����eQ�{�����Mi&���{��b��(kl� �zP	�d� �k�Y3�q�	�o,��N`�E
���1gy�2�?�!]��V� V�L�s�61�� z��80����0���:��7�D�cs{;��{{�,���� _~�Y+���?�����
�X{���w4��3��3��;}���Gh'��U1��@�-@ӗS�a��Z�^ޙ*7���u
����s������gt�uS[-}�����6��9	�^(Z�Qj�y��n�b�jfW>���p8Y��u�����L��ϵ���{��:���g	=��  ���=&�r��m����g�ǳ9#��$���}.�q�����8�d��ŸŬ�u����D�{��%����wHnH�������k��뵁��L{�����7�"�z���+��pu�C�dc�趄����£�$��A�!�I�~x�MӔ�ǉ�YK�Or���޹U��O�-k���:�ce�Q`���>`�
#��s�9g���,i���`x��簴�+��. �|�z�ǣ�O� ���� &���ݷZ3��	�>.$u �tgz���dg�m���sf���{�-��4��7�I�j�/�\��LUᛴ��ظ)���%�|:sMl�.�b==�����Tra"DڇL7���ۣ���bll|�gk8��r-`g��=��]e�:�����u�����iO�	���qjg}4Q{Y�̨tN�"}ǼT|Ǎ*�6��a�*
7�6�0j��E��d�q���c5�ќ��ȝt�����(�ܶ��	�!A�Iv��v�a9c/���(������n�(�&���b<2B\��^���=Ҍ��k������x� o����i @���$�� ��k ݤǮh�=8(����(�MN*��	��a�Y5��j�0uk��e��o(&�/rl�ȗ�x��/��Z�y'�g�.Rwdb!!�+�C!�γ�N�oH����1_�� p��/9~�Y��j��8N�����.�W�@c4ǻ+�N�m���`iCxǔ�n�{Ev�ۓ����� A����,�P-���x����Q�9�~�����\J=&a/����7ٺͦ�԰ %ſ�V@���Ҷr�l(_�M䨆R�=�~Ni���=��>�mYʚ8�s������2 dl5�N�4��/�r��)�P}c��C�����3�h�(����5��������4�x���pϿB����GJZ�j����%���/z�g�)z�Zs=SIy�	��[��s9e����2�Ł6P�+�ɦ�G:�|����{�s�_.:������?���=ʤ�P{�r\���h�Y��nre�������2,7��a�A#��K���xH�����Qg�݄�^a�#�Z|��֌5E�����A;F�H��wD�z+#�5B^�Χ�
���c��]��1��~����9�:e�CV�L[~�խF�aj�g��ck& ;Q��n�ӑի�Q�>�մ���2�O"�+��sX�<ｘjr��>��Jׄ�UX������\V���ˀ�]`���*����e�9H�0����?"��SHq,�ɧY��E>8_��z�'��]|����-]��K�H�h�'�0������<I�r���wԤ�glp�|w�pZ���ȧ��C��ݰ*Yi�n��<�i���E5S��L[?�Q����i;#�ϟ?];��d���𷷷�<��3����)��$��a��Ȧ��]-ф���U}Ҁ
[ۿ5�S9rp����z0�Y�Ko�!��ԬS{U�y����$�3"+Z�os�N`�A�$�ҷq�|w����L���Y��^踽AZk����\Tdd�ǆ6���W�X��w@q�/5s��Or�ij�&[UbU���N�SƖBW	m@7�|�Sl�)�����ᛊˤ�}���Y2�[�YrM�$kq�� }����l�x <F���>a�w�����; **���OR
��<F��z'�]��R�e��V��G�
Tb�r><���ZI���'22�*-9-R���k*㻴���hBm��I]��� Z��|z�<�@Xȹ�'�.
�/�jG�c���,Z��D�ƼW�-�H�.�wjYx�m8t5�Wx��b��f�@{mwAY^S� ��:�ah�^���i�ݢ��r>�Pi4 �)�c�khT"�\�q�����hGO�v��Kǅ`|����H��hn=�"��/	���"t�fڱ%�Q��|�9~̳ܵ�� ��8BxO/�b����[*d]��ŜkQ�񰴞�!4��ss�ewj4u��u���h��{Vwe�$�9�E�X���>�9���{�U�hC'�R�����q�����6������{â��}�.�P1a�ȳⰳV�x��Y�H�;���|L3�����y?�W h�'������nf�uML����Ff��p{����P����ř<��FV�C��ca'�&(����p�ɬ�s��7�ϑ�8�!�ok�LoKP򽿪q\Oz�C�:���t�@��?]Ƹn~|s�˻��i�Ա���.`I�z���	���]G\�|�8q�����B,r������Gu��B��15�dt�K�|@��Y޸�P�d�c���,�����VRڿM�a'�y��n go���>���(3}��A�-M��#� �k�!S��U��r)��R�\���ISi���%���Y��@(FY�rV\���1�$�ت��(��y��霢�����v5�#2��~��M�B�~�q���4�F�,��� �9�����'~�x'8�Q��:��sV���TJS��v�p�sUd;����޼R	؝N!�Z��G��*ρ57��u���Kž���C"�3m*�Wh-�H=������\J�Y署�"��3a�x�I�h8h�7Α%��p3����[��t � 9f1�ٔ!�g�vvܨ;3(©��f.�+M��~3غ���1񖸻{��j��|�%��NoG���M�b�c��%�?�9a�A;�PXaC��
��.�p�_�
B��M�Y�Q�1�-����AGIEK����r� l���&^����B`��05���.g8T��l����j�ȉa�?10��@~�q�x���C��5�Q���O�ݦ.IA�IȽ���|.����0ʷ����h��U��������	���gѮgי�Y���KB�W��[��&�]4Z��4����(�B��^��w�!XR��������p��n7y3��m`������IZ�OШM}XPc^Q�GHB2��]�i�^�3$fz�"�˟PK��a��[��e��ȕ�kԁqQ{'���`�Uy����h~\���G�!U�UV�$轴 P�{�T�>�ٟ#:a>��F��:,{�f.�|��l�a�L�g��z�F~0b���얆�8{h���q��L$F��22�������2G7~��,��:-E�vJ<:�s�C�>b���j��j����+������z��m��T!9��Ea`��7�yZ���DU~����o�Ht�������]�������"w-x���̺��ʶ[�� �ӌ5�\0���	��/!����_&"�q}(0�,5���_���	�q����H�����3���XX���ĺ�Ԏ�ʄ��S֔�;��A�3���>!��djEF��/���@�1�#�o�dZ�k��]g��p�[wh�ZJ�] l���^�P�E�9L�H�Ѻ�ސW�P���[3�^�s�������c�|���-���1���0��'蘮ʝ[׻b�>zm� h>�V^��a�J�^���:�s��[�įu�,�'e��f�a���9ˆ��q]�,i�M�@�8R!wn����l�ov�;��z��TX��A�
F$���3��T			� � ��c��1���j��T���ü�K������up���CJ~/)�V���(��/��)$����}PV��S��s�>a/���g�ȅp*��oj k!���/��w���j_�n+��=7ί��%m[L @�����k�v?�aK�=�����N�ؠ�����v+~�
�3kk��ʾxFiR\�љ����~�}:?#&xC4���%��
J49M���xƂ��U5��:�0��K�>�f�j���5P#Ǎ���!�<!�mt��C�̇z�U��K#7^^Y�Z3���\<<�&�gF��bmr|U��?k�=0 ��&ۋjXr���Guu�*���q�??Ҙ����wl���e#��*RL���C����0���h.6�0�����@4���[�h�02�g��"�X]g�Q ���l̘:q�&B έQ�_����/ӂߏ��j�	 +d��lw��
�߯��9�7���n��u��k�?:>Q��7�0'��:�u��$y*P����n����C����g��a�<!��4�a`�2ԮDW-�'���~���t�|��;@�Y �ִa[�����Yom:˘)+
F�S�90��e[���F��b�e�6d���@>�G�e�bW��;��4��`��a���̯� �0'�l9��/ĹJ<��fYf�w�!u��μ��
n��`�~��l[����ՌG�!-?`�Q�>?�;.:�$�+98��]���vQ�3��T�z߷.����N��OTSْ�'�mj�?��9[F����C/����!	g�����ub(l�70 !�����g�����cD���m1.)�cM�������JJ�.�Q,Z��li�#�Q2���ђ�>ƭE̮z�{����VG�f�����V��x�l����Ą.}�!��-����VsX�}4�W�w���5A��c���f��hGƇ��}5 {�<�yC�̀�9=�!�`:`��sKj51�8��l�~�h�=Z��xX� Cͮ�i� ���n�4x2��"��-nd�Y.F�S���e{���?j�\�B�c�E,Lt��X�0R�J�����.�!=�|�R�`���9��Ġ�1W�+e�"�\��ȏ+|ځU�����)%w6�i"��������{l�z����}Ԧ�$K'��qx������̣�cz��(&?�����g�֘���Y/����rI���g�f��Rj(".�z��%�s� 2*
P:/��@��=3����(@@�l%'|	\�n�@P�Ls�nK�z�yۭd�i����v��t�[|�橛x��n�v�wX� 	�TKu��4���v�..}��}n@VȒ��/z�&���Uv��Ӗ�EZ�`]L�t�]�P�>����Մ���w�H�4�$�!���Q��j��c�ȵ��R�9�B�2�����%*
*v�%*O�=M���b7��k�}�2�3d (���n�3��m���v�b`a����my{�d&-Dؑ�>3��91�!��Î^���?%1��ALgko߹���d��km-��Ty���N5�D��4>?KQ)-]�\�~��_el�~MϺ�1�� x�vBO0xem Y���!�:<.��X*�c~K8LW�4y�T����:+�;Z��Amو�MiRI��߆�k*yټ;��e�0�1R.|Y����[�p������Q�YU{�'��6�Oϔ���1r�����NGz-wF�l�;�:o��� ~�MQ����7����?ޔ�n���X�/ފ��NS��b f#;;{s{[QM�
���`���C:~Y�r��>�&힟&4B�Wq�Mu�-�˭��n|j
��R��!���h&%�k���~`+�e��n��]ޓ,�٘ʸ~J�!&�h��|{	򿻸�<ۀ�o�՜w�.#ro� ���rFF�M�{��7��y���vd~��|�����"����:�"⟹v��	Jt�����B\	��07_:���P���ca f��g~��'�G6��kj����<�����v����j��$v��s�I���@U뮯#�?:��CF�#S%�טO��������q�c�L�Mo,��V͏�V$���za��/9��
4�6�/z?w�Ċ�v���h�Y�2�O������,U55A99����";HB9�ϭ����2`�l�
�����Mc��%���y�w�okk��D��(9Z��Z*=##N(ţEv���?`JPv���'�f��-HʧO���sXo��]�z F ����T�уl2��Bw�3Z�����I=s�H�Є�����"��J������Q?�d���G�!�U�Ѫ��"���B��&9M__I
 �(= }��-�)�{����.ˉjL�&���{�(}��	H��&O���!VR\TQ��bi��g������R�^7߳�1|rX���uf���gxQ�8�-y�8���.�xF& #sX��z�Zp��t3R���n���ˆ�:*<0�h�@�{�V�\ ~���SB���&b�?�W��3�贐���Eǝ��M���n���9�1`�m���qt�n�3��'+]��y\�	<%��7?���z����*��@ش�Y��{��*"�15�o/���X����q=8�x�탨�ܖ��kd,?�1V;�Lw�P�X�V��%�}'DQ��v3��E���A�P '+k�f�@.�w�bo�m	����t�!��-�9�iq8tu�	L��8v������*�׃%Ա�v�^�w.>��k	>�PJj*
}Ξ!u������S��ӡ�m��^�13w+�(�
LJ4�>�	���������f�\>l�szv����//ޛUl"6
- �[�*v�U�i��z;���j}[z9��yʇ����d?�)dlL�z	G>����qſ�:��WZZ �8�iUE::I`Y��	Ø��R�A�旅��υj%���{^�@�7θ�w��:�8��#��oO�r6!�~?o��/���U7%,0��ծ@��ݓ����Ɗ����kh!����<-����`L-��
\d5}0<b"������NQcx+��� ��.��s�	��v�-�^�������R��}�z�ñ��Hb�gX�ueea�z��3ҁ�:�)��p�ߟ�k17x��#��l�M�3NW�d.�!�K��Ӈ�󀠛=�q�镯�����J���n}M�r�曱��:�h=�L��8K���`ߌM./�� �m{�\�,�c<��be�y�r�C��)&�Y�����ʼ��6����O��+6� �w���t6��Nϖ\V@�zѵ�R���p�
���= ]`�DH���6���Ug��t�-�*G�2����l	���|�[�m�7��y`�]�fl�=9��/�'����e�/aiD�eDǝ��M����<J�5�O���+����Q�d=���� �r�t�L��H�ï�ľgVY�|�c��D̥�l"��!��/ pn
��-HU��gԳ�~������8U"Q 2�׏��Fo���i����� ƭkcu��7��B� 2�+��g�QFei�����T�j�%�����4E���c�t�RV�������Ys��ÿ13�8���p��;�	�W���/�S\��R'�C&�����9�3�i�gg�Zb��2�#����2��)�T[[���N�f�/:�Ќ?�� ��b�����*��1�v�(��]����<
(��Su�B���ؿ�����]�����#[��Q+��?/��O�ڒ+tGe�!�y�0���gX��20y7�|hHNE�u��Vr�/2�&���n1I�K���F�g����"w�ܜN[�%r�K��vF���+9���+�����DC����w��=>�,����ʪ�k���q;�[�2^J�*A?|��S�����p��,>A3��o��IJ/C�;��D��ٟ#��@�.p$B�!���l�pש��t8���kM�]��a7y͠�����V''' we�:X�)��Q�n��2�Qds���.٤1f8<T�<�c���`�
]9��J6�##���o�.���lcNT|���&oGϞ0�z6	�]�*q#y[~�C�l�HD���}���DRNߧ���
��|������������
�nE��@�����U\��*��sL>V�q�^Q��B��s����4�غu+)E�x?œe
-�Y"J�}㦦�<���yï�܊bsL�Ē1�H䁜;��'nSؼ\�;���Dp�����{5����Q�����7*�N��Ɋ9�6�ea�m)K���Օt�pN�^�*m���P�0��'ŀ�j�NSJ1��}��1��y��
�a'��u���V8��{^G�^7�����P�ii����8�$�ɵ�9�[��h���s$5�A�"W>�g��?׸p�³خ�pq(���U��\D�I:=:�8N��?�z_&@ajk�]�B�q��|Kjii	H-^C���J`��\��ѿ��1���A���>��6��=&���n�����M{�j���\��A����.g�e3�I���/q���a��aq�7��Րϛ�/�#
���[h^�`9G��;���!	��s�gE�r�\/ (/S�j��5�,�����ߛA�}�$�z1�0))����
�4J�fB,���Y�?��&�d�E��<�ш���\���.y���`j���"�NU4G��
[4�tD<m�A%����QR��3�8���|��3Ab<s�:{������pZH�#�ٻ4�
%x��tȟ���3����o�(n����oPy�����e|H3�]TRwݣ���}WT�UW�����X��G���~����I��KX�)�#�I���{�}e��SF�����E�?��1M��^�1:�3텑���<}��9�/ƅ�yY��}�
<���o7�vE�!�A���5F҉���%N�K<bf��P���N�;0���*�wۘ�^S�.�妙4ʗ�.m��:<rt	��Jg�I���>��,�d������\%i_=��� ���4�y��3�����|���x/���h�-�I� !������S톁-@�GG �z���s��B^��u��z�;WgA�=io'�<	�k��ГAȑ�[�B30�3ꀩ2o��pIaFE�����壩�� !����0u|t'z��,���xM���"�|�)�����=*6�:&f�G��m�_�.g���H�n�m&��&�lV~�!������=%���s*"x��2��ߘ�+<����c���e������Y�rߏރlLDk�ࠋdu�#�F�.�x�vʽ|����A5���M[�4>=N6��@Q�� 韲a%Gg(�C�p�I}r3�q�^L�iǲHMH��m �{|O]��y&/nt����˜,]�'	��8��vj�����cofNf��%s�"��n����.=_usb�{�h����6G/�q�.����RzL��m�Qd糙u0,�(*=@�fZ=�k��v����^�s��>�'��#���d�Tj��<]��:����N3S��uŔ�/ßLv~[z�e�Y�T��^v����Է>�<�<���U������;���Q�{}�� q�!=i�jUp���������hh/�WG�|]_��`�J̚�C�o���ҒxQ��3��V`��C1P컑�	e(h��W��}t!K^rX7�U�&Q[*�->W�g�@D�&�{o.�������
�3j'�#��yqjm�g���SW	#:��Ej4���3X�=��w;kb����2�MJ�߭���}#�H}��iY4�bz�7:y�Iʰ��H���ёp���|lb�!4�q�[AnKwO�#A�V�
�<KJYF׋���Օ��@��ä���)����#d٬I��ԨA�jXtv1���L9�(�������O�c(w�6dF�+)�h�����u\7g�^.�)E��y�N�K�V���/<��Ǿ�W��(Qz�����;�(ʻ��8m2I�\(�<�:c~@8�w
r7���o+�_ׯ s�8�ҏg�O�u�4Üמ�z)�CR/����s�	��dk��a]�����+湳�܆�Y���$�h澩��4�ݬ8���nҜ��>=u!,��Bn#�3�s(�~t<4Y5�.^�uv"W(�cֻޅSآ�~���{����X� �eח`n����*\�É$PouP��c��?��n|����@����Q�.b��}���r���|��Q�����0����a��2���M3k��wE0V��G���	�b�lS���b��&���TI .Q9�������J0�Qw��&^�/C���Ĉg��",�� ���2W���`�U�>땻����,���%�����|}d��� ��?}�Je�)<R�R�Xt�0�x�)	��(e�^=��� �p?������-J|L��Q%F���?�'І��������'���E�����*h�s�]ٙ��� f=®�q�8j� =0w�[��ӨB��H�C}�	��љ��~���|%>�<��Q���������k�;���n�HiҤ)H���&�w%4A@�� 
R�&��� ��Ih�BI(A�=����˛�a�F��{�9�\�����ۿ��<K���ht.����"	QN�*��p��)�����՗R�ݽ�$}���/�u�f<�����c*4(��4�6@�`<##E�{08�Ϯ�$r�Y��Uc���;�l�'����%���_��^큳��v]��n���g�Y�>էy�O�lSW��u[i�S�zJ؍l����p�l���g�޻�8s&�[����ZP�U���>�񪕭�#;9[T��d�h��Q�#;���`���>zT�W������������o;d�
aI(��(�6����U#30׏اo)ޛ>��;8zfs��"�nf4[��Eӽ�!�^��M5!讷��.�e�h���6}d����� �+ܷ����%���炣�WXnP���gJZso���}������η�����=�rk�������7�,Jݤ�ކJ/���������b�nBk?�X���o��j���}�{E˭�� �`ŋ|��F�2�u<��ci�-A�t3��4^O�Pؘ�;N�u� fbW]�S�V��8�6��|����+_���wmxO�}�2���>#���Cj�0��F3ڗ�;lV���:{�����\��R��X���3�<�uc�nX�)}V�
P'��՟��C�ZGa�:���瀑ac�sw�p��k+Ò��	5 �`G��T���K�����w�]�6�~��1򼆌\A�f���:��׮���
{c*�3`w�t��EbG�]E>�׉nN>�~ȕT���	�_v�zz�j�>c�*��+��Uv�r���C=�8��mb����6��+�74S8f�M
˻0��o�����O�)����ɤ��9��9�� z�l�����J�a�������}����K��a���x�7����)i������Wb�+��"?�"WR�14�G/y��~�D���	�l�D��O�*�D�������f)��w>��
 ��N�~��nc,������$�\��$�R�
ѷm2 ��h����y�Ω����W2���z��-�/{SQ���V�+~v�bշ�d��\^2U��JR����(���\Q>���T��X3���1p���aER��d���x�8x�=��A��J�R*3�7˻�ք���<_PO�sMX����X8#u1��������P��OA����͡򟋧x�%�ºOw� �Lqɩ|�1/��wT�uG�ֻT<��>�z2K������-��z_�pڔ��I�)?�E�C���'W˰����%�y��m"0 ��hg�N2�6d0�X�uU����<���2`�6<����16�F$#1�l�#�;�lI�h��źS���K��K��Ffg��S�; ��u��`4��N8j�<�i��C^�-�O�X�M�n�OA�2�\��x�a��-��L��L��zqV�xH�x_ ��@��W�^��'j�����g�r�m�bً��eڞg��H�D>��ޝ]9�zB�(y�5_1�I� ��r#�~��O�#ۃ��������T��zߛN;�˳����4�����C��CNO��`Yœ�ĥJ�$B�3[��\{�g��\����zE����6F1`5��4,Ai`�_�+�':���p������e��1����ѷ2���X܂��'���J+j���Ey��{��U6p�B���t���y�~\�\<pށS·��" �w`LޙM_�
���X�CEa�òp�c�[�xk��UP�>��qv�N/;��O;�!�L;%0ڑQMC_���J쏨K���ʹsڻ_)�]�ԥ�N���+�J �*�0�(K����L��#5%���V��L�jn�bއ�[�#��s��Zʾ�ʹ#;h�߿"}~pɪ��PhO�wP��s�I��UOk��.����V�zaQ4�iַ�&�٠�2��Y��7h~K�m��G����W?�g̈\��y��-ғ���؜���/_EMkc9t�Hi.@�7����+(rܬ�`�(�Au��R=�,r��ҤxX[����͞=��7��S�}���4�Ō׾d����ټ�y��� �Q}Z��=#���U������O���oayQy���dۢ�[~�q�=<�{y�0[�S���7B��!ݦ1�IbQ���p�&Q�}�0�9)ЈBa��� g��v6;��0���.ϰU���o��'?�/�?Q�8M۵���b�� 84��P�AIz�tj��f2�y<x'$ȱ���$u������_�3]|����f�ѭN<��xl�|�s�Uty�}?+��Pp�(dS�ЋM����^Rq騏K`�5dag��h�����c[�לa�Ls`�P�-��Ԯ���3r�@8�B���9����a���/�%�<aS�{'����P-�?�)(�L�)���̦��@+����g�	x�����T@n8m�����k���ƢΉ����:��&~�GA�KCd}ξ�i�{%T���e(EN�,z��}���&O߭J�?��O�4b,�������������7��p\�mmgƥ�s;����\�^���0�.`��z�x����_>oA��n`n.�t���y+l�kv�萫?+߼o��q��?�G��ƭ�GA�A��g�r&��?tƋ{��T%����߈)�ٮ�_L٨٠��Wy/�y��}�pPab%L!�Q��/U�n	f�}�5�q䟻��x�+�<�q;l b���`n��v��E�b⻏��t|b"���j�Lup֋>�s�N�Y�nЯ��i�.pL/�r�B6����2��@�c���.��E���,���������w.���z�{�,�Cҁ�FG�mUb%�O;>��kb �O��犹�`��BS�k���k�Q>�޲��9�j� �߶~�Ŕa������ƃ:U9=cɤ@uѤ�/�/k�����BHݵ���#TFs����=��������/�Bq���ӎ����Kh��/#b�����F��ſ��]ئ���}����uf���%�˄�i���n���-�'�(�R���7��NO�e���b��rZ�	��[=~�_�I ���Z�QWx��ٳ�z=��|넘��R�t��4d%gw�"> �ʹ@�9�+"�z�C��7�@�ˉ�*ǀ��WTQ��Z���ѯ��5��zZ2�E7��[�}����-U;��'D�&hd�KL�˳[2q���1��|B��0�|���#�Ώ�2��JG�r[^;�怡���S�ҕ�#}R3�q�	��Z��ª����n���ɍ��d�PV��t����6:��z�d�m=�%���y3��X
��z�P/��51Y���b\||�p��P�$��
�j��7��^^c{�u��u�ן�U��d����yDC�#?B��X�8���!y�L��$�ρ���s�3x�d����?}=Uz�,P�\��#
'���fl�ή[���{��޴T�O5�sr�@y�;!�����s���@O~U��� �8���{���=/�H�RÈ����8���IYe_�aT��cFe��T��ߊ��A��~X�����#�*��).�c��JFl���2O�\m�ؼ1}☦�t�~$+����8m��?/J���1�%�p1�Q�E�Y��~�Hv�L��囓������p������ʃ�[*�5
�Ъ����pO�������Á�K���>����o�
i��覉UO�3ԸH�_[s"�D���wqw�tM/��鷃, o���@ؽ��XZ3�A�U(v�y-�n�pTOg�U�����o����w;���jE@�!��U���#!?o[R���m���W���^
+�*VQ�H*���T�zl�����R�Q'��nE�(�ϩv���>������<�	y��Q���r��pta1�?/K��j/d�]��S����YzF���ě�ra&҅�5����8G
�׮���خ��>k|�;,�u�u3Smm��)�:C��7�fX��Eg�.�4`r�<-9�~�L0�my�z&����K�M	�n��&�#��G�Zp[.`�ڌ��|��2����_�Ug�/:}/d20� �i�P�M��"�$O��(~��
�~|/,$���"l����6Jm���!�X�Y��^ ����]\]��������{�	[卍���*�~�~�2�u�J�ejZ� 6���JPȲ�s�r�]*�3+�J=�q�ڎ�0�K�Yuh'~�F^��}Fɪ8^)
^��o�a�^U��;|`��6�������V����:|;F�v�
�V���z��a�i��P�v���fc�*eea�'�@�ח���O�?�pO�~v/@���K�;~T9	{~^��NLL��Ɩj)���j�h�%=��U��𐰅�9��b�g{��Y�:D2��
9�~a��k	��p�X���g��+��oVɴ�=0��qP.E�ĥ�l�%v+��_Y����������j�=��;����6|������"
��\��o߮�>ZDJ�Vb)���p\)>`����d�r���CӢ������]�t������s��y1�'����Os�ӵ�m%F�!�}⯿2�6a�up���Q�:�Ϊ:M�f�iI�d;��lX%%�-ۄ�F�(��?��{�/J����b$A��Wb��@��E�fHx���eѫ��Z���U��B�ߓXo�e���V,)�d���q�G�����2�fdʚ�"R�HǶ*��x"�%N3*���>  A����}R2�0��~��Ù��s�r񻘬�N��2z5�t�ׄ�'i����N�Ҡ�SWS�>@��φ�_�5�	{"��E��b"�i|�Mu�`�C|����s�W��O�j�	�q��ƭ�ǀ��#�w�)�r�F���)���-���k�X����Ё\�O .&;�]a�^��3f�#x/�7.�<��0x��e���2Z�х��b��.�Q�K���XWOT�9]4�JI�����U�$u�#n`���w`j���y�vx5+��ߴ���(Q�"Rc��ܐ���Ί�=�\z�&�J���6K� �f���1�斣<��W���;�A	�>�p���*qCr��IP�6c�u�fլ����ũP=(��я�{�7�QQdȌ�Tcܕ}��~���85���Fأ����	�f=���$�H�-������n�Z��!�C�����{�|QO]����/�H�����ϾT�_d���-	�=���q@>r��m2�e�Ѹ>�JSx�mKES|'�HM>������)����g���`��-f���:tD�_lCq����1�эzP�@��gkgl#������
ߪ�/���b0�uj�����H�C᫸+Z���o: iJ9���HʓjF��DR���Oڻ��hC�\U�g��$��s�H+�\+��j�I�[���>�]8t�]��_2n��X���,:��-Y,�_�r���1�C���r��{G/+�u�p���O$7�����&%r���;��&�~��/E�\E�F���y��Y�t������lve�z��k��"^�zT�5_��N�xXW�ib��]�H1p���|�s`�O��1�-�Xxs���8܂�Ȍ��O�Zƍ��5�J:"\���ߤMW�.H1Wq*�cp$eV�U�+Eè�T�os��h����eq����O�fm����s��M�2��������d҅u�gjs�T���t���{�����m2�J[�	9*+�s#��F�,���b<L��CQvC�J�k E��le���۠�m��T�<��:ܨڶ�g�a�ߣ����< ���L���D�}z���������#6�S+[ނ�� ��Z��Na�9�����vp�\*[]L�A�6�BD�^���Qўch1��t}����\&���5a�od�9�G�'&T��Î<G�e�@_��&*B��n�
s�z�.��n~�Ӓ?�1F�q����-p74�n���:3�mz�#��[g�?h�b��\�$l�*q����¹�����ء&A��$�iE)u�����k�7Nῆ{�Eu*sf���F�iO!<Dd\�Y�$��P��n!d�u�WkI+rtl�㠄���������Ϳ�39���c��=�þ��\��	�l��]x=���-ʑ��
W�,;��Y|zRx�sy�;6tug,�p����k��~rT�>L�i�� G}��S2��3�C�Z�}��*B^o�糮3�>��/1�x�c��c�C=����$�� >rJ���|��B�y��ؓe���6��6��D�?{>�<��`I�ٙ8?%˟��ė�/rT�i�r�BG����*�q��2N��;[�a�߈V����̓�k+��1Qy��_�	�ȥ# �räʖ$+�2"{�7�bE�*�����k<��f~_�8
;E��v��5�^.H��t&P�i��\�Ou��ؓޔ����Y��lz˺��a��`c���.,��SK{c!R(��뒸.m�����D����s;���I�$2��e�Ӡ�úӘ��V�m�#.Ц�7`� �E�����>"�a�pP��#BPb!	�:}~��"�r4��*�ĉ To�ՙ�h�hrD`��MJ!'����5a�p9����sKTX���>;�ep�FϮ�1mt»#ۊ��5�5�25���m�Q�#W�b ����lo�?�ܶW@5�� �O�٩���|o_�&��^T�2���dU&��r��.|�%<h9��'͂��IV��f���z`�`9��&�l�ÝꙌ�f��&���i#�Ĥ�횓3�v�}&P��u@7����"��(��.����O`n�N�[�u���Į����0�1���!-.oN�D�Iw�s����gҊ7'}h�^�=�V&�F�[�u�~�_�|��@e-3�0�(x��]ce����P9w><����8�Y�����nt�����,b+�Q�8OgeB��������3��aZ+��=C�R�zۻ���b�>A$��c����#�O-�ñ�p�\S��u̅4o	�~mִџ���G%o��'hC��)�p���`X{H@9�k�D��������!�/��[9��(���Ї�z��`޽ۣN*!�磯���0�i^��#��p�(���W�_�U�}�l����u7�+�0����wu �7Y:��C�[' nA��pWݱ�2rpڗdr�o��!��6e#  �Z��z/��{��)�{�j��p�'���~�;�ၮ��;����b7�D����1��=ٞ(�P9�P#�\���J���5��_P�q��ν2%�1��+Po������0�x�	m��z�I*=
����3��7�y�I�|Q����X���ν6�D��)�uI-B�A�fu9s;GnIs�C':X'��@G�z#�E�ŻQ9f�j��&-#��LR�8�y
��2�j��I��#��4% T�nG'az�O}~�@�����GO���-�`��3Vv�磗��'��[��bʑ,e�Q[�A�3V�Nv���}���(�!�_	KоF�q@p��ȼ�S��m�%2LeK�������9������s�m�����M�|��(p�NG9~�[�dI�����4���3���#G@x��1����������4޵���C]�x����Ɠ��!Q!����$J$?VB�]��'D�j��;~'�xa2܇���бpQ:E�#��J;�����ȼuʙ	2��~Z���ݓ��̱��5��cIp�PNп��v29��o;���p�_l;(�LC�b���#� H�Z�ke�=Ѩ� �~ӿ3i��a�p�1�sӭg���=4�O���e�~:��ީE�������W�rX�G��|/�,gi��G^�[���H�3u;4���>�q���	�	�J��|���j�:��e
Yawm_&6�ǂ��u�����kD׹��G�\���`��eF#۲���J1��FG��/��v��.v�	��z��H�_�b��_���T~X��e�����*��&� ��m��[Q�4RG=�ܾ^?/P�l*p^���A�v�J�~�߅��^+|��[h?^'$�SJG(*3�k0�K��_�������󌽆b���XU�`�VL��%"����G�
`s���f�>.,(���sO���҄$ �`�b���S3�Yn!t{�|��dUs7_Ʒ]��Z�R)�r�np6f�&���*�&"31��f� �����#�\C���R�� t�@L[k�:Z�l���:����fΘ�	=O�Xr/�&�vE�����/nG(������
����e�����9�æ�٥���e_9��Kpŷ����w\�*t��_��"��e�[��N�1���h�//�.�O3�!���=�݇x.���儜L�H����[v���.�a�y�����G�'c �j�3G�t���r®7�3R]�P+�m�ܰ�����8�@��Zt���i��o=,O8��҆mZI��Uo����$�����:��|�\.;߀�(�@-��"����Կ�Л���Ϧ��Q:����ޏ�P�C����m�5�I�`ۑy���`հ���w5�Z~ƍBӇ�<j����]	G�Z�cD e���3�eb��=(���F��zj�"���w�&pI
�J-���[�q6oi"��U�`�i��ӱՇ��FB�K���Zܜs�Iћsc���U�`��'D H	�kΎ�$�i��#�$��B�4��=OT�
$��a,���i_���JVxh���'�������=�����IT��\57N��
D@��=�#�Q�UU�v׎�?V�.33�i}��gC�������n��q�?��a�qj���I��#�b�ښ�X�[UT�A�Xd���`����-�~��O��$�Zb|��9(\�p���s�16�����4�{X�g�я����D�%pe��,���w�;�K��H뢁?PBNB�Ph��y�+�޲Ӄ`�-�B��r���M�+c�Sr��N3���EK�!>�}}"�l q �+N�sJ_O釳��Q×��
^�DP���p+.���)k�HHO��!j?�IvUC�K8�t߿
�v�M����#:�}	�?�@q�3��9�[����֙@�!�U�r~>Ȓ%��'��G��FK��出�:�E��g�a�.�m�p(B���z3�U\ѹ*g�0ɛ crT��׈���G�$8O^���T���>9	��pa9�j�<��'�`s\�|���)�Nߓ/GO)e��L)����1A�h�h�S��fbv��5���0'|��ݔ�"U?s5�=L����}r�a�}A���S�v�H{F�Q��ř��O�"$�,[Sx���������]��JK�k����d9�p�h(��fn��A��Ĭ��0��⢜��-f��d]ϒъ�&��@�s� �����U��
�p"
8Ucg$��@�j<�	�&�Ɔwn���Fjp�5ֺ��s*҂�@/�_˃@̏�Ӷ���	���5��8�?w��|�z��.-�:�d7<��Mϙ������C�F��(��ef"��	)�$����e�Bh:�?��c�l�B[F&�
	�mW�2Q�|��[_>��-m�]�)Z�8W��z����yu_�84~:�d��T�� {������4Z�%@�D��x���>P_����J��D�V��c��3�@�W�n�S~T���6	�o�|`�x�/�0�GRo�ձH�q��?\�"n1䝜�_��g�9�;���@�I��� h.C�3�|�!b����&�������m�$B����>k-@��V��n)l�u�����^'*$Z���Z����a*-j�޶�([gM�3-	R ��bB�L�I�lB-<�m_0A~�.�P��!�(���~�gfˏ�7��n��j��?��Nd�'�*&��A'���DpC2���,�/s�a�v<a/�WmNhϗf�*C�0F;���O�`"?��9s��.%)Y�yX��x�5�r�����!A껻�����Lo�j���(	 ��v-�����dL�F�^�rjO}�;&����j{3�z������Qh�=i��*���f|@��$q�]�/�L:^��F�k��i��=���>���U�P�)>���9vi�>���Tbz���R/�`s�Oq0#cnۣ�!鿇�6��OWk�휂C9��*���Rw ��7��6g]Ź�9P*���C��$�_�T����ɒP��ż=��wͷfB��y�����!�/��yd�6�� G8� H�:��lM�~���=a.�4��@C��_�m���N/;��%�w����aa�ax��������q���0�)�"
_�g��G*�&9-8:�]%��-��A��?��n�=����0�8��S� &V��]�TZ8�la�=}���}���X|�$ՑK>��6v���_���3��]V�ҝ�n���F@�7o��;}΃�]��M�-T����?/����T����n�Yo%Z.X�O����Z2gcj���i�A�q;T �J��� ���Z�C�&<ƼkTG�K>��g�>%mO�ʏ���0Ki�2_�^�2t2� D�a&r���ڞ�R���Gf�s�4�H}c��"�6�=ˡ�Bc�j�L�� ��V���3���^���_?����!/O�`��M��,+A�PU���2����ȏK�Y��~�[�/��sU�o�U���K@6k9̟$G���9Z�ԓN�j���.���ٺdDwW�xS�@:�д̍0m�4��/������\�|P�k�C�,����uo�呿�P"-P2��"����$1��G�倦;���*�iH�pzjF �3W���3���7Y�#K������i�lOЀ@Fd������|��]����v/VC)6hY���I<57������mqㄞ({9��tPn���u�������V@��r���=uG2e�_�u ���=��E�*�K���!V���ݽ���]j��^|DC���\����O��+.��t�"���u�?�����mxK�v��!卂�Hh���C�����_K����7�=6^�ݿSU;��� |6�\k�;�Qfx�_Տ*��z��;���Jh�<'�
G��ٕ	.�Klβ\�c����iw���Rr9�ٓ��1��lA�B�6�b��+S�j�B�eS^��/|�X>τ�>�9��+��5��y���l��$J�էy�\Ϩ�9%�
�n�gA������>-�7(��Y�b���W6x�+|��O.J���
�j#^���"��o�L��f0����|��q�"��vK�F4\ѻm�م�ﭤ���:�g*���*�&LpM�M��t������Q+AҲ8�%��lm��Z!��V�b���>����*��&/���T�'���'y�>�ܩ����gg܍rp�W�M��f��hh*�8O)��]�:n'bg��WٲJ5&��±�)s�N��oy���X�p�
E={��6��kȖt������O�F�R��M�hm�_O.�
8��{˦���Y�OG�d�F�vnxa��˧���/����8��={DP�u�eC	�Z�������i��!%��ϪG�(n_T!�V߽H�i���*з�zs�[P6G*T����HH����1`c,F�k�a�F<���!r�]���ӆ=���[����!���@�����h�:p� ��=��3=4ؒ�ɯ���R^��=�}�]���?�|�{矘��|fa��#���cÌV��`�� ��|,PT>���y���r�/�fɲ���0�"v@LH����Q��/�厢ðS����l�K���B���r�� �D�}:�v�a�r�v�L*؅�J�����:m�������h�2p8��p�Ds$˕=�ƌ�!\w�z]d|Ѵ���Y�5��i!!	�e/L���:��g(,E�y뜬�ւM��8`݊��e��3��G��	5�3S��m��礐����-Q��H^h0}�L�_��cC�H�U!(�Pr$��K~���]6��Rn��-2u&\~�$ܾxثU?-�]/؃c�OK���^`4� <�K��(LP�V��;�� �~�ރy����Q�.�N�C0Иh~�����D(�u�Ҍ�U���:�$�}���D��~��Sh����J:ˢX��(���-4s]"K��A�⎃�����m�����b������>����Jr�P;V�$JQnA��wjo�@��tGBWiCM���e΍" 1����i9�Ƥ.����od4_�P���&������>�'De�Q/Կ�8��d�� <�Huc�n0hEFu^Yh�c����!��Vzbp~��1���ُC8O��Ƿd�MV�f����뻻w�k��kȏ��@ �;/ ��lY�_4�$K�I��V>>�k��1�\��ɟGv��q�y���fO�Iq��Kub�l+e��C�P�,��\Cj�˭N��K�����,z���m0�� P8���M�c��ٙ�C��⺡���,6���E�Z�	�z�3�N��3�oU��X��f��v 5��t0��O�a=����EJ�ƨ�[js}��E�ٌ��8b����p���)"��It��L���*ɭT��yw��ن�1_VQ�el�+#���.n�6��L�E�y���H�^���2��#de��CѡRI9HfB��Ԁ���į��E�{Q���P�b_j'�t�y�7z9���$o{�n�e�	��V�rO�I�ݓ5�SůS@j
?u�@���{4�5S�#�-�W	�ک���mIHhU���}C�s o��z�ߍtF���y2�:��/�D��f-�c+�A�m���{�g��H�~�m'/��_���L�����9���JH�R��y�}���5�~ ����(�>ʖ�وݷ1%���� �y���" �1 c��?xY\���&�mk�c�l��2��0��1��*Ztt`�*K�E��[�O64Ft�#{� ÿ,1�5��;T�ǟA���	�j[D��F୭�gZ�^m<(���6��OY�#��&~�z<3��B����+���lWIp��p��CR�ukX���HC�L@F������8���F�n��.ش�!K��kļ��*>!DUW8Z���of���̹;�����(�`�
O��>�Ͻ�WhP������F�<tJ,e�龰]=����$E
L� �����U��aJ��㉖mMS?�o�ً��-�vn��U:߾W�	�.��:QpHk�̘+��#�׸�`=ق�.�L�P���<p2{��Y�S����QlL[�B5螎��t��X�M�ٵ�tѣ��p�S=�i�����?��f��<�Suo��"$7psX����H(��L(�&_k�C�[݊��q�k�Z"��n���_El�\�����-R��~�Z_�ңs���5.�rYL���i���5���o%*����]CfRt`�m�^�\�ㅟ�<���n�R	}ڭxߝ���5����?e
�S����"�%��I���a�d��ѣ�Ͳ�����*��Y�'��/�HJZ$���S��(�F�s��?{K{��
<շ���x��x)�5��һN��E��ٿc�r�=������tY�����ڬd�K���UZ��٨3ӕ5"US���cC��b��U�j����7�*C��_W�4D�￧B��d��6��O�=+�ƶ�.�Yy��H�	)��q[;�>&c��66Iy�w�ꋬ+v`�kj��L��&r��VX�U"/���m�ʜ�9��I��
�U�:2��	+��*G��Lo�a�5��U� !�L�w�(����k/�� "*$a5��z���C��?=m�7����S���H0�����iS
�2\��F$>:��	iU��a�6��ѩg�5Q�p�d�����"����u!���
�N�-O���7L�kS��`hf��}���^�QآNF�j���)/����iw��П�y>�9[)0 � ���?������)�%e
����84����x�a��~���y�CH�8���a�����!�c�߿taD�=�Z��qB��sC�
F����d��E~��?�����|�[���A�{s<YJ�F��v����5�_���D>��-�'@�j��m�����	����?�a���q�!t�<�����I��Wm��,�`����͓����fR�Zz��f�Kt�ɣ���픪6�=��A�b���7�>�o{o ~�����$�t�$�y\D^IC���-3(�\g��m�i[�N�0���2��m .��y�����́�|ڣ8څ�y�ZTIY���`	者��`c,�&,[�#�{줡Η����k?�B4Qh$��"D6ꃩ����|�o�@��V��h�:�y���uO�#��q��RS�$lf�I���㞔�R�YT�����X�y����u�fpy���0��0�$��=�2�>��W
�z�F���*�֍t���&X�,q�Ϛy��	/re�(E������U��6ݭS���╅��W�>����YTgnh~�!]��GR����˹Ļ��vv��Ҝ�����Ø��p/��2��-P"�'^�ί�	f%�6
A�A�<�`Vb��ҀB������,�I���b�����^���U�(��C��8����o�e8��4��2un�ˊpKa��.�5��h���B
���O��\�QL�v�o��Kp��I�M7?HU}b
�_?a.f�u/|�w�b��xr��E��Ժ��EX`Њ����d���~V�(�_[pzKݠ�)��T�`�E��-nO�Y�咦ؖ\�'T�+�1�9����,9!��b����	�C��	R�j~%6��>=g�@KBW j'���P�k�Ï�\%d��ǹuOjP^d�qXM�ڹ~/�b�lY�&�c��sDs�%/������i- �Ì�6�c��G���M�I��Ւ>ߝ|:ٺL�d��Kn���t�"�<{��b�镐��;m�5�z�Ny��iN�iBrS���Qwr7�oT۸VͰ3��:��TO���X!���nݵ�t���F?�9t�蚤��I���4���	�:�Sba�����������)/	���lZ�����e�Ƙ�Y�2�0��R�JqD)�i�;m�=��f���2)A�W�v�����һg�T����M�ͧ�nd`�ϱ�	S\q��IG��I�x��j�Z���z�e��rf��)�-������0k�-������[;3C�������=���I^q����^�lҵ� �!����i2��(dў������4 (H�_a �v��5:BY��e�BX�Z�ZS4��D<)�cx�Vz�x�T��}3m�t狤��]wHj��[i��m����L����6����'�͸��"-Vc��c��(���, �Y�,��p޾4u�v�@	**��i5N=ywK<>�����q����E�hm�c)�e&�����̇)[ˆ(�iZY*��,��)QX�l���Y�O?0�p��	rݕ�{Dx�^�%��G%�?��{����=�����}�_����YXNy��j�A�z�媶�PK   ��!Y�;�К> � /   images/277be1dd-7489-4b2a-8eff-ec6391927629.png�{�;���w�t�QI��PI�T��pʾ�{ن�M��T�,!{ɾ�ef����1�a�ӌ���ܣ���{���\�_�뺺�ܟ{y�������D�s�=v��!M�C��Q���{����q��o�4M���G��ߏzkX�:������VWc�x�O������n��t��t���:�{;���qɤ)�:t鐦�}�'o����&�;צ�p熏F��_�6rgLT��I�.<����6���L$�<ʋ8�j�1^���ߗ�
��{����ޔG�'DD��fN�Hn`�3ȶ\g���Y��W�SO������/��X����������l�[�$��6>|����}9�������7���~����?"����#������2y�g�L)j��b)���_��8�n������]n����H-�opm�Z�`����}Qq��S����'{�2
�X�|��Q���wx�yx����̿k��ט�Иy%�*u:���QRR�g���A+pƛ��L��A�ĆqUk0��V�c����c@�9��i-b�xo�Q���Xj�RNB[?��ayyG-(H��G���{(��HE�A��iDU̐�~�CUT)�\D�ōJ�L����ߢ�c���?$q\lXZ��a̙-Mv�D���==y�����Î�J���(�[��73���Q�gS��q8�F�n�HxN�"sRT^^��U�LLɻu���z�>�M��)z\lf�R?�yY�%�>�z�:�}y�m����I^�������j��beu�V���{!nY�k�PI�����id��q�9!������ؕ�Fۭ[����[*y���w��z��v[����J.�sF�붞�Q�����Bjh���ۙ�z��e���
4k���u0[���	uXJ�a�C��cN���AOPvXRhw˫ciSSͺayY����ؖ�˹�i�V~���T����no�|������9�{y73�ԩ,B��F����vB�0��!^���;/��G����{�t���q�Nk��rr\���v�)��<��p�oUCl�`c�!��;�e�] m����eC�
@/%r��볉V��}��>E	*I~�j����g7_���F�g�%�=���{�C\Rλ|��}w�'�"
rN�v���E�)� a�:�c+�����9�R���F
���6������+�c�����i�};̿���Fh�.*���L��ѧ�����wj��dk}i��A�9�~�~}y�=\B_�]!�⌟揖ɺ������eeGq�7�W���v�RU�ii�jQh��q���U�
��`�ID� �˳/s~��V�~e��`K?�@��J̮&vw}QO�gU�O!�k�'�&�ؕ�����{Y�D7%���1�0��� �͘8��/�m��4��#,�<�p�Zh���m����(S>]j��ߗ{�ӵ���YH��?���FB��B�?�UT4�n��+�v�idd�������>K9G����M[�����y���������o�֥�F�U����n&��au�g]���~��� �m�cnB�`G��y&i�E*2���V�j��mHL[���ꮩ49B4��"a[��G��)U�X��v�<�i��<��f��3�A�Y{��q�Yv}bt�c��Z��}l�O�[���[7|��9���hJ>��D�"���>J������@�/��].y$@�4l�%Ի�M`�|�1�R�i���R�?�A\�V��ӕ^��~��7�w��]L��p0NJPg�y�X�LJf���&�e$ܑ�'�7�/��)��m��S��GŞQ���-8�]�O�h�ߚ����8X�e�jK#�^Qь������Y����5LK��x��ڹm���$�ቷږ])��7�s^M�R�ep���a�0<�퐷KoT�W�u����
pl��`!�g�@}&�S��C��Q���1�')A��=Ć��[VvD���s�M���얩%.v��ŭ���иcc��m�ـ��w��B����dG,���6�[�a/(R�
�HIj}G�[�?Ѹ�T;�`��`�r�rq������B�)l����*�����)���q
/Q"�>ջWQ���Cwe%Ey
�1�I�؜��0�b@^��|�$���>� ��a���7�>�-m��_bF�<��������g���X�R����*��C�h�S�oiSJA)�O5�$��q_ٺ�b4�h x�ʎ�r���A_��«�hV����w<�8R���@ܼ�_�Im�����hKk��ߠ,��d�>k��?��S
�S�,��ᒾ��y]�`&��@�t�K�@N��KL����䞄w�z���cbc��n ��S��?�ׁl.��z[�={������A����<�;�+ai�6%;t�j��N�����?x@����sG0hw��$�&f�<bbc���+:,��!�j�ǌ�����[R~*5�a5���WӅ�C`�FV::�N�6���d���船�Ɓ��\tNur������]|�2ڍ,Q��c��D,H.����W����N+O[>u9yez��������^��M?�\��1^�W�c�x�2n}�[�^m��)��}�-_	��M��+�x�7�*A3zz�X��S|�5~� ��ʿ�E�@q���;�����Ǎ�I��sr >؆�����VI�d�z����ܯK!�lV���5F׮���//?y`��Ɣqrq���\P)�ٟ��54B��_�Qkc3�{��z��_$d�}�W�S=".�1N�𙖝Q�A���P�� �����7�4�xaX��'������>9�Q?l<hW��'��|���g�f����^$$p��#�w7�)@�g��#2���H`ؿ	�#m|n�ꞿ�;�jF ����H�q�@]_��<1nC��SOb���P�
�J�� mV�xꊫ�v�ʃ�j�X]ի�~JL���$�HTdI������y�r��d$�3��b����/_��<�\�3�+f���-HW����Vh�7��
ţ4m��������V�#x����E�߸^�K,���1`Ja^�a�j��V�ab%��n��۹oѭ���7{1� ޻/��������5�xt=ca����,OX1 T/���+<����F�OLI)���'x�ʿɎ�Лۈ��I�tP�ٱ\�2��׊D�A� m��������E~#�k�zw�tV`2���Xejv�h-�k���\�a�QL��O���sFv�j��O�����5�֖����Ic�Y�f�yJ��f�h�n���+ڍ��B�хFl���m������fڛ���f$�{�p��� �C�C.����mЖ���	��_�l-�j�9�>dPDJ���Pϒ���nVf(�"N��A���;Q����W]�Wø�]����!ƅ,�o����.��.O9��i�d;L�,���)]�Q#�y��]��K �*uR$z�AAʈ�q��c#s x�qAA.'�G���-�,�o�����������<�B���ߕǶ��|��ez�P�V6���Y��Kn�
�t�s�uF}K����I�1"!��㌠X���ܠ1��W���н_s�����+e�ew�C���]Y�d����(��Y��O�io��Hp�*��������R�����A)(R�$��844��{C�������S�Py�5Zj��ޤy��H���yD�Wdg-H�2�]�y���j���>��0���*�W�A"�'0>��jϡ��r1����A+�#Ϻ�ǔ_����ָ��'t����I�
	k�N��C��md-ZP��8�Þ���K�C�MWة���v�6gQ�# ����`�� �C}^.���S�.��3�k	F��Q2x��E���K`Ѕ�g��XQ�m��e����㯵`_N��d=r��,9 8����gմl"�^���ߟ\̔qB���� J�UH�
�c醽��:��֧؟B�p!v@+~��I����'��7�P$Jb��(���>TJ�;1� >H��c��:����TB�V���͛���(�
�ߠB����a����(#�~����Eg�H��D� ��'� f���]���Y1��x�k�$ r$p0+�#�/B��r�T'��B���,XvJ�+H�f���U��E�W��
�&c�f��� ��v�z�D�aP�\�\���Io���M�^��F>2gg��F��A��S0�PP���Ǘ���򙦬P������")�]�ƇՍ���g�2`���	�A�-�XR䅊Ա����4%��{�K_9��Q��65�s>��S�+ː�X�dUhQ(f;|�c���[�{W�#uڿ�h-�:��,����80D忧�I�"0�a��I��&`ď�[+�/��@��������f����F�ݏ#26��X� ��N-�����O	}���1���%u�I��|�3�t���#�"��ĸ�-�=ok����~�
�X�3^47�a�J�*r�0��c�uKZ�Y��+�a�X�T�]\�5�� }F:���D;X@��+d��^%�)*2� v-3ϑ� ���HA��lBH�����>�@��u4������{\hʠ�Q5�4a�_��?��al���ķۨXk@��5���>�!J4��\
�icipҿ�l�i��`.��?DY�my�JX)W]|���Fc����"U�r�%�ս�r��A�֪���n/�wF����A�6�^* ��?�\����C&h�A9���0o*����p��<K��� �>7\$���(���zy6�����E+���.�;� I2�!�²�j��`?�V�,�5��5��TO_���$n3ǥ�l���������%A:�M���iD�@Ѓ �-��{���;tO�������Q�H��>�*�����HKI��#\z�x|�7�����{��w��CVK
f����h�i��ݏ&"��aJ�/̾��?��D�<�c�p�6�.ض�>'����*�	`��e�|�8?�G|qBb��}�H���eL���(Y�m6�FB��3�V ̽��z�y�c#��$6�pF;��"�g�]�ܱʉ��~F���%�������-,��*R�S
9�2W��|��o�Wxlx
�S9�۩���
Yw�L�Ĕiщ�#��pϹ
��ŸF;�����<0`��e�b�|Kn�.Ku8�x���}��֗n�A]P<�}�&d:b	Ҡ���UT{���L��X!==O�Ck��HE��̝�^@2�m��gan���$&�����6�����l��48���՛+��$ �O�I/	 ��	���<G�V��Y���z�I��細������&VVP�k���v�%}���5���,��C��L�?c�t�(Փ!?Y_���Z2��TI�֤�ʾP������gU��Yw�k���Yh[������F�S���N�kM�Zn����k6^��r�r���a�����{�B�ю����ej�,@ҳ�S �&�u�_�p��Y(<����?��;~qO��3aH�<��2�2����6�s�-É�唉�G�\u�`�+��9	F��e�/e@j�'i� ��b�����{_����8re���O%�&���Tk3��c�څ3f���_O��������\�dK/����;��q�"��8���D8�Q�	Y��u}�%�x����
/����̥�-��}9�������!q�s�)�B0:O<>)�����5��"�7^�5�u�Y�#�:)�.�T�!S/�Q�B;X g���m�lG���b���M�#2��Yo�дW,7���Q��!�
��*h�����E�V[I���^�!s�y]"�>�����T]k�턻���o�C��{:�J� �7xc�w�rFz%B�z���`N�A �OBc��\����[b��3�엤oW�'2��_�w1������n�V���jt*�yn�s�'�Ge����L��j�ϳ?m7=����s��e�Yav�Z�?5ۋ�<��̫&�V�nj���o��E#=F$�|�*`,<�ʩ��S�
@�C� %�:�b�;�  L�6R)M���Ky�qEN6T6-'tl�����!J�<��i��[_�e�ͨ:�?�������Qi�J��
�g�=�$��~*HJ�X%�&�>��%�k���vQ��o1��K�;�PD�Vx�m���/\<k��n�oZ����s�G_�����/�XU/(���ȟ��y/ɾ�t��q��]~�|�B���,�N�a�נ�f�����q }�e�&s�S�+>*ǘ�B�#��9Gؕv��[w���0���m����:���:�����7�O!���i����K�[5qRR����;Ь3�W:.C���ŀ)W~zw�m���%����Y���Y����ͺ�oP��E:�BL���;�>1�!��9 j#+�ʨ���}�e�u	n��	�9
8Y�4���'V9ì�m�gF�N�1���zK9f�Դ7��=��Z���W{G�@�6��l~�x�
��UzY78.��V�g/g���Wp(��X%��������{M�n��r�1��y��d�n�5�!�z6%��4�LOK���Z�w����S����V��|���94���Ū��'Y}���3+��y�kl�<�]=SQo1 Pf��z�ո�J~����®z0����j�	y-V��H�0`[��<��RS�Ǫg�w�WT��ų�!��mqmw�4��ǉ(p��B��99,�$�ɞ�B	<�fa�w�v'�zI~�~@@�SЍ}���<	�;�6��P�B�З�hM"�A
/͌M`�1��UA�s��?�B����D�VA��$9?	=�C�W[��1x�6�&&�����ܔl\�ל�e�5�f�V�H�:����]XG�P�ǳe�ˋ�kc`<#Y�����$�;��k�u��i�B��!�.�(�Lک�D��k�o�4��� �zʰ'�04l|!0�9�#��#��S��b��f�{�)AJ>��G��6[��a`=emKr���z	�T��@��4�Hb���	��Z��d�j�O���'8ٖ�� ���<�N��+���?�?�i [�X�B��+]��ј�]! _���|�F�N`�� <w.��@m�tG5tRAi�\�I�U%7��S:�8���J�q���.��
�%_�Y���ܴ�(�	������.��.��ҙ��D��ob�Ԋ.�=ٽ3��e Q ��H����'�$(�2���k���B�&dy��Y�x/�:7��/	��#���^z��Ma(���1 �O���B�s^+��!`V�/�kz��l@��)yoJ~��K�-'Y,ch���5q�r��;�V�R(L� ��]���s"�C���GA}_y�� ����-�C���2\ܱ����rk�ǽ�]1	��m�}F.�Q�Q�dJ�����E������&�l;;�Y^,/T�ـœhs�_�D@Qf��g~&��D����/K?�Q��_�9������X[S*�����>���pH�zmT��䝟IPbaL`�����e	�SH��#�B�}9�i�J�"ېyvP�k,11��JJ�Dć�D�9fH�"�&.���k����> )�7fxmH�dV�d�������F�4�����GJ�TJ*��0
��v�>e�B��ɕ��j ��:�q!1�=��봐��@��M��QI�-��*5t���K�߬��״�y`�[6<<�����t$謻���y4�2���7Q��~е�햏�Di��8������	<�-����aLV���݁�Y�����9r���B�#B6g��h����<��	��\�U!������l��Q#0��xw��rx��dk�m��܌,�R	���࢓��5!Hq�Ia0�^i?���"�>;͊��ů�'ݎ��KG߁�ecË��[�l��r2�rNK�W�����l���`��~tĈ>�b'V�ђJ� B����p�{,����Ŝ�K0L�o�AV�;E ��$0�6�G��� Kaw%}߿�[ǋy�$�_�B~\�a2����������7a�[}Y�:��I Ѳ>�mTYr@���R!�߸�:mx.�(�y@@���O���+�ќm�5�r@�����@A�<;u��F�{���$e�B�Hs.�$Z#]ɍ,X<c7��� =��b��E@_� ��.����ėD� ���
��;�IWi1��^P�.�[�.�fBt�m8C����X��y����^�G�6�mtན� }U�;m�}v��u_��u2eW?��6���kk��/�=0w6���<*K�C�w��h|yz��]�-$��=+�7�ɗ䍥��yΒ�E֦^��j�CjK�cN#y
�6�)qƕ�MjfT<�!��޹�2�U%u�6O�tHMt��o�v���tÿ�a��x�!��?���F#��Dݝ��ڿ�v�/�����vX1��Pa_�ʹ��cI2����sP�g:��mI�Kv�6����s\HD��=CZrs�l��=����HE7�w^�>�qFX�NQ�Vb�W����S��N�=�O1��,bX��q�5��,�؏����T����ۤ 4���Z�X��\\8q;s�ۇ,�E#A�F}�k��<�"Q����:�=B��
V�){e�"�;�x��Q�)����y�Q���S!kˠ4}��
 ��VX8����KT����v	 )寄��Ȣ�nN�*�g���'��
Rk����2�*)�N��SK^�cߠ.6G��XO��2O,I���a��3��l�������J$a��J�'�jSݺ�W�iף9٥�^�� ���e��=�s�Ajf�_�Ӂ}�& �~���v6]���d���n�yP��f���6��[��?ޏm��VN���}��Bt�`�P�EFiq��σ���/���h�]�q^Ƕ*ͳ�嗝�?N��n$@����T�$&�1�Z�3e���_���A0�#�x�8�^=�i�)��@<n�(����C���淹���ԕ�� �_Sb��x�� ]��2rZ���϶�	��QEW���Tq������dy� ]/+�9w�6�Ho��lձ�%�9t��6�ݿӀKO���Bt�P��P8}���j-�:��E����Sjdf��Ϫۆ)˸f\�'��:��Ֆ���i���l�ĸ�'Z�8~�b�b��)S�
�Ӷ�N�H�,|�.������I�nkoĒ�o<�����\�Z��w��~cv��U6����\{)�_j������ͯ�xn�@��Ft���F�.*@փ�Ocn�|���%�,��P�xa#.4��$��9|�"�]���jz��X9H�Ț�VR^y?dj
�c�׻�BA��
�6{�}-t�*5���s�	�[��M�~cvq5ږ���c��Xs��t�Dx�v�N�Ǟ�?x��c#q�NpH�6���zl��c:9�C͓�γD�$7f;�6��"�V�c��i�-ń9�6[�3jؖw0�d�W�Q��N%|��_���O����`K��ax�n��ؐ���e��h�*��g�
f�5�Z��!�����������Iḽ�V��6%[�����e��3_O��c�k;�+�P�@߈ �����]S[�R�+����w��=�)%���fd�T7�SK��/Abpx�
�kXk�Gf��5�/(�х>+��6��م�3�T���,tD�R��Mm���h:M�N�;Q2�m���:�e����%���Z�{���x� &[���y�B���R��EE:�l���+t{%ȥ<S���|��6�L*����w�6ZO��W&&���&N��a�����3���a-u3�e��*����bE���§����U�*׻�E�/(9�#h�8���z���W�묢���XŤ/$-���H0%5h��o�s�$�"���j�>�zGY�ʋh��/mYp�)�
��}2�+����`��l�AVc�����>�z�w�����0���=�b��t��LG��6�6��u�=�Xij�
�+z���c�ۆ�[whB��<�]�ʼ`T�Z�����4<|\�Sb�YT4�=* M�� 
��*�=8����|�4?�T�õ�/�A�J)��@�e�b�X!`5��`j�w�(���6z++�ٲ���()뻇��͔4M��+�A>Ѫ���������Z�g�<���>��o���|�?�B��r�����Q�:Ɓ�8�#d�f5;)Cg��ҮI�P�����{;�r���\�:P��l�ҵ��}��2D�3^����#�
�Vx����<���M��5%����lrYu��ǾF��rx�v҃t�Z;P�M��J���bڃϫw!K�P)�m#BGr$�,1=�M��WC�Ҥ6���n�FF��(%��)jp�i~����]�����c3���'��K4�fL���1l'���_��[��mK��?Z�T�KN��2�)S�Ġ~T��oU��uZ#�i8a��w�:E%!�I�ԴǛ�����(OG�6��f�y_ɏJd��P�j���j���L&a�s�z�(�9�k--a>����JP�xc�:�������n�h�Dĭ(w9�I@�,��*#�_3���ͦ�\����
�Y믭C��2�}�����F�ꌆFX�l��eeC�=j�j��>�I��}�n��̟�v3`{�z��Jʛ����=}���sQW�^1�S�����
���u�ѨAkHp��N�H�)Zڵ.-�M���xQb'^��C����Ү�l�J,%k���4�]�(���a6ii��B��^p�Tӽ�t����ף2�}:��l�U�n}�g�	�5�d����M6�*�|�Q�ǶNQR:��pˇ��A�V�t��5�R�B�r*���ГШ}�e��d��m��q�j�ۤ�����k~ٗѸ��?�1��R�	�	�v&+>=J4���q&�dG|}9xș=���o�K��c�@�u�����ѯ�HD�O���m�E�!���'�N��o.),��)ݻM{,Us�!HWG;���	̄O6h1#��������*fM���nN|l�x���w�XgM�
VqinC\�Qr�S�I)�!4X,�� e�gRr�x��n(R����=e7k^�ڝ�:#�f����E��zX��p$6���3�b۰r)�m����Vhх����h�N�����U����-�4m��j*>ͣ�{��A��j岰���?'�x���}��hx�Q�s��w�R[�q����K���d�p�?�E@;U�>�	�~��Bٔ�K�r�SD��?
��2'"��R]R�g��
���np��X���g�sıc:���2~�w��h�3)2�q��F���x��x����ۖ�w#�7��3K�*��L�����t�o�Z�����r���Vlo�:M$�x?hE�p��1;E�G
���U�־wO���㬗ͪ4˗�-O��*���3+\�0GW&U��xo��<�m����V��~S���x�Ksӑ��+��p�q��� Q1�rJ�m���ԑo@,�R�Y\f``�]�,X�?���#��
�m���-
h3�s|l���/���@	�6��;WjM�q�B"��r��9Z5ݭiY*x�i̅�{BSθM���OE�z���	{�=�A�	zs�m����b�~0��-��:!r&ɬ"�um���w�^b���X�x�9�&[�u�za>�~EƏ}]\���$�3��٘��;�#��t����r��N��~E��d�����1�K�0}%��iBG���MC�U����˱�~�,�q��|C<��2Qk.���� h��/ֻ�q�$ڼJ�3ʋH���t��S�red��쪸ujd��8׭��eg�I�l�����:�K6��Փ��k��>Ƥ�����m�T@c��y�֩�MMX�K��/�y�B�:����5]��&g�w�����mq��N�G6^����'%T���{9�3볨U��3�%hg��XF�q�/�Ƌ���m�����e$��%�y(4� 񯋪N&�%�)��줮g����۶���kn2UvV������u�۝�?��@��3��ڂ��P7N�{��d������kfw�u���N���S��~ �N�C�E�'�>����>����9��T���
.�2�i ���C�М9�b�@3}ȏ�"]�5vR�~���IW
~5�KX�0(�>k�#*4�����J�Y4�,�b�m�99y��1b�
�^����?�R�Q̇]	�F�/�ΘWR*�V�������������Ju�P�y]��aL���?�ڙȋp'��B�u򢴣����淨�����*<��ֆ5"?���ύ�a�6�
�D���uR�U�Ѯ���3�ip�*�$��㲙�u�} y��5;��̓��n�/<
�Z7�ix%���%�},Y�9��,���M|��� �:�昸5m���O������T�ml�y��S�&�l�c��J�=�<��K��}�xh�t[�E����2������Ql�37_�u��U�.JgEw�����E��.��Q�Xjc@�Hi����\���w���p;u�y���Ѷ*;�2Kye��(b�`���m��,��A&�b�V��A�h\$X���Ҫ(���]��]���5��:�LZ��#N��X�K�[[���6�v{��Y1Q�unl(F��ru���������)����� ��,m �/f�LN1�ʹ���4ͮ�)_8Ь�H�W̚�߆��v�t�6�\+��fդ)�k�Jo��!�Kb��9��9�I��M�j���)	�,O��E4m����|��R@�_�"ƶ���g<�O�v��/��y ��κ���D�q�ų[i�U���f;F-��*!�>{&0�ڨ��ʗ(<Ŝ~�EB>�؟c�$j兒�h�m/r�}$���w��N�j��{/���NE��I�j����佩j�������vA4`��w�[�(J��RI��X���wL�ƻ�R{��KQ��69;z�Z%�Y+��#�C2�r][~D�0���?�϶�o�s$(y���P)�i/�T�ݏ&��r�{��"�xG�S��c�b��������jT��#�;
'6�ͫŞ�o��n�(��T�t���KG�1O�R����!Yq�~z=�x6� �{�����5��G�8)A�x�)4�u(}���)��\W�
c:�2�@2�f���+�C��!^bG������w	���s�%BZrh!K��Q�!����{��s|�t��P�{�X6�FaN#�m^Dn�Ŧ��Ǧ�!�Щ& ��[���.E�xa�d�~��D��U�����u��&�r���v7���:��ڿъ'���%n��L��xdF�0�m5��Q���k>�˲��_���z���9����ڨ��]=K�Z^��+���O�h��}v�3y����d���_��!`�(eDf�a�y���k�p{�R嘱k�6���<"�D�{�����əs9��B]X��p����O�l���l��*�A���T�Z��of�q�vH�����g��,GtA��W<��?�N��911�����MXx�a�����^�P�i��]�k0��B�ޒK�*{oR�S-�ے��JQn�	}Urh]���*Q1�b���LU��2a)z��u�s0f�����k��1�K}EN-�������&tX�m�_�l��^65��G�OFA�	-� ��*� ��Xa��-�8U>��� ��2TV��WD��kQj>�D_鷞�%';��{�6f�@�������! ��ݢ�
7��~�;�9�%{5�yQX��ً�'ى�����&S׾>�4�CSw7��06c�Sx�����/H���Vf2�G�e�Th���L���[7\�?���k��C��pٛ��#PG �H�?^Y�A�FX�t[�M�:𳌋O1W ��?��%��k�'̛����D�8i�0"��#��xN0_$ߝ)Ҟ�y���n��|y��.H7,M�ïΩ��O��*��ϴ;���lh<�C��1l��i'��!�z7�tԕ�ɯ���y�nurT�Ӧ�x�����9��n��_rº������]T.������vuؽ�:�Ծ3���D��/ɒ��@z5�� ��&�S�`��
�K�n�m�'kB�ê�Yy�ƚ"W~����Roc�E�cܤ����Ld�����Y�H֏s���#�K�]��Q�|[����)� 雷��A<?��-�Z��}�v����u�7��a#��Q)�Z~e��g�~ V�s�4�A9�\~���6�5;R�Uq`3�6��2���[M�²w���F�`�nV�k~�$6܎W�j3�%�^�g�[�)F*s����M�O���d=���t0��.�^����d׋��W.4H�=�q��כ�tQ8Dma������/�VP�����z�ΈԠIUv��J�R���f�H�����oƺmu�{v�c�q�fh)wf�JpZj��$�(��%<x�R]��JL�|��<Δ$YVĺ���Ӹ���>���7����3���b�C<��`��A)���m~��Ł�Ɛ ��t�Ǥ]��vV��l[^dp�$���1�2�`�l���d���V0?_�������\�����G���L��`L�X��J\ߎ�,�ir���T��y	�Y� �\'���y�w�qU�WyG#�pr�Y�H=�Ev'��&x�}��\�o.�V��gT{�"/П b@6�s�]�ʸ�v9����v�q����[�>��s��+#5�w��	˓�rzm�)eL�'��R"^N�~�LPK��W�LGANɘ<�X~S+�B�6R��t���i�-��@��z��\�?V8�:P^�{�I#��ׂ�b��G{��w�@���mk��i�5���q�����/�6[�ko�h:c�"LZ�s�(����tr�J5��P.����O����-�n����1{zn���m&�%�X���6��vP�����v�	�[4z5K��L���j�qѰ\_qW���S��Z/Mˏ.��kh;x�쉢�5��M�|Y(�C7н������4�Nٰj%�R*�\�j�ꨡ����#Q��Ie�]wF*�
nf���\���(�[o�!��kڦ"�3�Kl�k�۶��Zq-q��N�q���x�2!ĵVeC�a���|Gd�#E�s�?�����g�h�C����rp{�B���z�*h3t8\�+�ߞȈQ���P�h}L�x��⏈������q^4���.�s@Dv�P+�
��<A�|UM���4=*�� ��|D.&�,9���t�����f���������k�ˉlI��bS1�g��E�/�����#A��d�4�(�ea�BVք P.���u�;��ȴE6@\���^9e~�A��T
ؓ��y��2]^��Yg_��w���	~4�T�x�2B;o�D����E���;���S���_~(k��@���JJ=~d��""%m���۲ćxw�*���A	��GH�+��kǁ��qV�&qJ&y�h�ZhV[�i�!���
�c���F���\q��ɦ�	D�1�z�!��K�?e����Vmbr���s�d�
�FG�>�9���{�.�y.
��Y�R�"A�R'��͓_�Ž,vb7�}�RE)��
/�X۱����D}�h*�_�ȓ��kK�F��m���[P�Ӊzw/���豯1ޭ�ݹs��ձ�X][X�9I��߿�k��$���7ND��k^��i���b��ɹu��/3��Ԣ�\3�j�Q٪��a4z�����[~o�#8��߹�&�9��ShV��y�eu�$�h�)�L����$�Z_N����xu_u�.&�}��s���,}�%1	����cj��$�
�g�3�.�D�w�m{�f�:˗i�,$����e
'���L s�WB�V�2�AXȭ#�����}KЀF��:�.�E�N*������sKn絮�eɌo����\D�M�L�u���.Rq��C<{����7%���&y9���^�7��l.�_O& (2���=fo���ߪ����ʏ���ְ�C�^Z==ɩ�b+_�o����wX���{��%�V"�p=�Ӎ:�j��ݶ�*�b��]{SW�.{@~��њ<@��\��.+�g���<^�$H�~p�Uaධ��N�cq�ԻՂŔ ̕�-����l������bS�Z����.f�.�t���7���$c�C43�uw����t t�x��4C����D/%�b?-`Q���Wj��9��r�{^m�����m����6{��|�Nm�^9K�Rt�ˏF[ t�\�FsB�RĚ�#&/"��������N��F�j&xz��~c�O������U����Q�tr�]1�i�?OĮ芏��&����-��N�v;���l�\��z�#,"���">�{�u�o,$°��0���ő��S�﹍�11y�vH��N@ WUi"9Ú�/��pWR�>Z��;���~ʎ$�s��-�Y��J!�q6dE�;���8<��}P2)['�6���Lά��N��v�����s8.U?�׻zo|�23�W�W���{�1	E��\�G��cl�>�]��z���`8���no��%)���C�Ӑ�~�zo�Ѵ*o~��p}���+U����_�k"Hu5�?3r�66-N��H�J���=��Q�=�!�_�~v���"*�|Č(xIHY�ї�Т��\8q��y�ܹ9��OƉ����5Q�~�'G�@.j�-�*$��Q�?�q���z�/,��L�&2���̌��ʣIn�c+���wt��3N�W�e�|8�ͬ-�Ӂ�ߨD�>kS9�ߠ���hg�Y���Y8�;ʝ�(�BK���G�i.��?��{��d��^�f44��U!��i%������"�Y>��4�Gj��ʒ�|eQ�1[�����J�o}Y�J�q	޽m�&�|�f��y�R7��L{̽ךV2M6n�I>���a��Su�m�eJ1����?{�u31J���_���|�͹��Z��z=���aI'�@��p��աsMa	D�e���,���X�׷C��jު�~kܾ�G>mV��7�����3�L�z�!ogd�x�@��qyL]q���58��v��׀g�j��6����<<
4�v.-Q�!*2.����z7xJ7����M �॒����� ~���{��#Ϩ�+7,��9>~}��C��`��� %V�`z�;��������	�F�M�@p�<��������-Xp�w	���5�{����s�}�o06�ꪚUs�^�W,s���д=�L���wה��h�f�c�����{+��i�"�5�,�3���\��I��y�Nv�iD�09f}������sH�	{�F	즶�ܱU��c��2�t���S|΅�ҏ�|��w�(�fb`��{��0�~��P�v\?GK��cZS�>g��;>y��K��O������A�+J��>*vGA�J�������V��k���[0��
���ҢΌ,�����!���������:L ,�X+-���3�\9j���m�(����wu�Qb��:�Q�K�5�V��~/B`�tC��5���y^�CV�ls����Vr���Z}e��l�{�7���5�[\�cAp41�K���ۊ��kҟ� ��BS������g/��3�#���U~vd�?�����̋� ���M�/�?��7y���k�͆�g�����)}�	��!� ��װ8B��������X��,Ѱu)7߾byȺ\�@�m��,�f�J��sjk�6�L��_㈈�7?��@��T���f�;�$ +O:HE��+v��H]��Tu��W�iN&�-p�P�7%�'K�4�n�Ǯ������?�pɳD�~� �;�5�N$��Z�t8ﳮU.-N���0~�Gi���;����\��05S�=E������sj0MΫ�ß?�|�
j+�V\�ˎ�b��ₚ�HX��a���܌��&4�`�=N��L��m�i���i<N���ڪqm�*K���A�~�o��]�l�4B9�{(C��������B�,`�ҲE}?������Ĉ���#8ϱɻ�|��y��1�s\x�:^:bJIz�ʷ����~��աm�޼J�n�Ge���f��ǵ�^��"/(��n2�m�\�ƕSP�Tx��c�Ֆ+�9��NA��lB��'2w��{��C���F'�j��c����b���\�5�֒��X�K����[M��M}"5L<Lw�eR�)�޼F���^�L�B7��Ol8��W:�Mzŕ�B���V6�k�&%<3*c��\�%`�d9g�y�>訷��RYa!��n[k��&�j׉���ݢm�.�6f 
^�����B�=��4�&�R����D���fF��$��]�Z�x������uWE���ۆ�K���c���t��[���`sY;�ڽ�����Ѫ��_���M;���>��?�>��WMF���>ސ5M9zk�.��?�yz��^KT`�+��0]�/�q'y�}.*����:��,��i^;����
�s�������9�ez��ǔ�n4n$$R�A	x�w7��<?���kTap��2�}d�"!��&�0�VEN��������i�d��>f��L�ghYY�9rO7���{�*	U 	]�\D"8t��.��ci���&�YG��Ύe�$P������w�,�|�b�T5������]E���֕����@�*
*F9��:�5�?W��]��0��dr5���G"q�A�]����9���*-��P�ni�^���}F���\#��&�q[�Lr�2S��}p)�y�E���|�Vo��a�RV|*��*0��M��¤���5x�y]�󭉭��·C� �f���(�g����Hzv��S�8���bC>B�v+ʹ���[�I��E��R<���@��ݭ�]լ��w�a�����xߠ,�<�a��8�3��3U2g	��V���������x堵���:h'kFB¼+ʨ�����
�[��N,���ޥWGT��\8��*���auz���O�:��D�0�K^BХ(�[;>!̍IC�;���tx��խ=)(<b�Ń5v��3�@��}�u���n��K��U�4c[�5rNӦ�L�3��Ⲃ:l����a4u�ۨc�FX}�U<��C�u':�xu�{��$���k~%�4 �;��@}�ʆ/��	T��v�:fl>(-}�D���|��y�BXl��K� ]���~�R�M�<>�.;��Z�U��[	 �br�NEF�>C!�P�������)}���r��C�3��T��1)^��T�n��-�t��Ʃ�X�E��Ï��J\`��fp���7c����$���d�H�|��0��
tm�+���T�$�vqD2�Z*���fD8&D����Vݩo+̲'��1�$�X���	����g�M�ǻھ3s4��Ù�&]8�a -�Y���\��#�"�.�j�h��'ٶ�M��oi����ή���^AOm��-��'�����'���������g5`�O�tE�ޫ�XPн�K��!����ϼ?���M�»�K�N�%k>��]����[_|D��?��HD8ؠ�+�Ҹ�D A��&��)�S<�?<ZX�H�E�"�T�m{^��S�[���K�qmݶ�D������&�o�fj���7�N��s�:S�9�	�}�d�4=�r�:ij���5;� |�%�����Ƞz����j��d�Wq��$� �a��]_���\zg���`O����%�	�c8����N?F���$kT,m�B�s{⮜����n�]#(,�bΨ{C�{i��Hp��c��F-J�BUm���Ad���p�,+�gz��۲��f�ju��XlP�Y,��[D��1��f>�8��
�_J�nS�cc��3�V��hq����;��}$�TS��8��������@�l<���ېL� ";�o�,�� <J66�3 9� �ǻ�p}��O[�E���R����#�8H݅���c���!yM�ڣ��ބ/N��ҁ�ٚ��b{P���2RRFYA�¯G�8JRg�]3�;b�b��HS?e���5�h�m��IO޸c��ۮs&��uaW����l�S7'�XS�����;]7�m5�[��g~�ccGs��;�Q\�ug�e��Y��	6Z����n��4Z��
A��I�6σ��hѿ���ߟZ���=����>��让,��}��WФ#`bJ{+����,����HL-l�;�1aݫ,$ԑ��5|�*�e�צ�U�lMX��� �R\ɩ�]\e5HC��_�*j�+���Q�}k�+}�7#8��d>jJ�q�?Uӧ`�:ɷ<	�s��1t�`[���|�qyp���'�@���M�|Z�ek����!al���2���;F��x�AW$��l�E�t�թ�����K�'BN�z��O	 �+Ub�Ԥ��a������#)A(!K�أkĖ֘�N�7(>�D���g۳��BS[+`�n�H�4�dd �U&2��6���@�ԗ��x�åL���ȬC�OD_9��8[(J�j�1�а��Ŭ��_W�-��B	���i?&m�>/��4k?�1CL�Qj��A�ۧa���Q�#{=]����jy�G彘#O ֓�6Q�|ڃ ��Zj�|T�(HU�)z�)�x!jg�#*���[cc���c]�:B����.h�3� n�܈�H�`yZ�������غ��N����^�mC�Hi�����n�;�\WՖ�� ���T�Oш'�-�k����gg�U�K�ZՑ����܉go�S��k��2�����@��hX�
���4s�"A�H����R �'Ezu]�P��]V�4а�t��5L'vUJr�� ���?�)�G���UQ��X���B܊G6�S"�A���v`�B�=2��&����6����Y�b���>�zm�>�VK<��8t�$ xL���DqyIG�[>��*"���[��\=3�s]�#����!
���ښ^Cf���J��0�mU��q*����ك���>a��s�ш�I+�V§ ���(���L�GgG�5 irT}։�j|A���JW}@?Y�'㎬��X�\�-����_��>,3�n{�p�>M��SC{����R�	����GW���G.H�;?)��H`W�AC���'��{c::z��R�l�>��Բ�����6*O����l��A�O���Y<E�9�Rr�2����s��ɓU�OJlt��=���lvo�Fyyo� ~e:͋76�Elq���Y��t�,B@'�L�GX�A����ww���Us�T���t/��[�Oi���Уl�M����%,W�@����^���d1��kz�#��ǯ�k#!��rN�@/�>Ѻ�Ң�����sk|��7�rS��=�0�y������/7P����#�!"q�Җ��C����[[���|�'a�̮̭���@��k��w��<���|OP���@��U�������jچ�n--�t	�V�U��+;ې՟�0z���A�Ѹt�ܼ��R���ު,NmG;�Ӂ�1�����j/�OcT*gR6�0�HY�a�����}�u�x��2���-'.Z�f
/����Y�8smu�g,Q����?��'+F=���@��!A+ȳ
):M������[�����I����	�*���U�5K��6�Jut�!��F��p��M�k:���"�45ß����5��;���脃� wE/e�0�>�Fʅ�O��m�_W��&��U���B(-�l*"'�`I��f�G��Sa��!ԶT~�gHϡ�di��84��sNlG���0	,�<N��5O?��>��++��kQ�T��]9��}��.B8?�wKTL�lt��\u�-�}��M�����u��Y��JAv�4������B[�큽(�\�[�Q�EE��R��[��}l7BO+yV�OC��"6�ϯ��U/��"�~�����%�3FB/'�o�%c3O��wR�*Sd��)��><5�T˵-��&g����������F�y����=�7�(Df�d�t�L���{���
U�͉RRVw������C�ĥ߈.ɽ\k4X���/�X���Q(����"d`��ݩ,��PRR7۞�KIMS�F�rJ�$G�ڶq�~��9e�LU
SV�M��o�FoW�ł������_��������?m��G�=��e�R��Z�w_&����>��ʤ���J���^.�����os�-��&V����2�m����4A�i�i �$�.7�gש  |��\A�5wȊ�!m��q������p��M��V9� r�bKx�I��~t�sp�ф9H{���lֹ1{�S)�d�� �.�z,=OT�	�HN��(�����g������~����{O�?�rs���uxr�;M�Y�����5a�rc5�%Zh;�h��v	����6���[��a`�Բ�w��1�D�������&����l��{4�6ψ�cbv����GX����p�OU�a֓1�շ�%уV۾��aŐ"XFQ��ۍ���-]��X��4is0XJ$���&I��K�j&]�����~���h��Gа����n���\l��R�OpWR���iCܡ��OeM��Bd��Z�Ñ�bj&F����P�0jqҮ��r��#6��,x���Κ8� �I ��1fE��������Xc��	���"�5���5L�خ�K�k�%޴�cL\��8 �|�����>�@�;� �Ya4��J����J|VϏo���=��$��(,�Y&�M��ς�@�/���>�θ�l�$�؈H�o�V))�����.7�M��h�"���6-H|�}������D~�����V�SN����G %:`��k��x�Q�zy��B22do�1�E(r�Tq�^B+�Tj�~Pv�m�� ��Ғ�f*�K`L�p�z�}�?�s����D��v)�'uI�����X�l ��G��I׶���N�d�́��#'hC����͔�u��P�T)X�>�g�x4Gfs'<�r��g�b0P���"pDO���}�?#D]{�hr�Q�{%������X��h�߈�H{5M�Ȣ��"���F���gK؋���t�C�(�n�ն]��+�kGV�ި�t�Wx׳���tU�nS��ocՒ��3�o�p[����9G�[�E&f�������́��G����y�{r��f� ��/��@�O�;X8tq���*��-��Fs_����~������6}B[��&e%.ra�����Ť; ����}l��٨Z!�:|��i�Ql�ޱ;>0�;���?��p�����^��g��gn\�n�DS�ͤ�H��]\8E���u"�df�j}hLs�4�����hkw7}y��Z�$#f����ގ5����x�aBl�)��\R����+ U�[/1 ��U2?�S@H�=��|�~���������y�����M��S����Ԋ���$�s������*��lqA��LH���Ԯ<aq���;�Rg~�,��e�-:v�cY�@�]U�G��+qEJ�x�_}�a�\���F}ߵTTb�暗�y&yŮI�K���!�:,�=�wSԽ���P�TON�>�����)��A��K�ۈ�����|�z�>ؚCe���9����'��H��"_d�3@49}}��j��g�Y+�`D"����|)%܆���P[nH�����s"DD0TJ$�C�����������x�'����oCC ���^�l�����|��>$�,����]1�{�X`�����q'x�ʖ�%<ڝ�b��/\�����]N�r�ַ�@��2�I��&l�z��ֵ��v��vh��Vtagb���{X��uƷ���X�-s���ygR��5���:˄N[	
�;�e� E����1a��1�GP$MI!����"5�H��Ӏo>�w��ۋpwV+h"9�	,Q��-������:�")��1�W؟��qc��@��H� �Ny�+��\�K�m�Ѕ�2 �"RJe�(*ﲰ��_�X���
�K軳��	]K6A��Y�7�Z��R�0 �]GN5<xKg]�o$�nL�F�J���m����oP���e.1T����~��j�,-�
���}u��!��4	�f�&����Ǿh�"��xl��6�N\7I1��(�]����^����`b~>Y���-4��0����b~��1�\o��3ޔM��&���ɤ����M���JZ���l�a�����}A���I87��9)��C�.�{��s�5����jA~�
���)�|�Qkx�:Pk�DH�b�i���=T2S��#���H����]����9�	������_��o4 �N�rԡ}0&�uy3+z��^b ���e�),hYG��7���$�zI��*��8�ґ�A�Z=�րp��>#x$�U���tb�����z�w�ޏ�λo%��/;S���ZX��C160�$LH *萳��r��C�%*&ez�
7>�FÔ�)9hav�W��������g?��?�˸��.�������eB��e��J�ZW�n;�����M�[kW��!P��l9-ו�ph�K�f�T��h����%�t!�k�|!@���у�.���232��|鎭������Y�BV��-��f)��O�A�=ǅ��ߒ�:���Y�U��;y��~ lԀ-y��H�4�Ofj�a 9����kjޮ�c���JL(c�����ydbd��P�5%�gϛ⪙���5���S�jǐ�?��P}2���¨-������"��s�`���-`{Y#{�t�E��6$L� �8}�Z/�؝ �FiII}31��̾�!i$��k���ǈw_���Έ��oQ�B�8Ɍ�!|�~����G}$>fʝV��dMf֩\�#��B��̏p� 5q�a|���J{G�5[�;�B{p��"��Sf(���{���}�4!����9Y���LE@@��^'AY��	�C��3�z�f8�K��V|��yQO�(�z�u-��� ��+ZZv_e.(B?���V�����Cg�t������#�x_���f��:U�f���F�4ڣ��J4���q�n^3�n�����*]���1�����@q����Zmm�[c�{^�V�1��j}�{c�r߰.�}4�8���k
�EYN�I M+g���a���i�da��oB�(��T������`4o���r�����8�ڤ.|8Q]{�-����+F��j����^�Gl�X�f>����h�� 8t<f&c!�V��ӓ���dE���F!��!;�J�XY�t3A���X���)&po�h��8�9�Ox���+,�@�ܩ��㸷���$'����kN7��kh�P�)�_��@��K�A�9ܴǟ�pUl	�I���`�,N�a�܍"�IY[=���qi@�G�:�N/�?iԴ��P]Lm�W��U�%�{ݟ��?T��ѩ%`���5�>�b�8�[o"���`H^����-��^�z����b݋���~�i΋���Y �ΗhU{x��!BF�F?��b¸_	��.N�
Z���v����MW��9Xm��O����u�H� ����s):�����(���^����y�:�ti8]���:8'Y�\[�
�¥BxE��n*�2��/Q�5�XZ�]$�AlG8��u��t������L��25M�A[P�}���ۍ��?4�#C0� m���v�1���,8��/�������_B�j\��,D��2�i�PH\��p_u��Lö����"�QE22���s���.=�'#��ɮM�q����Gv�+;�'Zf6��ֳ��ut�}��B��|e8�:���űNWD-�'�䳺H����:�S�b��1b�B��H["�6;z޺ ���uh/@9Y�a�l�#�g��^U/�F��7��[�rlУ|�����Ƌ��m�
�|�RC��k��:��Ms����|�&�����N�x�8�1K������?{r;�i�^��=�y�Q��S-9�W$T�|c�:׆�!0�W��9�V��!���xmKG�Ah@�-�LElA��?W��8��b�� 8-��v���8䇿��|�Rh���&����QS�EAw��t��"ц}���#��)rmJ��m&�h\������W/�0=�����N��ML�O�P�H$k�H��Z��&ī��8�l���*}�����&�+Q;�
� C��?�7��ןLe��7'������s]���~2|�QT�h`��h8�OKK�bK�n�� I�@���������K�!V�f�u^������~I�.�{�q�NA-��j_]E�7�`ωї.�&O#$!
'jId��'�t�-����;<�w����s"��>��&#��������q	3�`�dl�ɶ0M`L��>)7wD�W�����z�O�涎�3�n���-6�N(�y˺:���<?�3�|y��t�Tמ�,ڃA�Q��>��+cu3~3&�zP#�	}��|��m��EC��,��l\}Q�R�ס+yû��LOY=h���eq�>=���������I#nz|��l�cib�N�����������**�\g��"�$��������F��@j�_t���,Hn�'��޶r�gmϾt�<�\�}��pS9�&�gVx��B'&��oWm�V8����NAǴ���[�㚅>�9����5^܇�mo/N�>�M�_D|����ս �('fF)��RgY�>��Q��>o�zz�j���W���{�~:��'x0~��)�3(r��7GΧj��W5���
AjW{n�$C�+E}#���LF�`�,��%�����c��.%���J|͕���c����J�ЗI�j�
����O��UB̝��~7B����Z�J9�ׅj�o���"?IZ�qO����y`��i����ٳ�/��), �S���c��=�p�_�>��,���z�Q�,z���U�evLX��޼�v�Np�f��ni~���U�qxr�ے䦄�Àѽ'C����ff���v�n'*���P��VZ�Y%q	L��.�G5������Bh�Z���?�M�^�*~� �D�?�+*t��-un�Q,�D����!y�d���.���-������Ҋ�t��/�@���AN�r��,44(-�����Ǿ;�N	��M?&�*������"��S6#�r
�����ך,���f�����ܝ>����胡8��0�B����{����>�X�������������r]�~bCsV�cI�!����8��.���p���ݪO�}�`�C:�z;Yy{�#֬�"޿���v�,@~@��)�"�ZiՁ�Vpp�����|��Q0|�A�R��x�����(�����ϳ��nzã�B��P�v�F�y�^�i�-6�&n�V�N2��O���F �v���IP�,d�GDV��@����=J:�Y؜�Ce9��k�E�9�c��e�Y�I�Sڂ ���WM��)_kbN��HF���y��-�����+Ψ�P,f8���B�v=�4��GG�sؿe�/�$���Č�Yp�KK��T=�Z�$v{]��U��=�R��	3��6!�}wo4�#�;��U���Z�r!�ؗU��]��)�m|���;y`;:���$�̄Β���Ax���j~~C҄fj�N��
9y�8�QA{m��f�Վ�*������ ̓�@��e�ju0�!bԁ��B�K��(@�PR�l���
���� 	�~`7h�r֙�\�8r�5�L����1�!�e��,3���C���N�ِ�֦=�{AG��9�ƞ����!05�(�"SE5"�K7x���֘���ƈ�߿���"��i;�	�g�P��/Z��R�?�뜽ؔ�MN�D"0�� \�Pm��1!�;�
�3�M��g�7<�9���xL�MǷK9۞�M��v�����-���R�wu J�Q$��OWE�ݲ%Q9���|�>K�Z�ҏ���0i=V���~{"�O7o��sV6&���i���֎�e��V�?�p�`ԝ������	����w�8�"�h�� �ݼR:O�w�.��z�;�OF���ہ=�j�P��F�`r4�^2f�f��¢��&]��p�a�YJj��r�91�
���ϼ���b���u�2jj��m��t=;?�mm�V#HD�ڷ 6�x��{a� �w{���r������F�����7�\x�M�ɫy)iH���w:IJ~���L�^�I[�K$�^�=�0�w�{�		f�{���
����Q]��>��F����=ek*|J��;by���A�	v��Z� ��zr{��'��1XXC�&+�zrڄa+����`a�݇��,U!(Mף���{1�^3!�f��i<a�?K��5W�xo�1m�\M.��0����S����%��6�Cs1�8��}���-@l��>��B����#�qJc�%���e���xI����pɴ�m�uI�Jx=���Q�`L��rH7�C�ֺDb��g�k�
��;M�C�~t����պ�#�[�Ok�K��"�A��?�Z�|A�eLcx����e�-8a__�u{�_�C��S�pfʘ�G�w���:|����6tl�@�>`J��W^ݖW�|�����tKk�����Jnu^?�#�N��џ=�|�
�����U����GH`w�e':!�W{�3n���H��-��B����cc硗��Ȥd��Q�HAK_�,s�4%����v�|p���膮���q'�����3ʦQoT5FX����Z]�(2�Bx�biő[1���Ia�xt)lY:�ߞ(����s)8�i��M�?��w
Z�ÆZִ���+��59�?�������d�W{�4������G�&��>f)P>�ᯡv�O��46Dn���E�+�s����	!l&܀�
a�"�v�0�J܋�G�J��\����:��>3p7�柬�H�İB��ؓH[�����y����&�{/�ml� �'���_ߔ�Z�D���d;������V�Kz�-��8��v�N���[���\��M�M��u+E����ˮ��T,�?ѻƶ�ç>�˞>�M�b���IL�\���O~��q;��5C1��,��f2a�>�Ǫ�~�|���SE�L�?M�c����˝/�js�Fs��˚|X��]a]�"�ow��vqG�-�o���Aej_{�tsp�\�U�V��OwD�����:2��['�8��S�|b�O�W,�P���;fZ�Si�?&�L`�+�so�~,.�oz*7�AVL+#p}��e�J����7aXd�Aj��rh2E�\��2���.ݷ�ytM7�0dn�2��t[8�7��� A �7�Y94�a�O�"��n3// �0�3z���f���2��&F������b��ݻ�S�F'p��!���>{]�h-��Z�E}����ɺR:OY���Bqj�4�]GL��sN��LP�4�/��vS6.u�{r�g�Pu��C����/�w���noK�T�9��;�T�ʎ�)-���6�4oWv��=N����`����L���5���W�0?�@;�Z<ƶpۼN��*E�n��j�"e�Fʙ,!Lx�l�oƃ����ٌ���V:��\c�7��%�r��ԯ��
"s�ֻ�e�B�᮪�ᤒ��h8?��#4����w�Tp�v�ړUm*l�g�H**�<+;T�y�$Y�Q��uNo[%��0nt��o���e�n"�Z<�++Z�����:]{�Wan���#���\���P��E�|r%�=��'�~�qT��_�,L(�������(�vq8F�����Ͳ �V�W0Ҍ#KMM��Q������E���L�n�Y�:?�����r}��W�V�-L}�aq)w��!9���N��|>�籌ѝݏ���z�e�u���25���bbVe�?]eS��q���DN@�[�/��x����7È]t�r���s I`,����16���|z�0�	�9
ƫ��k�V\�������0Ll6Nm
�T$^��v�U�Ub@i) ߭2pZ�E�HH`ZuF{!��<D[Mă�����OR�V�)W����WT�U?�<z���
�#E��ӴffJ��&����A���ۚ2ߺ�O�l{7���ڨL��i;�Y�!7�����l�{��->�i�J`�e��)�͇JRADDl8�\[�jk���� �	
ƹ*@z��"�-�x��HX(��>�rN�wQT�^�
������)-Q����dyώ]��ӳa�Ѕ�|�2 z�nba�eJ�%G�6;��zކ�/FB�ܭ}֖KA�nPg**#��z�1��p��P����P}�oo�Gޯ���d�t�R��
�й3�g�̖W̙����ƿ�SV!P����o�VZ@E���ۋK�&e�±��OF�eR���hS����?Md'):�v��4Q��ɔ���U���ѠlrGa+rJ�̺.%�P�1.�L�l�2�:	��T��+(��x�	���v9{���6��ü��k?߸m(�[}�C�*���1��j�C�4�d�����|w_R|����D*�h�I�m�hO%1ѣ�(�͇;V*�8�gp"�ҁX�7��D�--ïmO>>
�21�2�A\��Ԇ]u���J��?u�2`�]r ��^���"��RBK��_in���C;�@��*�9��L�O�		���2�俖5?9�0j�����g��)�W7�,-�v�I1a��k�֬��,(�>�p�޽��C�V�V�isSH��,b}ɤ�YC�7 ��Isaj�G�ٵ����0)�Ej�𗒇��ǂ��^�L|%�,G��]���[�,;�3�Γ��t�G�-eō��hڶ��j��w8"�4K'&"�0���߳�J�}�{�h���thҭ�M[h����4������.J&o��u5K�p������^�<�Pe�`Z��t3�.Fi�Ek���o��hi���
��Y�>|PPT�����(X�Bp }��[(��^�ί{]su�Q��������"��.)IsK��G`��̒�qE���*+%<�2�;IB1�K�\���7�'զ�
 1C��5Ks}��us� r�r����NI̦�NI�R58��A�Yt�Z��������יضh�Ϋ.L�Ah7ߥmr��H%�+�]E�S� 4R���^Ӊ�vj��+z9,ٓ��'K�����*�=l��N���E\<Р^���l��?�p�|�5\�@j�:ɺ��tD2�U2y��F8x�c���e��A44^wZ���g�";}�ejX5�ynަr4q��4��@�o؉����l�,4�"�<�X�1U���8��D��dEoՀ��K�X�3�cY�|��L����A�]hP+����k<�G/��K������^/NQ_�X�c�5�y�����>�`�Kޝ�}��(E���nh"^Q�)�.�ú$�!u�KV-�	����ݗ0��nk�xWy:�x��`?Rt*���~���r4$�]�c������ܶ۳T����.�B�ͨBkS�&:�/));���#&�T�9q)��ʼW����cє�O-�V���������i����2r�۞�ԗ��**�5�Y=� =K�є��E��H���Um��fV||>?��Hs۞N�`ݙT*��2xjWmf�zԱ�����ַ뱼O�R	8\)�)�0n��|,�-[�������5��(�Cӎ,��ٯ��[ @Ȥ�eܧS�i�[h��ˋiyΫ���ѡFFM�MFi镪>�[�?<����xw[!B ��t�[4��&��ͬ�FtJ���������h�7���q�ʖ18���s|*p ���s����b�!UąA.-��Y��i�+��Ï�-J`�&�+a�ZMϔmg�|=���L��N�ൕs�������!��ɝ�|�����֚W���rAd""�	z@pv�wm��	3�'�j�]��6�+@<n��)��by��zd4�EBW�����v?�>! �lZ9Zp���։�����~$�_�r)�Z�߉)`bg/�.-��bVP����fqR�ǀw&�˰B�Q(���|~9��s�����GƳ���t�$��"51Q���|8�7vA�/f�UR����vM��+��%q�C����O�2�j� �N���� ���L��,�Z;������Y ���Gw"KiJ r"� �UKl�3��k�-i�)�ڷ�o�����'�V�K���I����.F�弯J\m��~��?K�EN����9�V��¨@���T껮�wӷ4��y�
�HG��@�~�w���z�V���.��L*�:ї�d�]��~���Jª��3Sd����/uz��2�R.{v@7,̩�.ts_bj��gPFЋ��(���de�=Wb(�Z�̴��*d��=~�����/D}%����Z)_<�e����p��$_n��V�x�~�����B
�7�N��,������1��#1��%�s�����H8WY(V�0���w����쥨|�Q���l�$񊄬�/rp����������7:[YA��BI���� �=(��J
.>�pdD�چW\m��'J<l۳��~�7V����iMP$(�jKK�E���W�QR�ԩ���iġ�	��u!��2��_Ǎ�8�� �s~u[{��4hqj�	����ul���'s�vϡ�R�S���,-$�jG�5rJ��ѳ���o�ܭ�Ot��DE�/���ZJ���S�l@2�$�	o���<��7��>q�:���H� �4�DOK�K�r�NV�<n����9B��CU��1�u9�ǟHJA�� �q}t?�ç�3^<���ݒ�4��������<�W_ܯ��sM���*�����2� ����N!��/��b�1�����׊X�3����m&�Ɩa
�3�+�)�١Ӯ�������SzS��;j2<���E�~i���s&�E��PT�`]Q�`'�L�����XJ�_-,ʖG��Rɏߖ��ɇK�}8b�K�f@�(���Є����.Y���^`]?�u9�/����	^o���1�F�ӾRT+#�D��n�pL��h��g�Zi<�~�F���A�.'�k=�����v��]}��A^�&��g~�"i+9t�v��q�z&ŋ�:9�\ۻ�>������ay��K�y`9��0�-���d���뙼��f�99��ʼ��:#�� =%�iK֠,\j[�dd<�Y��*ڮ�I�sa��:&3���Q���T�!2i.��7y���IW�.W�y�������XZ�Cto�c����H�z��޳7�Ásۦ�X��k,]��&\����-:0�
�zO3+��h�i� >P�����e����K�o����ڧ$�Kf*�!j�E��e�E_������g� ּΟ�@�|;����Eg�k�Uc&����V'q���4p�M�:��+��ߣv��zW��\�B�\�
�S(˶�SP*h�M $���5!/�;�|r�[d:CC��l�3���W�%�b�� �}�����̝G=$ó�� �u�#3��|}A(a���p���#���.��1	/�t�e�}�}�G�ܹ͚T�6���.0L�!Lm���U3`��W� .��j����^s���;8��¹O�Lk�=�u<Q�z����>�]��aV���jy��	��4��=�O��f
՛�چ�~��M��J���H6J{U:�F$�����$F�H���
��G6c��L�� ���}��NZWΩ.r���RQ���:p��Ǯ��Nm�o�<�>nq)�Ғ-�k>G���w��Ɋj�d�=۾ڣծ�b���Q�Tp��7�>cھ�0[ay��J�VT�,yY���[�R㿽ȍ��׬��if5�R�r{;�ՕI��:�պp����9:�x�g���<������e����?r�%ŋ�H)�2k^���5��K(M����/煊"7��y�-�����!Y��]�浛����uhRG�b�Ӯ*�2P7٪�NI�����w�m�,i"�r�[��[7"��,�OZO��o?���٪�x�-�!�� �� H����tw�t))%ݭ�tw7H,��]o������fg�w�眻3��G�	�j�����J�(�ɱ��"&],,�0<�E*�~��������� &��)�L˵����gl�<�'6|t�w���Eb�=&�3<	�]
W�m ��1�%��O������1
~�5~x��mtH<�dz���}-z�.�f�?]\��՟������ک����q|&^�qT��V�mБ�LVT�)�quJ�L@�
$��B�"Zb�wȑ։�c�T��� =<�MϰX9������	K;�P'\�E�i���M]^YÇ=�EDd���#� ��}b�t�/�����a��V�+ٗ�-	��;��\N�Kj^�ly�&�GG��ʝw�rG����f�bM��g��'-���4NR��(�F[[k@�����e<l�\~�")���]�T�}�����٤�$_Ԁm(���g����J���Z|�U1}MW۲;�ە7����5����#h�#�PKJ�w���:N�f��T_�X�(�݂՘[����/���K�**o�]�e��BS��K���ZYY�(a�Z������_%��gX9�<l����c^^�*��̏�s��8�XF��8�Fv xg����r݉9��.}#QF'���ޫ�Mʹ2z�`Ä́��PF���?;Ĺ����8mŀ��p����	\f߆$k�4��~ǂmf#�w(�&Q�X�0�JCJ7-��a%IJ��ޠ͎|}M� �Ƹ�3$��5��z*O&SV��zp�%� �y��T����K��S�80�T��N��g�l��32b��)	8"�s������- ��5�h��4��뜅��f���f[�*"Rc�4�0C�nm�V�b�h^�ȣ�hy�^����]P�";IF�=��8���V�4ˏ�ζ��31�g���tzY�Q����&��c$8�ŅY��-_�Ѩ�EDGkkzhb�!�,���ۡ���i��#2IA0��nM|�f#	��hP�D�d>
CiF�D�%��;|�\�}���9_U�������T!�%aUe��t;�{u��S<0�
1X���/g�8J���\b�;I*�$��3��2%+�"JP&笞Uj�l�TYo��S����T�����^/� S�� �49)��2뮑���%H$���;�QCA�k���uX�V�7\԰�N*ϛ���;�A�V�ѲA�սV�i��m�&0��aMTaICF���4�w����W��;P�y���ʹu��)�B[R�?Q��N�!­�p��������ْ+���~��%l��ƕ����B� 	��E��6����Q���O���T'Һ1�^�p�`�m��r!�,y��A�p�bwI���#�??�-N�ѱ��N��u�W�fX~n1��X� �}9����%�����ҿ��E���v&^�����P�.KPܼ���'�d>�}]	���N��0�4���p�B���E�p��<t�0�������onn����mg[���Iﮘ�"���w?GAFqh�`�ٵލ������E���
��~I�8eԽ��)����d����%�E���=H2�u���pT�m~P�(����I�z�&���Z�v�V1:v�w�zS�a��,q��Ǐ�6�ۭ�����o��S�/w9H�9�ֶ��I^�$kꆚO�0MyeuJ?a�rD�fW?�,v�I��vĕT����� ��.�^��Tx����9!�r$a��tډ�Z}�`qЋ2G�}�`z������m�lh1���d��z4���fE�ٱgW�̱�d���F��_&��<��V�΀8	�F��j��E∁�l�d�9eu�Y�AW䤂��ܐn/n�1c�˪����C6��LN�GX�ǵ��ş�f���oPp���o=,J^��yx�0�3��`�a�!�[���|���K"��$����m�����X��GA6,l{�l^��r#E�ؖ��2��u�נ���٦��*�Vs�J� g���<�+f55�/��AQ](,��Ua�Q�Z�(�Bc�	��5@P�䢞ŧ��ad3pP�<@��h�	����!���d���W$ʜE=�O[c�R�Yi�����w�z��Q��51�~G��E�)3є�(�!��\�xm�&�d���M�;n�xV�p�`�PǀM��=��O]�F�E�M����p��c�}��z���C�'e����+O�J���3	g{���������`�,����l�+y{ KD�.�s-��]�y�k���q}�jhqLeǁ��H{E5�������� #�/�ҟ�WO�%�npr2ǣ�՜�H� ێ��*&s�{%e�����F6$���_��I$W3�E�^(f�=�}|FԹ�M�W�q�Ȯ��:�"K���N�����"�]uKl���8�*��F�Ă!��q��q��,�:����Π��=�Xj�ܚ�ڟ����F�{�7�%�g�[9j�M&���G+�������ې������
��{�Y�j��a����i;��ZJ%A0�ʀv6���s~��7z�N�*���?�NÆ}f�-����1p+��iǵ���f�R\D"�@��짬L�EۿS�`$�ue��6�* 5�G�=�`�����t�~�Ӷ���˘��L=�S�g(�W�2��}/O!#RA�!�V-g�_�q��o���Y�������� S�<��i���?L$cu�@��I� ��1�
77�?>�v:���}�sl��n�����a1�t��3�cˏ�6�*����#]�'�0�]�*��zY"�L�Í� E#���>[�4$o�0�m!+%�)�.UH���K�3�04��TF��������@� oX������-u�+(ɶ�Vs��Ųt�]��ڜ	�A�V:����N�-����Gב[���?@�։l�O�־�?�{����N�"�"�����x;��K���^lT��� ��.à�1]n:LP6ݩ�Z���0q�ᄰ}'�L/����AmU���]L�L�ݫ�Yj���04�rS(
�~�p����6й�_�D�P2�1\����=ƅr��,H����Q�I),¦�p���r
����j�$'��o�WC�o�;9�a^�Q^� ���N����j�(y{]�χ�22�i��Y���|+/�+۶E%���Zg8������w�q-�u���h�G_ʗ`�an@�l-V����:���}���$���c$_#�i�#]�?�h0���Y:�oV� 0�b�$�&�Qo��GFm�U����1K`���3I!��N���o����Eޯ�B�T�ǀ�<4������ݫ�j��B*����ɌGm�AP۵�z����P^Kp˵�H}���W-AO>��o��X��ò�o�h����"���A��f �r�S>vl-g����&���ň
���:��h�m�͛�<\���|ϗ�������-�݃�!1p~�S����־Y��c]ȟ��gf>�yc���~wY]���śW��kh�H�f�:�n����CQ�LT��������[�!�cK�G�F�D�։�����&@q�t�ς�Χ� �]�
H:�J�㯒��?��k��Z�����J��[�����Y�g�&MӤ5��Y(�-�8����_�`&ѩӒc�$$ba�̰�mo�v�/�M � ?��y
��]*%�;e�ioK�Y˥$Keyy�$h!B�G���#�z��KtGA?�/�UЎ�V �t����4i�o%*Ąo�g�'��89K&H�HO+X$OJ�Γ�J�Yt�@4�s�7)U�y���G1�ۄ��?�u�ml�	�~�������j��0 {��à���f�6��=��?,�z�To8�)�;l�C���zUy�UP;c+��w<�+�a�x�M���3<���#�Vǩ��4^6�G|��q���|̃)CH		�_q��B�e�*�X�����:�gw�E��'b�2m6�0��e��N��<a�~��G�?���[��Bu��^Sq��o���*S+�3�>n�l�V��jϫ�ȧ�����"�8N����ĸ~�6����+�������%�]Q}vӌ�5��DE[7xX$~jt�U0Mΰ��p���#x�\�g�����I*���?{���v[�Q��cVm�z����=bUd���ܨ4�k���b�_�Z��&%�,��)D,@������)-*�2f�����o��Pו�ʳHy_u��P�.����d�ĭĤ�
E�<f��[��[[IaE����`��o����xi�Z8�d�B�D�ze���O������G��5�����V�i�z�^nlul�{0[�
�07_ǖ�M�_��kk���rp̿-��L"o����� �G�����t��M�yl0n���>/K�g����1�H�"�{a�o��8]��>[^�k��sB8��[�n����A�1�MO�o�ۮE��V^�A�� ���-����fIؗ�l���5��Y!�܅m�z�$@�Da�\R����I?%��Dy�o_0!������uF뗩����]=�"u0�f�%��=�"�_FF�u��@m$l;�+�!�/b1��f{U��yKkJI�nm����,���K��;�ëQ>�6Fzkݎ�R��"�+���nf��Ʊ4
9��lA�fzz���`Rߡ��B�`FG�z�c�{m%cc&֭��g��no��xB�1����Q]��:�8��_:���:�"`�o��4�m6f犒��j�[A�*gY}��r�����̾���Jc�͂IEU�Dk�O=���P)�T�W�s���w��*�cg�?�	(.���q��U�� �����;F/�N���V�Bg�FwUNW"���@�(�]�4� =�:���꟔WV���m�,����i/�_ �׮�X�}E�#����d��g��,Dj�1M��I&T5�ƞ�x�[�l�{�p���)�9�)w��k(�:}��')��]EفJ]8�2�Q$��&��v������`���Mv�c�Q�[a�灛��-�q�u�@+�����auD�0YF��b1>Z*�� w���U�}���y�w�K���	��X� ����Q��-ŧh���7��
��{��II3��_�������y��'5�����]����ۛ�U�ʁ
8(�~�l2�㺅o`N��d��/WJ��o8K�V��D�&:�h�LxFq�H&�,1��7�ʱ��	c[Q�����N�iޓ�6�0�\��[�b��{�۔o��\��f܆%w*��]	����3^��l�ӧ��+�z��ᙷ)�
�f��Y�Y�yG�RO��D��W�`��ex�b|D'��򽬌��.�ߟ�]{O��@��#���\����Kt_���ˬ�J^@�K9k��� zĠr	���{����7Y�hJ6�^�>W�L1��֬�O@�W�l�OxP������I-B����-~��$η���P�V�����G����]J�����+��VX`)�"-w�і�eoh+����Hs|Ӊ+:v�bn#,t�ar<�E��w%�;��u����C˩M�MB8H9{�L�PQ�mQ<Tˊ`�<dG[c�t{)���t���Y|�1}�ﹿ�q� ����4u�$3�	��7_�Ye�"�Y��>���è|���c��e��e~���ɪ��B���_��Y�,��b8=.���10I�մa�����)���/���,Q�ཕ6��E����],�K���q#M�1��l$�ej�nN�o^�Ɖ����A,F�h��>�A�+���N�z|�]���V��T��t�����z��ܜ���}��������h^�������R|��S4�j�+�������#���)�\诖�,�Z6<www���6���	utw�`ea�x��3~�����U��T�O=L'�W��Z�()���K��ΣϪ}:�SlA"�6�I�B(�ڦ���k����IѺ��W��z�ۧ^�.�$4��[MbJԹ�הɦ������:�m�Ր�Ъo
1����$���Cki{�0ޠЍ�uژqd�Wc_q��l6��m��ʩ^�KX�c�'&�L�p���GN�h�S���g�'vǞ�x�1���D��]8Lb�֣6k��"�l��������NϜ��~`���ɿ(��%=�/�I_ѵa�#c�	�<*�}��8,���E�WK�?#�,,T�i��ж�J2��H�<��MF]���I��5c��ݢ�2���o��ud蹒x�$�օZ_�����MV1/�f#�(Ty�YA�\���)P�Z`a#�:�\��4�$|�c2��[����+�ed�S
�sZf�'�����}��a{�Q�dXsҴr�q���|q�r��ɝ�6��,�o�xgX�|I���W��p���2i|�q�~y:��p�v>�1�Ծ��V��zc�\D��==�(YY�_n�rZ�8�x�&f�%Ti��ڢ��m�B��}PO6�ݼÄ��X	�L��.�r��q���a�e�<�H�������E����'��kh�O%�|ű�%�9T���@*t���a9PL�9^)��uZ2
A��O2��G)�E� |��}f��h'  &��SGkT�G����]a���8��Wo2I�i��<T����q�!�:�����7ku �t��N��g
^%���v�J�_��k���`�O�]᭪Y�jqԼ���>5e	�O��v�p����Z�d�݌s��_Ί�(#5��J������j�7qN@|�īF��!i�ְ	n��y��)��}�����谟�Rs(����F�����:����9�h���N��x[��6�oHJ���ay�di��Q�}r���-�����t���,�Rn������|�a�_������oYq�vޏ���Xƹ"��n���<���q�HC���XzG;v�����p��ɍ��%�����h+���ez����^����@mڞ�T�F��8~Sd��{��y��'�:�:��}�t�io��+}#ֶa�/�@׼郿�^Kks~�q�8~1eM���Z�yE����;P
ן�8$+�8���ڍ?�k���<��"�~
M��w$U�G����P�&�d�˞;�%K�W�k��Z�]�3�<��*�\�K1,���	���@ )k��}����5�y\��Salf���(8�q�r4p��?�/���`űw][#��.{��~�*�ozs������b���T�"t�E�[�9��p!����D���d��ar�Rr��hA��1\�Z�����3�?-E?|�sxY	��%�"'h�ѡ"��p�bk����.���c�[Dh��C��63>�����Lԯ;D�#�cl>���|�*h`��bʉ�/�{�oz��d9��wc�� v��m�U�\ ~G'��V�M+� �#�@I�ۣ�#�����^q�kT�
�S��]��k_Sr�'i��p;��]���
�kjS��/�Gŷ\�<��k�<z�@<`l(�W��G�o�ʳ��䀊f�~U�X�|��Oo;�B0���_it%�o7b���Ꮵ�oj�Vޜs���*قa�f k�yP�aČ����� ��@���'��82��ށpc��g�/ѐ�g�s�x� _g��:*jHȼ>�#��Sč���&�a�/Z�mqe�A���L���x�5�ߟؾܤ��Z�����)��B �$X8te%��'W+&�R�X�e��I�ζS����I��H�+�e���K�D�lM�������rER�߹|?#�o�@ uFa5�c)��;O\�pB�sR�֔W!�.��+٪_(���*&���Z-H1�*���-���^ ����c�gt^|�����<��*ې��H.jt7\Hy��SVyU�������	�w$��X�����y� Al�ğ���D˨�:ː� r�Ӡ�9�9��nک�-��Y�Ř
48��&R��Qd䎖�9����^~��>!�SG�K�kWJ�?��J�/�K�-g��th_�o@�g�����d6����"�ml<�q%��W`�t�n�`�J��;-��G�q��+�C�$�1G����c�3У^©6���M֥1��N���9Ʋ�#d�\�d�մ�M:�M�Cs���vO�0��wue�7Y]r6o�I޿gBE�C�wZ×<���}q��P���@���Qi�ӎ��.4��e���y��L�pl2Ň$�(�p�*)�S��z,?m�쓃�v�:�wfg��A'gL����ׄ}��bmc�|m�e�#�5�g#i$!�ӻ�Ea�O� ���DI����
�d��s��y/��"o�{�'������=	���)��5�<���$G7]:�����=
ćA8��&!b��U�L�z�/(뷲�:8��F��NКjw~n��&9��d���k�r����S�g�O}�6����Η��QX���uO�^���Q�=�O����[n�s�\�;�'�j��1����/�&+(b�rO���#��^��Օ�[l��B���@�e��Q]���/=#��U8f���-3CÇ6V��c�d�#<���������X�;�;������|Z�Eٰ��ko�軜��=���������Ԣ�J�
z�����6�5�d� �93l� H_9� ��Y�����æ��+.!��+�ey��2s�2��0�]*�졅۹5g�OW��.9�!��}��g}7�ʑm.
��b�;d��n������%�D;�ӐLJY�p	�iم��e�L�A���ƥp�v#��ψ1N��@Zp�1B ��f�t:\!��ck4����5��(<|��;�gD�_�`��`^n
��i�5=�j��ۋ=n^�u���|�84Sb�����r����A=UGtĒF$�T�&���.�-��|HM��5�N%�fN���|���	�Ȳ�����OΌ�M"X�,66GtI
,X��[�NMGT���XPmq
�$y����_;!����1xV��9;��b�v�􏛸�4+�ٮ	qCHP2D^k�3�T2�ӛe�a9�[Ъj�GyT�[b�4�2a,���Lδ��V=���--.�|*d�?�i�s��������p]hc�y��n���.�[�{�	P���EDl�1���Qz�ǝ�S90�w�l��T[Ƙ4&��[���au��vj3]�S��I���(�}9�	�榆����I�9��v�c�L��=��T[F�b�B%S;?®�X��U��l�RG_�)��%@�#{i�3�&Nq�~?����{;�}i�7�_��n1���9�b
x�to��[�d�7��SQ�D��z��;�<�8��}�ށ	-D4Z[0���G,�B�7�ҦR�sl��p�0k팖�[uW��S"���ƘXz�vW�5ͭ�w׌��5�}>����e!JzQZ�~$�B��0�w1�ak_^��|3��v�6Aɗ^��n72x�o��:��ht�xg�>ȢO����?NkL�[9 '�.k=IHE�o�:��%�oC#�.��-�B~ۆ�QR����ƚ˽6C����qh����d�*��c���	���i1�y�@_Iڒ�[sz���V��|I�T_A�m+�yg�Q$S�׻��m�MT��L����xпL���ݝ��#���@�Qx!�s���<Z�vP
\�M��c��Yp��HzEn��\&�u+;��&����1�~t,9��X)�E�v����7Y̝ʔu�ܲ�F�9�Q�:EZ6i1�~��h��Gف"������8v��N��_8�"�c�v7�G\���!�N��u\�rs'p?&c.	�AMWnŞ���f�+K�1���A!�a�S����dpz��V#9(����K�D	����,-��^zeJ�Хm�K��v��6�e�s��t�x_�N�_T2������w�HQdd0;l89p)�U��*n8V#)"ڸx���^��C ��hq�5(V�]�K����GYMu���h�ѭ8tc�`zb�;5����5WK�����SQ-�i���q��w���P��Yh�B�G���T7���uǊ�H00#b
���s��zd����� t���L��蹇���;���Ij2HBkLiF"<�;�Db���zN�9�kl�������S�r����ꙣ&�~tL=C�4Z�~�M���r�����cEX�>����h%@�ۃ���鴍n�yo�>.�_1�ٿߩ��?�$����B�ӡ��&�q����
9K���qG�M�$a�w�2�7�������b��I�˃����WfD��2u2%�
��w-�RW}ň�xU����:��r�*%Ps���-��r���m�4/\���eKp�Q<��D��p���ƞ�9&�L�|�|��N��CHg ����BB��>�����M=+0������,���A��Ȯ��O+0��_�&�?�ݶqi��>�	��,NkK�Nm�����g'p�Fitɣ�S˶1��@3�p��`ǘ�U�d��T�Gؠ_�W���nb���#.*(-�k��3����j��#T�����1�ͬĂS]ʷ��h��Qy
VX������xą��*͗�}^A5�����`Q��ȤV�1���f�Mw%E�uQ�;�<�Fn����L�nV��J����I������+�J���	ʲ)w^.^���OL�������r�ȼb�N�������OPt`C?��9�Y؀���������WH��)��@o#'rЊ�������B���␿K\%W�ل�/��]B�k��I�|��#�Vp6�����ר�Mڟ�\���a8�Ii����
bq9�I�Tz�N��]�֒�O�����%�~��yZ6�n_���H��*��@�$�]�cM41pZ1�Q:WE�1Z���4\"D�<h.�dk�w�{\έ�\M>>2t��CQ�W +a�p�5�ߩ\c�6��4�P-�*��H����3���x	�/���C��aJ��b�D�A���@�))�lp�T�&��8Y�L#�˦��qRv�f1�] \K~�L����x�����TЃuRRz�*ޖ��EW��X�;���2���<���(�\F�,�y�*��� � }iuG�����`���:��<D*����g'|� s�`�6d��
� �+�1�;{]!I��jl�8j�:����
u���b�';�]*����Z�9�|&FE���@��A}S$U��\_�hB'#"$�©FZU�L��w���KҔ+����K��ȏ���t�Sy5Mz"���3)}p�����::T,����䉀���j�G`���W�¥�|�� ��%�+�P����T�MV��V2�t	�V ���ć���	��N����(�h�h���̢�T��ce�o�U�8�Ѐ[91�\�A�E�pA�5j(�:,s���0�����Q&<?���#MS|㩐F�����TE���?sӚ��rPHl���k�t���C��n>z���wo{�ΈJp��\I|d�щY�r�Z�U���������(����eR�^Nչ���x�r�)j� �8^��N���<�ο��2�K�0
>-v"(�E�k������@��^6ܙ˅[��n+��=A��-�w��8V�~G:��y�jKnH>���Ŷ�E{D؝Mj��N�[�>|L^9B��t�M,�n�	�E�g��=F"#����LĬ)pz�Z�2��,N9�y�#������$]Sm�YXK�ס��+.a�ZZ"�>m���-^���"�n�p����Lݯ�
��4�Hi�XHj�ggN�5���==#��%[+� v�/ ȗT�u I;� �٦O�5�7L��`0�>~v��~*��~Jj�Ka����@1B���i�i��:Y�ޖh���؅��x�Z*���9�I%�55R�j�up:�����y��k�� �A"Z"&�2�f�	������r5�컶���k��Ia�	Scl|�l=�An�.����:���	�0զ���D�ړZ�F1ŀ�ü�����b>�
���JEi��~%7����oq���P	���5�.{3��??	�\�Q����S��+6��D^���u���h�pw���X�� P��,�v�%����Ϥ���IS�r3Y�v��"Ɣ�����7�E�&�ԠRQ���8�i�v�@��-?�;��1x��W�8;@��t�y1%F�n�T{С*�ЌG�$���� q3�h�k���^8��	�`(�}W�O��K���?�*j�R̅ ��(�^��e�
������w*����#>�4��p.��a�ϋ�F�8O��(/��_4���] �Y�4����I�� X�
gd��V	�T#G���+B|s��1l�W� �t^�oZ-�XIr�l�Ty5A�җ���L��Sy����OM��4�'~��)�G�\3�_]��v�����\�q���h��&��me�������͵���J�!�#�,}�d̋n����ĒW1.*$� ��:"�޲���|��+��h���k�}�7o�x�ɴ�����ߦ����3��ۯ�^�è�cj��B�l��,A����[�ykK�#FF�m��u7B	��sډ�2rK��N��O�p&\��¼̽���M>�JJ���'��>��������s�4��7�P�4��D#3�{.TB@M��v��h��2v~���tD�"�k�2O�$Y������e�X��ylR3}2��L�?��y��X]�+E�?�a7x�JjC��Ġ���4��?_f�S�H�Su���� 5/h5��D���W+O1t11q�g�v1t���Igּ�D�j��U������։\� 3^DwK�*���45��=&��y�@�5Hp��)1�������_<��+7�x�K]%1�"M��W��yfE�<������_ N�~1���˓QRi���^W��`� �hƩ���:���A9ңn:��0��� ���A�}Ӂ �D�$�柌M"*lN��w��!�T�O��bD�Wb�!Ob,�8#o8w#����v�}+f<OB��� ���3�H���gܭv?��"pL�<�j������,���%�H�f�8������Њ��%�5�p^���J�Kc`ً�]➺eQF
�
����B�.q������#��#߿O��[ƥ�7����d N;���� ?�xVڑG��M�G`�����7�C�80��<T���.���ԝ���'�E�2R�)FX���v��]��_o`���ё,ů���	��-��;���X��b���"��wN��N�鼣W�a�`c땿8CdG�n����kē9�E,7in~�ʩ�������Z�����,k�G�ƵJ) T�3=�~�S3P��]����n������V���%�h��T9�V	Uc15��~��[���YfyM2�@�nr�YW�ƣ�ؑ���+@���H��vop��a�Z|���zɇ�bU�0�@���5�e�%.ya:IVڨb�5�6� 54^�KJ���pe;��&`��҂�@b6�.��� �@�~ю���=��ek�{l�kz�<��KSJ6<1��Ņ��C�y"
��9H�S�d!ys	�N?K1t	(M�곟e�փ�V	���F�{$�o	I�ޟ*%!��JC1:�9i6#F���|VZ����~�BH��3��k��{%��Xى�2`�,( �*%ր��Y'	��h����0��m,U_��쒌����E�u��0�����_e�m^Zڬ:=�L{���|��<�wL���I��F!�1��d>�($O-6m?�0+02��J��j��ܐ����*����F��}�]dJH��bǹi���Ŝ\�)�gY��#S�MMe;("��U�`V�29=���g�V��Xq) �c� Z�z�B���Wy��?��)�F�)~�T�0z�7`8��:;�����Ɏ�>|�g��!�}�?p5T�oj��:b �##��n:h�W�;�
�E*�����,ek�ֈ`�o^��Q�Qп1ڻ���JF���͜���hVG]���vG�{��D]# U�gΣ�0j.ә�ߥz��[���E�S��2�@�������5��!�=����L �2��Z϶D��� �$���!�� �a'�ݦH�]��*?����j	���>���@���*��ud��a��d�#~�UW�Y-5H��h�z{�����13!�W¼�|s�#4���E����.Iu�,gj���(v�4�_��lhUI#��[>��@�fʼ^��7�� �ß*v�m�~�8����q�a��Ф k���Q���(�ɪM�ֆO ����u������E)��n�H�eR��g��p�)a�� Gv����&9�)�����I)�fH���4�h���[�):��U����`;ŐO���Lp�*�Fą;��k�D>�RF�&S����ŝ�ş+����z�fpXC���Ll�$�ڷ�"G���966/�e8�&yHHO~�Gb��^���o��G;|�F6��t�P$C�<��Wyl�e�vR�^i.�g�c ��㭖���oﰵ��\X�U��J9�K�?���=vP̯����-)9��j��ئ��e4v:�g]�O�Mqd1�W�w�ur_��v<�B𝵜���;�Xrg��\���j��ω��;���=����V%�ej�:��������f`c��,M�y�YG2>W��}�PT�M-�lgy��s��\;l�Ou��X�*"�O���;g��''�� }$\[K�!g�Y_| ԾG7�g��A����+�,m/�큙��4l���)dU���%�Xw�"��:��W%)��-O���s���R+� o�u-8vY�
)��)erGF�����d� e޻�rƌ��h�M�R��`�Ϭ��~�е�PucːX3� ��a������e��xr&+��נ8Ͽ`�ʪi��f�φ�]��I/�Y���u�%��|:��T��p��,^B'���s��y��6�r��24�,}t����B�ο����î��2�# �e;9���(�Y�������qi���ݞ�|�K��v��BԚ�P���a�?�B @�4C�%D�N�4*���� y6=��@A��h�(��5w���B�7LF������Qӽ��>~N54����i]��t|M����m�W��XP&n�!����EV�ʍ�F�SE]\��?��«<�ɺL���X�M��K։�d��p�����t�;���w, T��"ux�p�z�~�^�R�o9��e�&(U��5�|'��#Z߽�*��7C�"�u5Sޠ�Eٞ���ciobUh3K��-�ch=�BwU`̖O*�6�}�s�=Q1�W4�a�^�X�g�����s��sϦc�4����3i�� O(0x��aص����5tWu�'����UT��;����Y���'���5��W�ON��;�Ql��)�$�gc�;͸Y�L"�-�T[�!�o�����<躼��k�G�����3�PN)r�zfm�3J���FG��Vt����7o�Cb(����mf٧�Z��qe�bh/��8�@|S7!�Tr8YE��%��������5N����Ϙdd���	MX�������(g��V�`��Rt�gw�y��:��{`3BA��U�e޹�i�����~�ϵn��nN.ֱ����=�������V`�8&�X���S�eqr<���T@j������Խ,�0,�]ϮǴO���	�4�T��!7N@1��T�yݥU�|�����\��$�A1��«��.v��"����{�$e΃�F2.N����W�Ы��5���5��2��ط��ZV�j�Ȇ��W�~�TIXC�V�'g � ^Dq8g
8�\c�d̜�_J��w-S$_g��qm��u���O��&�9�pE3��S�D�94M�Y����-n�"�Bۥ���"10��2��~�N���J�  ~��� ������%�v���$-7}��JV�����P�jt�����U�
��ξ㝇�4L����}!�4�Xzb�66Mv��+���ʬ��Jd.�Zx52��Аm�Ĥ)�&�;f-�+m�+~�>����;��CevC�A����+}f��lx���IR�9j�q,s�ڡ���BС�ǋJ�����~n�蓶e^]������a�Jx��hP�_����c���![$����ڒ�ۦ2�^n��f���цn�����9����%��m��t��k���f��E2����j�M�Gc6�=�MM
�W�7L�g�s�e���:B7c,<�'Ϗ�Ue�}�^��&,�v('�]�\��s,�~��sB�[�Q�px���/ Z�$|�n<A!O1;��}� ���3���Vq̫yj�՛Y"��/~�^��b����_�c(���
�v���3��|U0�����@>N��1m���#��Xc���]O2ҝ�RA�g",��PَBV��G���/';jE����'�g�`bȪ�[�e�Ӂ,�,��Q�GV{6�.�k�f�13 ;��!7�F�y:z��'�D�ӌ��sz�Cc1z�2{S�ݟ�!�
n��cܬ$f-Ox�aԣ+8|�i�7��z���'���7�3����m�'(��u�. �h1	�ԧ���E��ۥ»�!�Y�(��IV��Y�\��CkTQAʦoc���W�1�f��[��$X1U^-~j8y�|CYG�7	8�r�Yέ�(�~n�C�UG���I�%�C���!@�஋��[ �;�Y�=,�����6�ݽ����73��տ���n�mA��G�`��F�sC�+�V�1Fa�kX�=,p�XL��;h�1�#[�����Liy���kܳ�TțSR���v�~�Hy��l��E'ʭJ�4᝵�=�ș�ƒ<D}��B��~	NY�b �n�{��ɹAg	O���p�a7S;�ώ�rL�{�:U���
���Iw6i��5�t� �W��ʓ�̣1en�~� ��z��NUj��h&�\׺}�^�h�O��$|V�9�Q'nAj�җ�%;���^��n��<d�~F^��_�m�"��@yq�ԫ1SuK�x��,�4(�w��=�?}>�Av�tln :SÓ��9z66����] �֮A�������7���#�U�'���H
�{II�ݵ�DCG���	t�������-X]^W�r�H�є��1�1B�: �5,����q��wO�����S��%T!�J�sj�=�"��Q1/1��"��V褢#�@������H��TT1?���-�#��MC�1J18β[3���'�ʄX����Ӵ?<�^M���-�_�����ȷE��H�f�-���cL��;�]^�ޫO�;`h���Y����RҴ[v�;{��k�/�v��;��,-݂�,)0�~_���3���y������a�-<�v��t��S��?�[B���2ǟ���ba0Q"���I	>�^g��Y��T�^L�������{�� �[4��	�1q6X�!�K��d`|��iZcc�+���xm
@M	LϪ��|'�z��K��_�q��eE�~k�Y���û^��S�,�=���e�rji$�=�ZL� �s=U��
j����������	-�z�^# :d�g� #k���5���1f��'1Se�R��K΍����_ۢ:j�k��b��u���T�zW;����O�����I¿�����ThE�� 8%{ٯ�Ro�n:��4�w�)'��шZ�(���G���TeǢǌ�8H:�����	X"�*f��O�V1lg]��8=H�� ��y'�yF�7�V�X]Y/N�$V�3�e������
�+B�l��p���X�R��#?#c#28��N>��B��Er�>#�U��җM����O}l"^�HqJ�e"!RDX($��;U�bO�'�������=�x���.�K\��Gm�0�@���f,.ƽ8�c�X�UŚ���9�zp�Q��IF|�Dm����M�̦����'�݉�/�ˎ�-��-�P2����0�M�>�A*���Φp�~�`W��s�0��aΩ�O���7:��u2��(��Uy1�ǎ�Q�d��\~?o��5XwM��G}�lHIK��� �1������Aϔ<�������WsU���{\QP�)
�K�eґ��O���?�$��i�-
^��ܘ4&���c͆�U�E�=s�I��D�4� �B�����r����k�YԢ�H��BcE��,�QԾ�믳1���.߭ �󍖐4��'���d�/5��=$6H"ܜ��,xP
z	�k�=��{��_]*�� ��J�/�i�H����6��V��v���qGP0��&�������T�8�c���w�pCq �%OhH\��2U�&�&�s�:Ҡ����ʲ?�)�;����$!|3OzE�h�p7Qd��x��&�p.���� ����+�82�}��-��D�j��/O��QQ�VXzb���@�N`��v��K�wˤ�1f�5��ԤR$N�����"���]Ku�+�d� {>ſ�C�ã��T>�@�0A�2��r�'�Mx�_��c�RZ-AFh��yJ�G�p� %<�X�R˫ǿmqڍ��u�8POO�9ɗk�b�	�<��BX��z��7�L� �O=����zY1�}>$z<�̈́�״$$��^�M< ����K�6A%,<�:Q\|F�ǯhM,ۏ���^# 5��:ƒ�iǔ+�Źh3���Bk,���/��aj /��M��j8�4R�[�I�7�v�Ǒ&��cC�{}uBiT�Ɣf���]"OA�Q����s:���Ǫg��A�<�i�qcMt.�#s�G�e4w��uhEIg�� pa�p��q
�<�)X��p�Ut(�}34�q\U7wf�/**��G�5�P��$ȭ�0`8֧P;���4$M���4Kי�bZ�"��-�9����<�?�~�\�*��N��7o���>/��l�-�J����Q(;4^[�vQ�<�Ne�_������S��(*Zj̰d:@L��!��������b\o�_Y�(����X_̡,*
(��Q��ZQ���Ґ�V��ef�C��6�a*�Du�����MJɶNG��QNƞ�:�L�#.H���M�V
���H<�T�2�)��ss���<��<A3���k�Eϭ[6M�v�[�z�ׄ.��
E5{Ppy�Ǫ2d�7E?&�f�^�9�֥4�Jp�� �HMkA<q�Ê]x�6LZXHL�4R[i�j��_���Kw��3�(OK�t���k�^g�	Q�� ��O�1F؛�P$�T ��IE��O�f���$�Z�%;�u Oi�t��b�3Pg��{��!�@��غ47���g��c*P�(�+��UtEǰɶG��[�b�t���D��3�<���3
.�j��%\���� �ݙ�� 霘�ȑ�vcM�[/�+�I�*;�:��\إi��$��wAF)>�:��9$��$�'��<�U!,����p����b��}gw,�{��= ����$��w*�|��?����U�>Uq����G�[�L������(�P�xi,�Hd��
��3�X�q���������8&�0�F-0U�z^/u���i3Ai�I���%
0_ 9��(`�DHfɤ+,�ڣyT������<,�k��K�(+ ��j����OBfT�$?�|����4��7��^T�@B�Pgr ��!V�\K���ff�)=��EԊC��1>?t�>��m�2(':��.n��͒�Φ^n�ޠ�~��d���� :X��Ȥ�FK݅�Q{q��Ɵ�HE�����u�g�k��X�^l�%]��n2H�Ӑ�	�h�
}!v~�"=5<�+w�+*v�JU�V-�e&��/�M��mM�~���K������������WǶ����d����V̍����\��]���'0��l�!5�a�=V�}���=hʢ^�#��lMIelX!����y,Ws	>��Zt�8~���~�F��7�za[y�Vر9Y���شqf�3��>*��;��(v�W]��L#�W$����A�|�!�z�q��{�n�w�iQ&\{X�+"\�	ڿ"� {�����ѳ0W���W�Q7�h���"�k������˯H�IWWx������9!�w�H3���C3 ��1�d�7��n��e�ˮKk~ؕ� �i�.�3'ռ��#�)C����|��]����̥���|;��	A��j'�I9՞�dpty�n���>�#���ư��K%��T�
�˗2l�ߥ�}��W}���
oP� �������抋����ÿ�_�01a���=��6�JM�u��>�ul6��N/(���sPF��	.�M�fdi��]"�����kĽC}S���d�-M[�$]g_�n��+�1��b��'Bm�ú�s�t��o��}�	�[��|��k��OC�"$�����d�%`���k�ޮ�-ʞw$꘨D��8�?���Λ���,~F�EY�z��7���va3/�k�h=�il��U���y�ʀ�
�@IՉMVxCyH���8v�r2j=�Й8k�u)�-͋�$O��j�J*��4��S[�fc�r4��f����򣀅ILľk@�9O#�B��s����RNDk�Ou���G~�6���V���i��u�d���#ɼ ���i�������w�|>�ŜÝ�KL;?J�7eX���H���N7��S)є�J,�(���:�>EO_W\/�[�!��~�s{����]�$7�%������OA�́�~����p{&�''���[�;L+R\.x�d�{]u��n��WXa+�G�0��rO��ȴa����B��7��G
g\D�Ie`�+Xr�^�5�L�$h�i4�RG�Jb�'�m��Ґ���5�ێa|�!�(h�3��W�2�Zu��;�NAPN7e!�b(�!~'ϱC��^��ݼ��e-����+xrT8��޹q�t0�5�F��믴�6�,P~��U>yve2�NJ��LN��3�S�A!�}�"Z��|��ů���/"P��0�$�0�Xiowc^���<��z�q__�c )	/��$#�3�[[%aP�Z���T����\��7J��N��8�9��\������5�fo��SWB��2�,ԚE
���0B�֍�j��v��]�]�2�/�k
#F�X�?%"վx�G�^��_ȓ�R[����`BF�����������r� �����:QZt�PW7��B�o��.6�V�Ii��!]r"��r�=<
k�1xQ@�����Wҥ���ש�6��p��GL21o�%W��y=$��^�T�P�w6��B�H�+~Y���<��G'����=��'��q6W)U_h���c�P���YrK����>�7�U�'Z��I>�oi@r[z;�so��)S���P��z��A��<6���%���5	�뺰�#�����4u�/�77�|�������r��8`�1�7C�Z�d\�~0H�b~��:�����tGվ>hE ��j��y�N�`ⱗ��Ղ�BӞ�c<Ɨ�P';;�߳l�w�gڒ�::��=����l+T��%���I��o��ӱ�3S>

.P�@��-��`i��n%TV}���a�<���x3 ���ev~I7�`aPכ�Iw��j踹T���	�%�k��|u�,i#�O��vZս�nE�Gc�<O�w�%6�3}� G�BXXkQ��;�ĕ�O�'�X0�cx��f�G��Ƨ�$S�jL���O�\Q��QNP�efD���ٶ�"fpUR�+����k���S�n�/O�Ԛ�`d��`����X.];�ɮM�!�E��$��&�4=�	���g��;�(9��;�C�6�؛��!��οMn�^d�����y�Ɲ��pP	2V'~L�8�\<U��M�G���Z�uI� ����Q0EIXV̀�o'�\��o����=�������:;���Z
nٺ��XQ_ڰiU�w�t��ӔH�w�,��ਢf]����>���h������:�0����U�Z[-b����Ji���ءQ(:�����:v:�A "	������䐿��5HP��G��CcK,b���Pݭ��|�v_�ua;3�/>?+Z������N߇T�y�K6��x�l�����C9���t�[�ɉ��t��TFWhմL7o�Gh��h-7aPل$!���g1�`�f
 ��l�g��Q��P/i`��q!&k�vmc���<�s&�}��ޝjp�?@`��|A�n��D�J���$��w�g�.�2w=�5����B��v�����R7n�RrT|�u1�>��nQ�B$L&��)M�����l�Tt9�������P�t���;��dh�\������>�&ĥo���:��&F��cB��Z���'��`�}}����i��D���6��U��ֺ0"�&����]���V�M���-~�����u�7i �U߉���@�bG��	�8�K&�� �>V��fiHr�P�ݭ���&��[hj�a���x)���;�e� �����y�=e�P��Y���<o�**��n��l5�����'xU���䧧�Z�ea��8l!��	��Yrg�~�_w�<:��ʑ����'�|�כ�F�<FM�i��7+��fG�|I���F�tQ������D��n��)`���ם��ӪJ�����zbP��Nᨶ��%}D(��I���GU돢`��n���� Зc~��_�NH�D�$%A����
�k�[+镟����.l��j0��ӷZ �n��H��5>�9wx�+E��'���I�G�+2��&~X�}���k�s�d����$I�<��ڹ�t�����!>Mh{SS���<��!���-��0�����5��H�1{�/����0NKhY�$94kӘ/[]Y/$�\N֘�,@�}N��ኁ�pqׅK��K����������M�#3�vf�������:���N�����YQ���k�)�su�K�"%xAE�Z^I�!q,�S4��,.e���ްc*ZnV�Y*�{���� Je���<�7�y�����bZzWW<b���Z��%�0��k�Z�}I�Ϛ��ݽ��b^p����\��9���va���~�_��E|���!���T�jN5Χdi"$�(QtЦ[#�ը�$��*���nB��b��Q�� ј��"�OY�Kڠi)�f)�<�5=��C�B�6���}c��9E�a����������-�P¬gH�A�#��F��*�;c/�P�ƈ�/ d�n9��x4T�	
$ҔU��BS��0�W�YB�mZV����*A޺���ŅO����	B �zY �Q�*	�����nD�1��4����bɹ�a��,͆S�9)A��@���:$����!���o`6ږ"Q��+`�
��A�Ͷ��4s�����9�=b�$�L��B�^��?�d/��Y��o�f)@$oOK��%����<U͉y�����������="D��jַ�L����~l�Մάcg�����7J��"���V��B՜�h�G4t@1YVݨ�N��E��h��HM���kε<��{���)��N����u2;WX�k�b�UQk�-�L�����UU�73��z���N ����A�S2b���d{՚��Z��w�w��JN�s��\�kEZ����c�ZzI(��8�|�ilY��b,U(�U�B��5аB���f��gi�:Eaϧ&s�6_�k�.���k�����ĳIF1e��Bce�lxa�u�����>B�}8y݀v��bD�
!�����@���xς�q��R OT��/p?nc���@�q�3ꀢ����((:����J^&���]��ڃW��Gy�;G�4�h�eG�.j�3x�@I��(���GR���w�/������{��j_�f��� �������
�?4˔��bz#bz��^1*y(50��t�E��e�/iY4���!���0C^��v4��[�!%mdD9��>�b+���`��-��(2�zv�}�d��tk`U�'2-��ɨ����������H���s������D��e%�����N�$�z9��a!�Cv4}|o&��(9����^�_���pJ�����>C�Y�G���HB�* �(��L=b�G4���El�za��]x���5B����.�G(�Q"���&����%�
�o+㪫'.�R$��!��1�\��<ᯢY���ɓ��"�쬢����bjjC�Z�ܗ��%�}̬��a���V����u0%����i��?�@ ��6�UV���UZ¸���M�*�u��3:G�@�ڝɑ�l����I�	�� �ø=뇢fA���>x�N &�.�����Wʪ3�FJ*%Ĭ�`r����!=�`�O@�}���5=�r��%���-mxqn��ɶfw�jU)EUU�߽
� ��K+	>3�����^jp��\�)!�4PK���lmݶO�b�'/(2�oA7 ��(h���@A;#�Y��QH��h�_��*���A�������A֫��,���b�g�_���gH�i�GIh�xgx��v�kue�=$J��U�����#�HP(r�7�\@3H~���8k�I.8��C_
��ȬW⩍E�l]XL���r�^Q�XT�#6�C�gq��s��Ф���w��,�0a��_�F��	6m[0��$��p��-���W��GZ�rn�N/�6㋏���_�����ky��������xPLLp}�QN	*W�'JG.Y����I�Qn��rk��[�N�0C���OVk}=��?CUF�,��bI��#6Y�����ʑ�RI�Rzk7Yi����V��a'�2�K�����I��Q�|p��*4wK�C[[7h�NʝV�U�8��:u<7ΗD���=��}�W׈V��ʏ*�����1-�u�lc��s`�o���ܿ��Z6 _�=���
��LE�$�m�D��R��^���s�,�
y����M�-��.f�Y�B�
����&A����P���T�u�ȁ֢���'<ߛ*W�!'[���)��O���BBsz�m�#�5<���RS�qQ� �@�4	K���E@W�wҟ��F������甆��q�J��pp�?�4�����х�Z�a���|����Z5�[�`_�,4��Rʊ!!h�$��Я1���I\��1���l+�ܡ���p��g�&�o.re��l22H�[:P�s>/^�Ό�����V����ݮ
�<C�z�' Ϙn'��*��8�/-�Yk�\�}DqqP�AO	�Yn�nTA�*��K�^N��qe�U��E��7���m��%���s5x����g�}R6�������IA�2V7��_�FFPX���Wu�_�xㅱT6�ڈI{:�SrG��/�]�lW�km�V�:�A��P1�>w��ZB��	)7�:Gz�CpK�+B+X�$�7��&R���<�֋m��&r
^8t�I~��[¹���f����-*�Y��_ ���0RK��#�J_�+x���h�a~��u��3�`̏	/B� �a�v���3�pp�UqؕO��e��A�\p;)B��ٮi'%�8_�rI>!M6B��䖓U9\W2�G"8��w�:7������9��zbj߳ɣ�sY��0N�ǩY�:�
�O5����t��X�=(�o�:�5�N��x3��*e���$5V��Y�T9��"�����#��i|z8^o'k��xz�����n���rډ���q�zPD�oP�l����L������İknN���K��5�ꦡ[؀`�#:b��.&��h�>�J���k~�՝E}�T%�C�?s���'�!����H�搑'kj�7��������P��}�C�3��f�tyH5�Hqd����l\/�Y����=!�1�%�$���w�̀���]�B���u�������Ol�t;�9"�^����?��P�^kXİ�I�8���'t���-�-��U޸}d ��d�usA�Rv�Z�3�t�Eã���.���v'��Qpe�99
彊o@ �hr]�MI�&OV"dC)��ŃbB��s�v�m�ⴝ{*�K��zb�^)�V�����2�A/��(>>��������#�����k0L�!�Ф�B7'S�H�W2��;��,C�}�#�@O��A�(�j_eP1!�4�s�h1�� }�����]�X)�3d@L�p~g��lx-P8d��y��z�:m���T��Pշ����i��l�R�=X�*64<f1��y酩˪��5P��k^�@��8xII?�~�T+�t�>�A'�Ҩ��f�F�He��d���ү
L��Ʃ�5[.��Ku���U_�iO�~T��mרz�	�,������
��ܹӬo@�iJ��o&	�pfw�@��U���l�T"��c���be]�k��KCWN󉱨H�ެ&�۰�L'):z0&/�+����r#q�(�A֯Y�T߳&F1q����Z�T�9��e��;���DY��J�[���O"�;Y�K���f49�q�&$��t)ATl8QSRc�Ǵ��X���b�#L�a'�&a㵖2܌�%��	��12I�q��m��c�_%3�;7�P��U��uw~�a������Ƨe�����;�O�����2�H����4��VW*9u}s#TW�N��伍��F%������TQQe�V��_5��/���M\��{G�K?�OZ^��qW=��A�F���V�����<UV���M��V��7MVZ]���bn`�F$J^�����-УV���K�w$B)f��ǁv�d�9JU��Ro�g��劸H�]\�����5rTP��x�������IB*zV�~�}ߪ��ȀF^D�o���J^y�x��	�Cb�۹C$���'L��Pnj�Y�k-���ܭ���0��sG
nj۹:�Y��HB�;�N�f����_�������j#��}��g~<Ӥ���꼃�C*vv���)�P��*��kw/Ff�l�f�9{��yoդo���9��ȓ<���d�9PH�������[:gp[׏�:}�Q�t��Q�
���V�)gP����^l���ɺ�r���8�!��?6�+�f�R���M FIϊ���S=�����]o�׮��NFQUFN]�O��3��O҂� ��9{���ܗ��#��N��_����ԕ5�UU>Y�R��OV�U"&U%d�'%����լ:Z�{ܛQZE7Ng�?�^q�Dko���#���OU�����cG�a�w���I�>�J	���Q��Č�����k1��F��V֋�L���_������o%��jL|��'����w�j�u��%"�=�̏=��Z!i���LQ�IYsk��;p!:������%u������ڸ�deӴg���Q>⊾�?hֹ�ۢ�[(ΏքU	����^4
�%�E���X�/j8^��"y��<�>@a�h�޻����9<K=+&���H����i��^�3U��%�|K0*�t��՝.��|'9�Wi	y.c�W����F�\�H{�*ص���aϳ��6E�*��ST72�,8
+[al2��j��Z��6\D��l��<������}ԥ��(�q���B�ίG�ǅm����[������7�c+4�*Z�m�Y�Y��=A����u���q�b��� O����\y��<��\0���^s����U6�<%�
ծn�ѷ�m�y��H͈h�ަ��b+쪕������A96�ps�/*�5(�o{���f�4)ag����o�2�`��n��*��`K_�ő�}�(6�2�Y��m�̓�����.�Oa.0��/5,D/��#\�Z�^�VUx�fw�{����xt�W���?�hV�<VoY�Ԋ��u��^���;UJ��%\1�����\-?OM}��W���*�9�:�SPL4_��ef���a�E���G0x�S�ʲ��+j�ۗ����wQ���ڇ���Ƀ���zh,uY�&��C��?�p�x�0��~Mu�����N�Ш^x�
���׮>~g��U�����N�u+/����B=\Z�( ���m^j���7AZt+l��D<0�X��B+�Z�\�*�������U�V?V�)�.6,��$^?E�iF�5�k��.�)*~8®ҷ���C/kfl�E�e'�,Ƹ;*r���u�lى�߄Jޤ�t���r�?�0M�W�������� {�qV�'�$���$R�<�c�;
�#=/�ݎ����� ͵<Ά~���Mz�P�2S����1X��Ē��)��W�iW�TŔ�_����@�2h3��� ��Ơ�e3�P
�W�	df#d'!!�֟�2Zb����m�_6y5��/\R
�鐞'�掩�<������Y$���v��Z�ɣMl�M�Uv<O��/�l���{����ĐO�*�	�F�Ȟ8ב��׻�)J�6@�S8�V���6#U/��ߙ/�}l�("�'��Td�uw��>���ֈ�8���6�4�ij���A�=^��7����?_��,:�G���~�p�4�햊�MO3l_��_�=?5L�M��i���:=D���i�����Ce��mˣ�]@������6Cص��jQrb�t���� zl��ܮ��`�����N���]"%��m��o���7+|ww�A�Oڍ����������l	����ދ��t�́X2ݟ���v�����1�HVF5��}�h�IV�
Z+�ْ�)2�y��3Et�}5&���ug6hI^��le�w^���Ż���ɬ�C�4q����LH��	x�j^Ș l)㆖в-=�>>����ј�X�v���0~t����]�S;�}H��Lu�"e�25��������z�a�K/�a{���2~�b⭳'ݵk'�Y/�Ζ#��iW�~���XY�Ol�_n������VEr�u�4�φ�})��Y���#����?���'2?2��ה�..&�g�.�}�'M!��JJ�挈�n���Z����
ɜ��<��EIc���6xH�T����O5G��.&�qde�wU�����t&��*5ORy�vǸ��|�hG��#��&ufp	����P0��v3�����@�ҭK7lg'�S�x��]8zj(��լ�.�Ji�:\�3|�c8k����:w�YP �F?�������0�̳ޗǛz������Ԑ��{�K�1|T���g�N�uV�4�:��o֗#O���,�)�)Tl,�ɺ^78�#�л�
ac*h����ԗ���������W���	%��-��ާHt�K���8MkFz9�O��tc5��E�|�~��$�n}%�_݅���r�Y?L�h�3Cp%��X/����*.hg�����6�sJ�	ˠ)��E�S(55R}3}�)ܗ��ݒ�޼�g�Wpۿ���
�i�>S���d��0<�D��D;_I���!Wm����b�=b6[�|�?��E�w�ob��[]���k^(ao[N}��އ�쇂��]�Q�������ح�ZT�������nQ���Y���]8�*���|F%!r�]ZA(����..יx���s��?LN�Y:/�q�<����0�G���pI��
G�K�=I��z(&0�<�r��|�K�5�#��݋A2�ۖϦ�{�FN���nUe+PkY"��1n�E��Yv��A�m��v�S����tJ]��g���x���O8gu�����g��z�i,��n@�H�uu���d"^?˓��L�>H{đ2�Fљ0H�b�?�+鲧e�^����6�>�ʁ���5�C��Q�O������%�(C�Qwn;v�s{w;�������;�L���4/��<> >��շ�vV|W�/�����uVI>=�.��ݠi������&�����_�}ܳ���xּv=���y�P�3�)�_�utl���9����}r�����
\q?7�?
�d�=��"MX�2����7��k#�����W������G}��	i/T�*t���F��`%��1Ϳ�D�Ae2��o/�aL����]��4BH���M�;�*ڠ7:��h}����7��ǜ1⥮��$V}>_�Z�rV{�����;Q���U�ϛ�ovkoL;p�cc��u�����ɴ�tnq��g�@�f��iN��{���&䁡H���\\|�	N������w;�L(����zԶ�3�߅|�=Z��6���[���L��v�U�k:�9��ddvf�K	��/	R�"�y5��gN��*
���|��t�L��|t�y}'j��5�jv��M
�[#b ��>�<g8��h8w���]ڪδ�_>�HJ�P�ɒ'�q����j86��2��B�����zw����A�i�䰬!Ę�C�gK�k^�醴��~�Je�O���^��$�����M�G�X@�{��i�}Ӊ�q���77�w�wsr�����'�:u������Ȧ�j�j�ֿ�~y��ׄ�5Ѩ��@�a�#`ޥ�?�[zF8��A¤[>���V^��d��2�\O���}���|Q���#�3�u?H�ml8�c��H7R��E]�$�ْ�͖�c1X��oƚsm�2��J;���_�H�U������u���4Gm�3{_�m]p�¸��h�]키=���9��f�7��!!��.��N7�ޢs��H�5��� �Z3�6c�f)T������w,�ұ���Q�p�f��Ç��k ��pw��#�=̲�'�C�&%I��
W�] �m0����������0������׮Uv5��PZ,�9�;f_�V��Ҋ��"��ٱ�*�i��t*U�C��&�Z9\���:�1)%"���2fM���K����ӝ��0���(�z����Kh(��y[X�zJ���8i#8~�J	��dG�&�[jaV�����sN��u+�0L\xx
G��#�R��ۅ_���������pE�g����Ƴ�j|C��?��L'IIǌw��Q����T�v����fL�<"٪ρ���1�R)�Uf�k�i_���s-����녖KN�~��@�3v�����4y�w�ηa��w�x��^kX'=�(<>�k��
ЕFi�|�[������b�܆��~'�NQp�m\�ۛ��������	���#�E!��Hg����qа3�G�� ��3��	��)K.����dO��?����>�]E�^m}F���,z
�h0Û���i��r��RE���a���ڿO��:�1�Y��C���kLbb��O�AQ��"��q-���﯇�B�������5*�|�,rh��2�$מ7�,
�TL�.�#�T?ݧ2�K"WT�ɥ���E��~���9IvQ�sm0���"`�Jd�D��a؛j�M�%��
>�;�<�����W����t�������<��L��D�N����$r피�����"��|π��U����>�#1�D�~i��� ��64j��@y��<P�6$y�gDFD�cd�}�A�D�q 34�b�͆ �����5�,��kl�΅6oy��{x��ޟ�,3�~@Ŕ�WTi�&�.[�I�I������p���-ݜ���Yo��_3d���m�����a���=���Ԯ-��khd@\�`�9�?X�9�ݏs83�-��*g�|���5����NO���>��ǓA�Zfݭ����J�T5IZ������h����.`�����Q���ӯCy�3�aHv��TJ{���Ŋ�g���$�	C$�eΧb�`�,kF0x�Φ����/cȋ��^���v�dM��\(��{�JE=�'��ML�w���q𙧋��v��<�rU�`�0]��&5�k&�-hh�#a�1�R�=���ľN��#��1�4IRp=>�Щ��da�AGA���FAh��v%?R�=��(W���/��t]�6�QA�W�$%x���x�v�w-��U��y�α9mh"��tHܛao�y���rBFF�g47�a��Ί���FtDE�2rP*��OZB�b�hQ�S�q$����ř\�m/��L��ڣ(eҸiʜ����.�<c#(X����/���dM�?(�ۭ���m��,�y�D�C���)%�#G]�А�����f,��y�;21�)��o�յ����M�X�|*+ �V�ޘ��e�T"��6��>ж�D������mf?3������g6�8�>���`X��|N0�%��p���A�M���v0;�]&�����5ʴ��*�vh�~U�Xs� )�E�;y���2�y��<��03?��-U�l �V%I��M�т� l�����(�1ޭ>�q2�iup�!�چ��տo����
���������s�� ��/5q�O'��4J������{,+Mc�����.�� b��e�ӭ���v��U�~"|޽fN�S�=7LD�p�x��bU�牖wխù��ܹc�Nާ���V �FO�C�y�_�߹,̝��~ް��|��x72u��gS1:I�2���U�ɾ��V�'�a\�E8)Y�pa�� ��/[EH�{ŝoW�#��A@��!���}��\�?�,bsv�'E��;5Y'���AjMB��ٱ��}���ڀ��(�&I=g�Y���00�
EL-٨j���� k�gu��W'�ZF���es$����1���񶈙(�J�9s�|F�9����T�8］1ö��3H�<[(�/\�u�+3O��7�����N["4[?d�iG�tY��9�u�eHR}�<��ANj���kx�0��߮�A��Z,
r��]U�?�Ҍn�ྵU�y3�'��!�
7����<���k	��yӶr�^���,pf[5�ɾMwCM;ؗ�'����r�DG�4�,��FTa[j�w��C[$�~�}����Bh�Z��xZ�B�{7�����!A��ے
0�8a��	�wk�ZwY�pt����\�'�q���jc����^�l��q�=LI�r6&�l��U��m���}s/2D������#�x����_�J��)��eB���Pd$z������LA�``�<��dm�.W�eg��Lo�BË�!b֩�e��e������`�t��dV�a#O���7�����^1ۭD�wf�⩬�M�l���9�s�ejJ��/~���-����v!ܶ���g G�.Wh�T����1��Nd5�4 ��C&8�$����<�?��~��c����튠��q��z�A�?7o�~X������y�S��5^��5j94?���!A��H�x�y��9w��4ߏ|�8�m�Y��k�`���C�{�@�9Z�V���ND)��Utث�4�"���A���KurcW��"�ǎ���!�����A��wϨ&��mto�(
J�ҕ* �H��k Q)�$�((E�7�i��$"�{�B3���y���9������^k�9�ٮ����ccS,�=2� ��Q��%��6��4z�	�Y�/�@a�:��&Fe�����˦���IV�I�m�	X����:c�*N=��}�\fR�SU��s���������N�B�HӀ�������^�ݥ`YO)W�J��Jƕ��P�ck�i�싼���k�˷ێ��B�S��8(��+Y+[\t"**����i)xkjKߔc��NIIXb�y�����_�y�w��3.t���ߋ$�z��$3��]��߀^M�!p�ѨP�lw�I$�b�\�hea���2��y"0UUqO�2�������ģN��m��l�z�\��#~������ȭ�9�"��C��!��~���b��7�#���������?R�彜�n��BI��<[m��D�t�ew�橬55�++�����[�u�r�ydG_�%�Flp�F�oae�a��cv ��Y���A��	^�6p�*U��(��hr�� ED�;0��v�"t�bu�٤.�P�<K�p��Ի�yjV�?oy�AZ�
��7��Q�x��|���a������R��ya:!��/��P0֒�k���8�Z��}�!ٻ�
��ίn��PT��!�!�Β��d��#-��op���y�,�yb"�}�Z��Y�K��8z�tW�ɖ��_�bS���@v>�-���~�;A����q�w2	'zRK�����侟 �j����V�q8�]�-���<fK9N��ۯi|���X^(ht>ġ�	�YMs>�����qW�,r���X�t�������@f&cS4�	5�w����yz�Lq�9%�-����D۬�`�jբ/x�_n�&?���MaD'��=��0�88E�d��F�=j�l���u��V�Hw���¯{B�pd��	��C��֜Q���<����6u�^C���ϥ�_d�S^�[���_H9߬��/y�j��YX侩�5�����Rb�|�FoݙF{ =�]�������WS���j6G-Y�%���-0�߀٣ʸ��NE��^^�:{�g){����'�1[���xr�,_g�`�@���qII����O�h�CŭM�)�F|���+���XWdՆPw��ǎ��8�Y1�d,}��ֽ��Ȭ"���'�2[ʧ��ʟ������ݵ���Cנr,g�_�- ����93ߓ�I�t����=��t��������_~'��/h}jc����%t�c--ޗ߹�U�i�(aJ��@�3��>T:P|*���)6�#4�?̏Y{��qE�f�-�ԉt����ͱ���jгr��?]&�@�|�u`����-.��)��M���� D�o�#+T|��N�J�T�i�'��3����?�I�Jw���TDn����g���
XU���:8
F��/��B�߅N�B��R��j���$^���4rB2g.�w(8V� 2��{�q���X��s>/��6+ujm��AW����f�A�Q�����G˩��Gy[�5�-�f^��ӵ"2[^BA��OvFi�S�E�����x�Ȁpaoy0t����y`f\3m�{W�2B��+��]�,�0h;����xf1 �d(=���3>�i�zwv�)�2������Շ@*�������}@�$2��w:�Vj�.`C	=gF5�i��քՔ�;�{�`%��gr5�"��(�YQ3�E_�x�!}����%��J��(�sAۇ8b��Ե;��x��ߍN/������]�c*+;����	�����4J_B���eԲ�9��yC]C_C�'k�V��E< 4&?zJ�Hj����%�ן�2�i�B��eV�?܇���Z��Ǿ[�5���]�+�6P�Tc�����ē[�v8y<�U���!�w�Z܊��6�V����O���ڀ�НL�D��ѭ�����1�M��	��y�����A�<_����zw����j\ܪ���*��Օu;��}�"�v�d�*��Z��_;�/��*?��j&|��F��>�9���Fag���?��Vm;)a�U�pR-&��<�\y�cX;}ɕ�h+�\Ex����B3���:%R��tGc){�����\��I���I-H���&�5E�6�$,�
�;��ͶS���Z^I�����I/�O����Zj;}g����M�Ζ>g��r������%��쪚�贴�HB��Y��;�ҹ���V����:i��GS��k��<����L������Z�J�5tsr�Pj��>H��k8>�O�]�`%?$�ZLjO�J�'��RP|x��
��wt:����쟈�vR�Q9�;N�<�lf%�<�-~���]���N��Tq@�b/�aa=1��'����@(�K�t2�L�6O�X����1��P"�2��M�{R��*"m���� ��ʏRS��_�~lW����OÝ�L��_�RT�{}6�8*���maΏu?�/�a�?-d�Qx�Ls�aWVQ	�rȬ~ɣ8�1g��mn�������n�������愦㏔�O]?Vܜ|�8JfT�n2�6|��_���)%��Q�QA�d�Lt|����	[�Y#}��+aB����2������u,%���G��S��SmÁ���)�P���8���)*��+?��vp�C�Q� ��c�@��ޠ}�(%��s���_жO]�Vpt�޷¡o8�ꌨ�HY��,4�u�0ߖs:�Sf��󯵀� �ƓoT��ƺ�?���t��{�f����ǚ�X�c�CO5W_fi��R���y��]`c�G��K�ѐ�nɞiű�)���*L����SSy�k���߃��Y���������"�� �]��cVa��=�"R�������)D���,�����u��i��  v�=h������k,o�ս�=�D�TL�QD����k����}�c��uXV[��>R_hŦ����_%���
��\dQ�q2Mp�����7���_F�O�C�g�E���]�H�v}V��;�l����{�^2���=9��[��i�g��J������lA���+��W�^`6n��^ �����N�Uu���-��Χ/�=z,;�����ﵐ��ź#�Y�8"��G�=KEO���?��A(�;��_��h�KG��8����ܛ�^�tO4�n2���z»K��2UjoЙUhZ�z%V��e��F�3~��#��o�jU��9�P���9F����3��=g%�҂M�[U$\Ǌ��=�����&k��B�!2g/�'d &��5Pf�h|g!��w�6i5��u�l�������+�))�o��O�x�([�d�ʺM��#z k~<T�f�����J���p~1ot�5��vp�I���?�;�?��<n@,�m#=2�RB�����3~���Ǒ�$v�����E�IK}�G_F�Ά��7/�<E���lf�����d�G��!F�s��$�iw�]���������L.\����z�Y)��k�p0q��,v���wn�c��`���XY/�N ��՛o�Ĭ�''�P*73����B�As1v#�es�,��k�T4Kؾ�����7�)`T���ǚ�$�(��t�xx3 �[�9�B�ϊ_�Ւ�y��s�����H���}�������a��2���FN�.<�`Ɲ=���	�g۷'���k"�>\�z�S;��?Λ�8ң��� C�8c��}آ
���+����*����^�*���J�a�3�)�w����{���[����5���Lh**|�N�e��M��Tђ�YM6�q�J��z�B4$�nBc�u�w6�M�C.d��z���K�"�cP8=<��y��X�5e��s���������m���������}��-
ک���L�Y0Y�&�c�-1���?x�}��#a,�|u%�m��e�<茟ͳM��u�C.�2u���ixkC�Ͽ�p��5l�w�U*��-�����k�բX?�}�x��O���%�:{8.0���P{wB���9!���$��w�5���Iر�����~'#S��y���Gc`]����� ���|��jŎ��$L?
�������(1=,?:�q���䴍�b��������{�<�_�Y�F��=l��W�y{)I@�����!=7��r�X�8^���?F�-�g�vn�_���nzvXO}��?��B �lG�S%%Q�1ozk�Y�ׂ4^	B��Z��3��P#�l����Y�L>�U�)�����?���;0
� *2�Fg__ U\ޮ}�����������EJ!΁�R`a��Ӓ������y���t���LXh}�}n�g�`�?�����-N�_[��r�T��II�2?{�h�@�k�k{��$��*_L��0hi���N�a1�F�hvH�?�3�ѯᖝ�����o~�zh�%���[p]I&��=/�3���ʡK��&qq=jl��)���)�*ζ��'��OL����3���lz���F��/�h}uJ����b�!�����Ɔ���w�y�Te�uB��~���a�o/C��Ц��Wn�p9�ɹZ�y.��H�Fd+�����h��y�.	���%v�����e��#�іMw�c�O����H���PUA78��@7U;��l�e���N0��������÷����{<1�&��y�� �M|�<�v�-
�z0�y�Um�� ��xw�����ė����u��e~�]���ɀ}��skQx���S4����_	���EU��4h`��,�k�0z�s�ҍ|���=+�}Ǯ��]����i�kc9B�s������ՠB� � �61"�v�\iT�I�-l_)3ߞb�!e���o��&��%>�(#�����ܫ�2TT����Q��x�E!)����^�On
�=$�0��M}3G�|�[�F��.��_P���{��w�i�s�B��l;�z-�8y4�?���-�P
���b�}5(�d�*n��=��7���t �N��������*Yx�����~��u�46��s ж��!�	�r�4�6m߿giu?�f7�	�!D�"g����ࢣ�=j�G���iGa�ΰ�h;T�Ni5F$��ɓ��j_��Q+]��1��f��PrKT�U�4}?�9z,/O%6��Q�g�7�:����][҉8��LKS�����&�hd˃�}}�����Ne�5)5�/|"xB�M1�T� l絤��L��������O}~�[-/7w�c%�WJYM��&(A�JuM���L�a5�6'W,]��H/��DX9�����F�x��������T�]�Ṗ�b��������,���}"7&�*�@&�	�4�k3��5J'���e�c���4���d�3�Ri��{���^�!�!!���4ϋ��Nv~� mc ��O�߶�O�EaS(ګC��Sl\��<x���>�d�u:���������B "K�����&�4:<ǳcsIO�Y,��.ͽ��A+�G�X�h� �To�\p�0:�=#ׄdLɖnb"��so�ud
�<U_K=
ҵ�%��~he�v�k%���r����uG'� d$���{]ZIl��/��duQ!Hc��k=Sn6u<������hV{��ek�V҇�;5뎀��KBx�b��o��1!�$>k��AZy@X�W��x�1�:EM����7@fq�[�*���}����d,�~��m�j��ez�e��g���{ތ�È��|��,�5�����׶���s0�0(�0 ��j�Z��;�3�λ:t���B/1�PH�2����;�{=�C&Z=�
����5"h���
�*���자��5�Ӱ�&BK��+��޶�%������W���<��H��'5m�Qri���� �����c"j��~��7ݕ��B�J/.w�}7�J��[�pڮ�D& 1�[~��v�tj�ٽ��H���`�:I�z
�y<����FG�_Gz׺&#/}��X�C�y ����s�V�P)�(�?9����%t���V�nDf�+�:�O�I�A���{y8_d�p��R����w�<����8W�	K�J��<0�hv	BG��]�;�P1�]Zw��-�X���q�IJ[.��~��Eڃ=ը��^is�l�=�^qpN��;d�F���usf��:D[ݗƽSRR������Akw��y�>�J�q0\P�>\�'xo�":AA���I�0�T~/����9wˡI}H�����@�w�-
4=�E��k�Ǵ3^�sr�����H�a�	A��1���^�%���χMe����\�͆�  \,7!X)!K���˂��L�C�-�&RR ���g�9<�Oo��fa<ʩǸ�Ϙ�%^�`o�|'c�ly���V+0�`}�t�+�`���tx5� K;�@� �
��q�-�V�y��儒[݌_������/C+�J<�}+.@��7�Lb�L.pL\w>�+V�FK�o8�5T�$�G�h���z~t�Z�^J�;����e��.yS�����W�M.���?O��8�O*Mc8�]DT|*Y��͚����}�`�
mmj�<{=b��QA���UI�o�nd.�3�M�^�����4c� bk1���-�q\R���q;��N-O�J8d�ğ�e�~�����;��ቀ��/����X���诈�kv&M�����\pZ���V]s�ŗ�����Q0BÔ5���kD�C�213gƧH��_��&�'i��x���\��/����7L��8|��j��5�A��
n9��a�X�ʿ����AE���f~�)���v{�5��[b���{Q$��x�T�5@<7�HG�ځ� 9�|�s�?h���s9�ϕ�<��k�y'�P���-��V��-���-~� �{��ܗP���x!�yS�	�@�[��X�m�c�uM$Z!x�i`�oZ�IY��U���Řv�O?2̤�t="��H���(�;�<�g�G�'<2ΪE���IPO������h:�N�ͮ>��Q����3�<��Qgr�a ������z����9�͙�vmXX,:���#*�.Qc9�~)�<-fx����� y�ϯV��nJ�m�NPk��nڑ&��G��b�E4�pa`G9'$��ǻ�d��Ϭ�D�08y�?2p�c�B�`����0��/�H8ko�"���U�����IЃ@$�M������ojOad��\����b8,��2����P���x��)!���#㵸ر�Q�X(��&�~'�rFΘYX�i�]����H�G)�r�'�������y�{��?F��|���#�9���i���N&��`�����8K�qT��E�hr��[�?Q.��!��Ȅ���R��VF��5�&��ja>��6���(��M�_ae�M��kU���?�rr��=]�Iُ�� ͘�A�yaO�}�Jz4/�*���b����I����=��ъ]�s�?�9FV$2�姍�lM���������O5DçOo�w��D+�Y�^*
O �s\�Cc�����E৾�$yS*����=+���@�R;s�o�c��+���SS-�h�<�(;�J��7X��ۤ,.{�e]*�k	�e=�$���Դ�"�_��ܫ��2y0m����|
~9�ޚZ�80��<�e�iq?���UY�f��8�oj�˰'�����-.W2n%�zeք] ���X_;�C{����7e���)��Ȁ�G5\��q������Q���k[�廜'O��_�	����jgCQe�q2�D@����ۭ+!kP
YN���d�ئ�}=�$��ؽrީ���n����?��Trc/������]F���ȴ!cw�lϭЏM�璳��4X�P��_e[�Ui�c�ql-�"Z���omw��������
�H�?F�xxI���P�U)��4C(���޲ys~����5�$ES�{`���"s��0+j��@�<!�'#p#��y_$��m��2���|o�~���ᙨ[�{3����q�ݥ��E�H��3����E����y'�i���y���WeЏ&�EeXm�
�~ӾS�I}Wy��`�I� �3���Y��[�O%g�0o�p�;��w�[Q��u����Q�xV�]���N�R|V�?3z�NVИIʜ�u�0���}�٩f0���	��hH�י���d��;��]���8��a�����ba-E ���\�?��m��������ȝSWo[�
��V�R1���<!��Pm��$kMPy�=q����	�|%?��5ғ''X�
[�5VX2�A��kk㼝��"�����q�$��^��@E��~�-m�ĥ�F͈����)C�Tq��Ü
:���g�&���!}]�,}�K�^{�`�9%{o�J~���Q�ˢN��+((2ؐk�q�;��u���_Z/zv�<��W��������'+{��1J���mw<��PaQ��>�%�� 0�4���F���Fv�ap7�.�f�JQ Z/�!�(�`=՜s�/,撲b��feH-3y���}�ɾ�5Ğ���(������=��
��d�"&'����6`U}r�Vy;g����PvƕM��oX&g��<�
ɷ����|u�\����	Ԫ��N����h�v�(�!�%J�q�94m���f��� �-My?$�/_\grd�vڇm	.��t; �4-7��4f�a֮�YIkR)0�D�|ҹΛ6^~�?�5����u���i�{QQ�:}2OFJ�fPG�[S�7��y�3��K��4�������K��)�]�چ�x���kKzG�K9LآP	�W_�ص����-,��K�w�&Z��u�*0�#��&��<é�Ap�D�>�*��O�%絓��d��|�RS�����u���̌��T�3�mS�������Y��T�0b�7�v��O�:�ޒ�E���/�qw���)��PE�:�ae�/W_@�q��+ف��b�&�?���`S�`mM��?����D�|���WѪl#5x�Y2�����ݿ�����/�����8��]uIO]߿q��˱��˺(E�\����q���-�\����O	&N;7H>�Z)�F��e��u�� M�i�]g�v1��H��z\��5:�U�����g�a�a;x8o�Ʒ�F�z�/O�(/�p*�[�ㄼd�}$Y��O�#�-�:�8*�/������k��i՚��)4n�y�����fГ���$Y��jl_}���Km�q���W�=��BA�����W|:�N�?,��Y�o
�V��V8Ђ�W�VT���a�c�+�_�I�.T�=�`(.Jl�#�/3�\/a���k]	��9- '��{�7 �pNaZ*s��_�E�&
#xyf|ZV�
^٬贚�4�4�u=G��ޡ�m�y���!lu�NX�4L/�b�N�˿-פ�ޛ�G���ܲf4j�uc��8^��)����9��>̧���`n~gVJ�W,8KN*��3!�� ��\Dlq��Nf�<;�kY)	_.�][�W{RO7�=A�j�'�qW��lu��eChՈij����'\>}��#��F�G����Q�SW����:4� �=	�a����g^�跾�қ�M'ĳ0�í��#���5������5�:�-Jo���{�EKi�J1(�S5��x��i�K����{�����S+M�6�]6L�ivky� [2҇�8�)�^^x�s<@�0�5��4�~mQh���k �{��}2�IZ4to'�`(RL�f�OW?m��T��9���Ir2c��T�������@vӯ?0WE]=����&S�yJԲ� ׿�����DY�»�2���:��uT�#���2��Jd��t�k��[=�K[���٤����W�P�%
!�:H=�e��v(�\��3H�,`G9�Y�v��X��1�y2����ӊ�w++�f�#��%�ޗ������Ё�̾Ul�
�c�6R�`����R�]U�Ш㸿[�$��H��5|ʌ�8�v
���*E�B��Ë�AcC�ή�Y%�B����\E�-]k�p�ŋ�Lb@�;��_z;;Vl����v��Oч�a]�����ݓ"�����P�h���l�;r��y\�Yû��V�7���v
S�ɽG�'�J,w�~�sј|m��}'�f�Y�vsm¤�`���m�'Y�gi�j(!F�|噏Әp.�Ojk$b�lU�=�r��u^k�E�M��Ξ��{�AaMݧ�����^�[3o��H۔.�������	||���Q�
�!g�"���Oב��&��U����s���-j�Lx7��_�ˈ�8w��Њh�g='�>4����q]�O��0r2����'Z@��#U��T���ӡBZ44:_�@�V�j�ܝQ#��-�g�Ⱦk���$qvC�dj�D(Ñ�Wa�-�MtH�uz
�uu��5��Z�HŖ��s�SmQ�~z>3Sc;�O��$�w57����`[T�#�	^�LoEyK�nߤw�:�bl|!̺�zdh(ϣ7��CG����k[��&LZ��,��u����߮L�y6�Ⱥ�����G>��O���K���l@����i_� �_;p��R`uj�Cq�����,���>��q(|õ��H�PK���O��ˆ|8\1�ܢ�t�sg.1c���:))�z�}���)�zԄ�����>�3<�-����]E�-��Lݷ�X.X��~4F�)	{���n�N�m2y��u�������\���~�����^����^�BT��Y(a�A��]B�(�#�C{�ș	������쭻o(jn�r�jE?&�Ř���1g7nY5:-��k�"� ezS�~+��
1��z\�E��Tݛ�qo�?���oPK����@fY�ǂ7X^��q��<��^���o�x:1r��Ꙇ��y�S��	�L��`����2q�I��� B�M&�<�����j�9�?�
��'g�{�(n#b�ױR� �?�R�ԓ�R�1�k5Gb��{���-�CZ~�����d�-���;�y���t���e�c��an���� 3IA�%6�:��}�g{K�H^2�	�Ͱ�yA�-�"�1<5Xdl�C���:+C��ؚp�:QFf���O�Z].���)q#$��L���9�W�w�K�Ͷ���ܞ>�K�ݭ��&Z���X& �[l����j��Y�ED�3c��--s�Nv�7ak����np� �Ce��y�w�Ma-��桮��/|�y�4�Ĺ��&.�m`�<��"~�f_����D{��˽������X�P��o�Vk��$薳��
T\��>*����YW��Fx�����Z�=�ɮW4h��U��D��UU�RfX�+z5�}B>�b���t(bfa΀�O	�Q%Ӌ��QD�,Ƿ\�C�uѤ'b3᭹R�3�Bp���$d�����;�Py��Z#=ւ��7	�XL�M��/�eO����^�x0#C����KiUp扊��<O��Ծ>#��N�?��~��*�J��C��<P突���Sb�>:�K�2ŮɸU�f��+%���X���M�g�Ըs�ԭL]���z��b�ReT.�l�)�B��K�^�c]���1���|8�h:	���.7E(� ���h��k�4{�v62w����o+w�����]�};�h��'jO>^jQF,�Tnd��ԛ�k4.f,��N�9���v�{k��R��l����qΒ������s^��vJ�X��.���Rϑ�����J�	�ح��`���qF��A�rO�L���K�v��.����>���dK/�g�����6�9�Ν���Z=��>zD��7y, %�( [-��p IA�J7�S��^�T;�M�%Z
VV?!Fzc.�������"�#�r�����SC'$&�8v����@�"�kM2�g����K� ��i�K�-�S�;p}�{T�TCG|���#<�|�9�5�X��8]'�Z���LyC\��D`�L�Dsa#���&��D�P�ޡ6����Y�Ov5s��X=��	���>ė���.:*(����hڞ��.P7i�\TOCs^�{ߒLߙ�
A")e���;�4��"�R�'��ͫ6�*���+�!RcM�/����G��Հ��]GK9��c&�d_Z�~�)�M$����W��kh���������Y��@��Y�Х�d#d �̶FH������ɋ�u�ݶ��Cy��Ek7V�L��9Ǵ�,�����s��6�Bk!�����/�LFN�>:np�h�3�4�n���;�|�o��d�$�
	�3�a�Wܪ*�����
U%� ~Һw|�=��`��P�O�??z���l9���1?̦�+V\|˪D�'��`a儁w�$sw��ʥ��&⏑Q��=Q��f=�*t���#��w9_6���'�4f�܆]}g$��3�>���j%'
���'�>�i���v���T)�!�d±["�}};�^���7��r���VV%���o�y%�c�T�+zRX�B�� Ua��{��_JX7�j�����L�.�s�Iq�=��sE��y]]xiQTXkԨ3Q-P�'�7s^˲�,��k"3���w�rg�F�B��6��S��n\&���	ȥ��9��"���2߀�d� f^�����7�O֏���&C[��;vm-a�ٲ�Z� n{����*�4!�UT�X��6�׹Go-���J�O>��"�`踶/\�N�S�<��=̗�N�"k�y�U��W�m�

�'�c����|�����߳��,��
��u���c��!e�JB���� ��
�$�#���9I��ǎd�=��,~!��d�M�}+J�o�u��x�߼�/#�������B�@��7��\�/�%d��+=�~�O,N��A��,�5�ϾtnGZ�"|u,���

5 ����RbiWK�<����9�LL��[�s+3��ĺ{d��h������Kr�@�Z%$��	c#1U� ����ڛ����H�.64G	Հ��%恡8Tjr����_�L��K�D��``�Un(0}��u��&K'�(��O��zl�z�ZW�,,��Q�+M��@�s��F8�l�����bgac#�]���ﻮ0�p
���-�r~�l��S�d�<�
)~=g�@����ڹ�^�ǺI�΍,�� �a��R&�=f�h'�6B��G%���9��W�Tʺ}.����ʩ8��WJ��Ui?c���R����k������:zބ��6������+[�x���	����f��o+ٺ�!� ���)�X�ZfU�s��(L^�S_ÿL|���ߤ���y����Y�3 I��.��c.7�Y����X)sx�=�[�W�\#���*e��[G�WF�ѻJ�{4*%����Կ���@�I8�Ak�a���z���w9���>zN!����J��,�h�*��ȸ��0\��_�ap%��9���.�.]���L��4|ۯ���܌>	G�J��ܚhA��w�Hes��r;���2l嵉8.�˖���R`�ڟ[#�?Ak��p`��x�Jv@�򽰳�}/�X�/�,UK���^�gb��B4I}�9�����@<����9���1֜��vu���m�p*3�V쑛��p�~%��or�e��Ii������?�����RJF�Z^/���*Vj���b;�6{��{�����W&�2�6���m�����/#�M���jo�n�ըr(�o��Z�vM����GUs9������**W�~
+��6�a*e�+��>_���2�}2v�����нﲩ;�	�+�������m��c���I�~_��=�^�82���}	�W�-%7>pӷ��]Z!�q�7�����cY��[�o�k����<<r2��'`���>��,���zf>[�A1�8�7��p�/���5V�M��3/�Ꭾ|�6�ӻ�=�
��$�
0E:c�U^���Z��ҙtt�TZ��L\_���,)H�*A��y�tw�?���qc����'*HF�L��7��l��z������.�>~�ssWV���>���<];f��z��n �	��J2��&��Jȗ�sX��V�a`O�V ��W���d��[�g�m��l�3ӫ%ƥ��7E���ԺF���&=�����\1|���lټ�AssuM��U�W�W�ޖ$�x�}�����|��O���8r�95��v��7�!&�T�V*�W�����bm�B�����DW��l�Tۺ��$�D�2�Hk1%����n�wOh��\:�L����-;��z�Ѻ�ݱw�����P�yM�=�C%�ٽ�a�Fd�z���7M�����E�[��� چ�}"?'Jk\��<����|���k_i���XiU&��W�v�>Rs~�����U�W�J�c/�W۱�P&^��g]4&���L��>4a�3�W��#���i��LT_�4���@`�n�:��*�kR
=L}<<�KȜ���=b��G�Ç@��Q�����XI�H;t�JӷU���������+>B��S�21$ZN95�с��=�+v��у���g4���o��!������G����"
�����eu�T��@h���bX���]&����
2g���F�� ţ!���V|�uC� n MeA��
Am*�E5�7N����ˢ̄���TIS-�w/ɯ�ǽ�p9���_�Q�
�8(��n���5��U9�Eg��ځQ:F�Yv]�������=�����	�>ܮq�>���#�A�#�e�w�_s?`��P8T&NN�f�����t���PF]9�<�ZY������C���z�M���H?�0���;E`��!P�� qd�ގ��P�ۇ���7$/��Y�-�v��_�G�o+K*Ӎ� �?����̮£�������a�5�l��̌�����#�^g��|D
�W��sA�R7����m]�@�ޖ�ں���6ΎS�̄Zpp�R�<q�ɦ0U3��p���P���-h&}�GN7=�c[�'5���e(����[h��=����=lӶԇ�����C�^���,�w-�q<�����������V�F����#����4�H��L�
���1�,��������vG����p�Y�c[8�2��nj�\�"鏲)(H���$�����(`�C��`[���{qЍY���vc}}W̍U<ѽ c�4(h���)����褳�2S��D�_A�8+�\w)��2��f����B�C�m����v� ���ckR�vR�b��J�!=z]�^�S���~/���rk�y��)�����|k�duU�UAi��6���u4����"��j��_���l���e��d�����ה��* ��	 kE4�\2����l'��o�#v"3�OF�@8R���T}��Τ����<�D���b�+��E�	�2���� �;���4O�n�o��r�GW,Mew�؃/Q<��ۡeW)�x���]��߿���Q����7N"7	�qC��y������|Ie"�ץ8Tp�豭 1�*%pQM'd��]�´(�	>L����G�g��S�Gө�!a�+� 5��/�n��/A@�vb}�J���o+��hV�����wy��n�;q���m�i^ߓۼ�ϵ��L������Ym��,��tTOي��:|s܃��z�(���6�5G8��'���"��dB��=���uj[��@o-�$���͑l;>"1>ڠê"�`c$zљ�L�y��䷎�<���6F6ٻ!D����FX���O���؆�� ��s/��M�?n]<42^�Wtc�(���Y���FP$U��`�;��c��\:��	�l��w����ݒ��TH������B�g6�����iΣ=y�<�LA�E�L/�-L��ib)�ٝ���^8l��B@b���uE �og�'���������϶Oe>zP�>|ؕ)��sQ��,0��:�.��y��
�
����:��წ���)��=�&�A���V��G���>���?��O�>L(����d~J`5��8�Q&�yߏ��ŉ�'����Vi2��q�(��Y�Bt�W�?���.'��d����(��j�k�;d�-Gbvefs��qd����}�D75lˡ��-@��>J^l����`�_���a';�!�wW��F��M�ۄ�K�u	��Kc\���ݚG�Jim^��]�V�Q��.��g�H�>��;cy, O�Ӥk�E�v���L��K�OpuSnC�0��Є�����E_h���síl�o�t�|�p�����ƪ�=�bb�����c-[����N��bR�u6��y��;-�[�S���~v[B
I��y鍔[E��{�uh�^�@��#˷����[������,��RʧA��x�lj}@��5�ˉ�)�J�+3�R�X2��6u��}��W�P3⍢D�#���'�����@�2�6���=Ǖ�&_�ɘ`_��9����L�{�U%���q�@��-e��K����ns�#�e�ھK������!������\��"��1�9A�����0��:�Ӯ�iL���ŮYJ��$eL�����q���Q< I�Ô�1��QՀ�>�q(��q�}r�&$�P[�C
ڮ�O�~�Ů�E���n�"�!#��Y}�}rE��:���e�[��N�����G0�.~�� S�%VΧ�j��\��&����3u+��'�-��k���'�`�[	:��/ס��b��f3-] S�6Λ=)҆*�jX�D:[�~k�4Inh���Qioi0���_�y>P�z��Pp�Y�������7�~HQ؉s�3���}}(��x�M�?p,Pk�;�/�R��F|*(���>ej4�����\n��ԇU�&�6�%V�y�I��DW������맪f8������U�ep�IK��7�.�����+Wʨ���C�	o4�1y�W�OG˂��,����<b7v�2�o����I��?�B���Ne���-���X�T�r�qВ��W�q��+p��BF&9����5��EE,�y� �փ�9��|ĺw��K�o��G�*`ay����m�+C-K�����s���aՎ9����z��ss�O���� 8�fՍ��I~�4��W��Aގ-[HXxlK����_�
�4P�'Ykl'����Y���yS��E���b2���UԷ5(Z�q��e:��m��J�	�����D�:�{���}_ǌ�og��^� ;k]��^��$5T��t��ƄH�!�9$�5�e���ۥ���
�WN:Q���-��ۄW�K���29.�������ǖ;8��U�
"����������sq�������d��;:�#�����+H�&�A�j=X�MzWBG@z��@�%��z�gF<�������r1��^k��^�}���7���X9�HK�+�ۃ��;u^?�s5��p�S R�h�mGX9h�m�rn�����J�=I4�Bs9L����w8*X��'|�5::�����%����%�I�j� v�oP����M�`	�e	@(a3X�)*Z&n}�ɉ���:A�,.W�����R]/����ğ'ih��]���qr��|�|�Y�ڎ3��&���p5�`���m�f��4@A_)��(.��,d�ѮNpȝ�3~o�pF���vǇ��7�~D~���9�������F0�(4f�ٌ��i�'��_�@u~��yI��\�xĉ���{ ����8
p�s �\�7��|���㼊�Q�'j��N�9�&L��{�o"���H"}�Y�x�e��@�	v�*w?����P>�W�O���绶��#=�l�1�3������>��F��Q�$^��}�'l�ǭ�׃�cm<��P0���s��O!O8�x�'*���F������C�s�X���
Dv��@�Ni<کP �>(�3�S�� ��ZX���=4�o>��fb-mݚ
��[� �~̽����
�$` ����ª����g����f�|��,�/-KCw�o*z�8�H��+'��[K�5��:"�3O��_8��S�	��� T��ym�B��� �À��᪺���r{�3,���t���ֿI�O��T`e�YN���Z[N\E��;����N�o�8��{7�ir�-��x�i��]	Y�bŝ�Xҧp=����9��4�\��x&�r���6���Q�H� j�`b'��G�%����D5Ի��_W��v t�)N�'l"����?߶6>����� �/�0��z�Щ��so�F}k��+�}%�oON(���tv�t��
�6��-W��I�����|�[��Ք���Oe��#���N�<�jL��~��]��g�D�a�����:�|]�-��$O�-�p�t����Jώ-��asNr������9as(]�z!GOF�`�G��9	C���%�9�~���\J�^B�fߚLze�*S�i|݇���5]:忳8�\=� ������n��p���#� &�k�~#�IR�s�6���w�U�5b�PvN��.���o^�	�7�ȅ^�����i��_��{��9�*�zz�V�����ߖV��UI�<B�:�Y�f!˵�*�aXqX�_OK�iv�8�+>>A\4@;⻋����&��ZCX��'�|����e_翿9ʱ����x�hzJ��D�y�m>l}��D��VD �	CE���MsN���h��{ߠ�*Pt>�jK2|�qL��
�SQrYE�d1�Ψ��xm}W_z3�So��
�Q�[xY�x�S�"_��݋����q��B֕�r�2��ċ޿�ɡ�X�f�x�tF����S�]Z
�yз�ϯͿ��P){��qj3����N��$���o� �Q��ZE#�D7�>���O{��ԧTDvܳ='��=�_%+V�g4�i�s��o��W���Wj�z�)}�|]�3�j�'N����ͨ)�סrЗto��|��r]��繹���kri�!m2�K�2�6h�����#(����Ni�NM*v���,低��^ f(�l��J]����E���f�q6�\R�p������u]�7DO� �N)(�8��s_��*��G��M��<����wD�V�����.g��������G6�0���
`�m�rC���������:T��F�:_i}U�-\!TޖTa�׆T����s�h��338�aE�(��7u�y�`Qx��MV!;�s��^�pvrť|>�%��W#
j��}i}�t,�qJ���p�t�\���d�4��)썢TrK��-x*y��|֔�[CCV�D�ia�w���͒;F:��0��5�2z��%/Z�]?�xR��ÿ���Ϲ����pO֞�HSdm�W@e;��RjʻJ��"�/�~����5M�R"����P���;�9�竺��V�>�w�q���lb^j��c��w�SS�������UNK��N�����̒����#''�f6������2m�R��Շ;��+����(���=R ��]]��E��������i5Cx��t������ތ 
s����|%��!��4�f�=S@��ُ��W�+\l�=��u��K4�he=j#6x��sNSƚ�.V������pF�Ԫ��L:�z.�!��B��Z 6��	����K]��B�b��nG�]v�4� �/gd�j�(QO�eiܴ�-��eB�p/݉	|�{U�)�G�+�XC�X6�]D����qmc6O����{)^M>�'�ϧ�B:�n��/4�\vl[iu [ǥޤZ�\��9\�)Q��EaU����8���b��t��,f���3��.���>��[��L�z6����饺�_�9sP�$��B{+)n��ԗN���y���S{�i+z��*�*
P)N�V��=ܒc	��ܛ���*י-R�u~}�bhY��D+{�g� �YP1����{+g��-$��_w�)�*�%)d] *5��J7��f��v���J�^��׏y��y�;RP�gm��$�����x���TT�V~+��⧸�Kg���}]���60x��i/{s�pAj�����Xj�N�ՋʹNM~kJY6���#�6e#m�i;�sz=�H�l������T�.�<?�YR8C���>�I(>A��h�L�{����[Gn��-�"�W)��kUJ�����:O@Tު�_5
�&F���yiP��,�%��.R���3����#O"�bqn��9ǥ�����J�A �ss󪥛��Ń>�|	�g�e�s��y���\;�Lt/7�9�}n#���f~����/9kFz��g���θ�����k鎗����k����L',�����|��T~���biq�J��ܜ0�����,�n�	|~���)�Ţ����VIf%4K�en�Po3j]��*�m�(s:�p�nP���r�~s���k۴j��{E�f��=��jhkS��4#D�4�]�s�%ר���Yn�� <�D��t������鞙+<� g-)���
}�K���'_�Zl��&��3���U���s�����z���̉�HË��k��#_@�~�����pk�)m����֋�ͣ��	�J3�<{��M{��E�a6��k��l�����wB�pw�L�z��Pd�s~g0-6Br>�R�5�#7��HӻeT�c\Tr+�,#�8ZW(UZ��ܸ]���;�_���(N����ǁ�>��R83�g�n8X�L��Ur��7v3�����F�f�!
�ˋ��p�j����[iw���{Ro��FgqhoE nҲ�F�s��u�l���(gI�d�^1�^G����4-�p��e���4dן�xYVc'6oո]q�<�#��痐���/��������JJhԶ]a�)�Ǐ/�a�قu;��l�T#?��\��&���pJ疕B��ޠ/�ঞ��k#�/}�J�K�5��⭵���L���cm�Ѻ���i`*_ܼ�u:V�a0�Ǘ�Dmn�����'�%�٧fN�7�2�[��5�O��"�t<~���*o���r��C������1���9=�8�����G�h������h~%�ǳ��-��O �p��b�����w�7{�~�;r��?zH�C)�����&�)|����B\��˚t>�E�<:6�l�!+�����/:�p9T�t�����v�R�P��.���XA}TQ���!����R�9�X�_��.Ç;��^b��0�|�ȭa��嬎���&>���7��W��{k=.��ig�jxu��>0�1�%Ct�y|�k���D�F�bd�p#����q�q�=��2&���,F�j.�=J��#��ֵ���L�z�1k�s�7�]ʃa'��0x��5�E����HJJ����4�7<[w�S9��.�{����
�Z֯���s�d=8�~��Ul�sNr�*��TB^{��y~+��v��6TATFn�����#��؉6>4�FZX���Ъ�_�6NUrXX�뢫�k����<x`=�7t�0�Q��88x�z�ͱ'c�{��͓���_��o�i�ޱ԰�G��w-���
s�p�ZOʔ��8�*l�Wy%���?�a��|�؃�E���
d�{�1���9�1���Q�����d|�+��Z9��w�>�nU�"�ty�DG�&Fȧ��5�|]�[#�>����t��P�ܗ���fHf�.�~�2�)�$��!�N��sF�~��X�έ����l�$	��K1���yx������Uʲ��͑v�}�.;��}����i�����_��si �Z�';�������n�%�\b&��f[���7a~�ܵ9���\O��2Z��J�1��'�ճ� ���8��眺��\�KBw'�?b���(>�-F��F@-�����0'|2lH��?[�d�(JN�uP���U���j�]��3��2,�V*_ʟ�u{	j�D��&`]��*�f{D�pKD)�P�o�2�C��w��/��ϴ�j ��%��.8@\¡"��K}���M��CS�/��U֥2�
$����v|�̵=���pw!Kt/����c��Y����U�Fȉ�Z�.��&aM�+2���͆���zit�_c�z 0S0I����kjGQ��_�^qY�ǚ_�V�陏�-�r����
k@/�2�=�w�e����\rsͪ'�pp��R�_���^�]���Ww�u󌷧�<G�ڴs�(�c�xk#"y��zȤ�ɳ��M��p��g0��v�ho?b�������@%�$>͟ي��Oh�7�F�%����ST4�t׭�e8���L��m&ls3�_�h������#���>JW�!@���|5�Gq1v�
$ไ�0qq:���=-��j�\8>K1 |����ٮ҂�C`^�bbN��ņ3-}�K-)u�v��=B��//��
�][i=S��Ao��s�%TFn
��81�;?��u��q�b�|�^K_�vh��L���f�������o�Q�[XS��7�C}�U��tS#JI,�aW	m�@�
��R������@�m(Sv�=�ytx?��7���kZ�c�띯K��뢡c�_�#zAYV2���u��P��ڳBf��IC �[���1���c��RG9|\[��$e q���B9*�5{j��0h��f��9HQ;25an��"맛�w�+�؂��e��ݍ�B�r'm�i�3�=��*��Waq��Cڈ�W�Y�<�zur�;c2�v�e�#76�剗,11 ���fOR��\��%+���_��Xz�����i�I���Hx����x�����z�{ҫ�	��zJa����T�w��Q6=�������
��:��n���|Մd�9�[g�KKj�*���>��X�b<כûeN,��L�*.�6-y�������J�r�ُ,���� +o��k6�5�:��1��*����z{�l2�2�\��9OHR��E��c��A��Y�s{�<Þ��1���c�N$��/��g��^[���Hd���1��{�͗��1�_��O��l�E��{�#d:1pQ��W�S=5C���1Ŏ��'��wh��H�K��{,��JY���G6F).Y���*���4�&2F�?�Fc�$Y����S��h'\�����
��ok�+��\��������6�m�y�i�,��Ph�[Ë��8d�Lڮ�R�h�i��"O� d
SOi_`s�u��oY �]h��7����*�
K�[v�9t������C\\��1�Z߄�Ϗ�\|�ґ�P<>����Pv����U_]�/�[0oO�U*�]�Ž�=�86�+��[�.W���r�Ŀ=������#qo
T�����)E���NҘ�tp
�n�d�=��4/����8��B�9:����7��C�#=�bD�9�	�R���ph��ۣۚ"���fչ��>X_�ă����_���J���ŭ�
�Ш���Eec�|�v��Y6_���R��+���p~��$GO�Ͳ�ۋ��z�%pߗ��ͱ�F�ӿ��;��_oC��<v�rM_�7�Ȳ��g���m���-R�;zv�����-h��� .8*��	���q�|K����
#g�y��2n%�I@ ��^����9_��e[|�Q�`�RSNw�r�A��Jca�͟�퇬��������J9�LKys1�`��➕�6�CC꧱"��r��ND�23���〽랧*3L ��Q���mng;��7P�u��բҴv�7^@,k��/�ܧQ(��d,���{3�a;NR0�r0�u��c��=U�-����h�Z..���ZqF(ZA���ʺr���E�/Ĥ�� ��{o���z$yѣ⛗�-d> H��.*��~��S�E��5���1�^��{M<�=y�*���<S�XXN?i��R�#�R������C]^��!����9�����g�o#�����-OOym��]}�6:-盰�����|h���o�Vm,�;����������`�qEZ�U_�������	����k�����z�}\E9פM���5e7p*����]/�2O��GuzQ,Q\͇i��0�����k���m���6�@���K�)�*����\j���u����w^�y#m-B��䔢y䲆~����A~���	��)�Lsu:�!��:c�I|}S�.~9s��v<Ztwe�a��mc�ڥQU3��B�$]:��m�dtM�ao��S��������D���b�A�"
�^GJ���Ui4<����(b�4�@_�af����A)�,���r2����ae}�:�Waa�@�qlBIpj7��6z$h�./'p���=���{��&35#f��Z(9{��b=G-��CG��<B�b�u���$�u�gC����[�lJe �*�2[fY�g��\���J�eO\�G!>�aѦ���-���=_�d_���f��N����u�����$�Ϟ�1�.6+�-&����ftK�����iI��\U^��S�A�ث�ùy�T����i
}V��ľȿ�n'�C��Pdi��V�sͲ�޸Bj
���\tM�*e�2P��Q9/�[�ͭ��:^Gov�N�C�7~���mA��ъ��7�o���%yD~���A8��q�3��μr�nn8��v�9���'������	�<�(�X�̊��+�WJ���=}
����y��q���Y�����_%sp�X��R���E����I?�Q�s�`������]��A��wJ��R��a/�+N�4{;F|�m������d��W)m������ǣ��f�c&GN������DQ�PXVV�ᬁjUn����?;��}����f���õ���5yxڤ�LS���n�HP�t�;�?�tB��1%�vEݼ�T�l���W�5r�O�1�t2�Z�ܼ�6�������pi`�Rx����x�ľ�o�?O*I�"��x���8�q�gynu���j�>cL]����gyyy5��ϟ�w�g����rϬ�w��/��ln[��U~�� Ť����v�}�u��^��"�YW�U��)�s �%�j����D6�l�'XTn5��@l��/?�;�-����Y�%��V�s�o?ؔ`kj}���?3E0��it^�f}�E�F�����gO��A���?^>�j�j�k�+.�w�FTߐ�����\k:��Sk����w��(9 �iB	$��Vk������x��V��Wc�u�T�U*�M9���YI��j_�l.���8��ʂ���\������f߱�$�9���9�ǌ=��
jȭ�wi��O��8��|�@Ϛ��P[%@�S�R��rK��|w�e��ć2�WP�!pd����bL�\1������:�k8�#QoL���s�H���TJ���Y������PB#X�;�wa��Qyu��pLai-��<55�$dz�I%._���	LF˔��u�Bl(C	���sV��rN��F�r I���-�p�OI+y3�.^��ǧ���;��Ԥ��j�)�����^����Hަk��Z�����f�q6����}%�3B�-�N���0]�lHH���N����T�f�����܇8l�!MpȲ'�r�mZ(z�U���WN��m)��I��ԍ�y��)�gа���[Ǜ1���%"�q��6&�oψa��R�Q���B���<�L.V��O�׷y+���{]�vH�~O�%��!����e��7�1�n|�[7�B/�j^�f&%i�L)���,?�q�l6i�ⅴIH�csꉯ\��2�C0Rg�l y�XT��l>>�/�&ƍ*;uJbogN�������^
f�+4_~��DNj��V���:�0�t�y�}�/�5Iܺ_+�s�~�ɶ�;���έ՜������M�w��d��gҍ���MY;�wj�~J��7c�&��O�R�60�=�E��2��Ÿ�+�~y��# р+ڑ{��h�O� "����k�ۨ��!S�����_sD�gw�r��B��ؼ��WJ�S�G������ޒ!�hc�2;J���>���x�w����g!�����]��H�Nmd�`P	��Nf ��z-)l�q�g 4 ����"�t�J�����?�>T�Q�`b�����r�5�����R�cS_��TTI7|��d���X\0ۑCҙ����p� ����O"�6wT`��v�;�E�8˨��z�;�[�zI&��lI�Q��[�[��:}i��� �ӶWq�I�k{ύg���?�u+8#@�(�� �B.b����VS0PW+5�Ch����J$�ĤFH��pv1���Z�\16!U�?¡"����o�~�������w���{��j�KYJ��ZO�Mut�������?|>'᫰P�B��4�녫��wUǯ-���v�k�0�xye�0�@�����O���~h6�6.'K���w��x#��p�a�Jfw�g��ň o��^�b׮���=�~��yA� ���M�������Е���9�ǃ��ۄ�q�a ���M��yn/"�؞�tD}�ɳ��n2��TX奠���ϿD�����L�-0� ��}��'���~0�1�q����j��_=`�$�`�~A޽��C����߯���������������z0�I.|�i�)�JA��`6��|_���M��J�ȝf͟�6��l?w��c��<�h;���{0�Ն�3p��2���
Jf�ӝ���?�ʬ��$gV�N����p�P�ȍy�c�-��x�u=���݋�S�7<<�g�C�7f�����܃r��L	;>(2�<�e��d��y9��k�8l�D�|���Ls9�a��O$��� wG�>����	#��P���6
 mbC��s�>H��t�v�^AVb���,OA9x�����[���ܰ�MQ��%�C
�?G���z�-;;���o�{����J�@��JG�iq��O���W� ���� ��s�Z���q-�Iޤɟ4�Ώ:���'�� )OM�Dό�;���-]�+��Q�M��0Un��o�P.�P�� �����������ab�Ә�����M�81��z�]��2�2��l�{t[�#
����\_�O�_WVV����)2����Gqƻ3<)"8o6�bĿ������O�rD��*}�aD�9z��(�|n�"iL�jfc��IQGG�8#"3J=�K���٧I����nɂ�����uN.��{����0:e�����
��a�Ua)v(//f�Ġ��!�3�W��-Yi�x�بhD�4���^M]r�b�� �}�A�����%v�e��2$ޛ��N�I`����*B��_�^o��~nY4~��k���7�2��ʉTډ1y���y����a��q1C5T�ݘW��˳7N�(/#�'}�..%E�H^�}:��l�y��,��t�]W2��Z8w�TW�+����y	�j������jN~���,�-��P�]��Z��s������i��W��%��o��L��Z���󀀍����i	�9s[� Yu�^�5y���w[j�=�,J.o��+х{х�6��������[��դN�!��4�\��S-=���4����ܠȄg�����[)<�NYcn�Yo�IR��HH@ �۪�3�;�^���P�:��9f%V1�z���L�R^�%���\��(���PA�D(.n�ʙ�'0N��z�?��՗'����@#���;D����꼽�a@�4��юo�q��Aԡvfr��5d��LS)�B�:I�{��/��o72u��Ȑ�<�)N����p�	D{�/&��ag�i%�B���60��g䎐�Խ����!�Ơ-�%xE�W��� �����ug�G�Vr�K�n�{4��.ne�5S+dkD�"fo�z��$;N:a�P
�Q68�8S�QȰ�^jԏ&v}N���V��VHe�� fB �E�q���ӣ�D��\~}?�S���!~��l>.򸦣� ��z�q�e��_'<SY��oL]����_����ĳh�ʫ윜�V߂+9���w�����ws�O<u��\L��3_��P������vIJ� ����}���o��(��/�Ԥ
T^ı�޿L�\�@��!�=�D�Q���Z�{�h�����G�쯝�R}�bN�{g��������-o�}磓q>s�Jg��?^se{�[�$�M�*W��"���Z[W+��Z,5B(<9����,��h���(����n�*9��5u��;]g���cE�:fH%���C>F���X���>V��~��޷˳
���BL��{;i"IC����e�E��G�e�A���OQ�,*�V1�h_3�@�ی���z�'݇�#&�i�,� �{T����E]9�0c箾��'1�I���8���;���^K��/�U[�6�)_�.|��z�b��I����p���eO����\	2F,pM//Y(����OX���Sxkp�@+A9���08Ed�`|^טC�� ���>97;;��3D�-�BdJE��5�n�~��?x-e_T�cr>�չF���Ut�z2�ޕ��7��Z�fte𗋱������L��Ɯ��,�#.7�򢒐ƕ�I	����&D��6iW�3d[�E�P�I�Q�=ʽy"i}�P�1�<d�}�f���5a���W5`I�Y�̛Mm%���}��Sw�S|1ߟ��5�O��<�頩Zr�M:�o� ���j�+^��o�u���v�����0uߑC���0�>��C�ζp!�"x��ܟz-����_��/mxüㆆE<�3�������b
��Sto�8h���ˋ� �\��'��K����<������rS��U��	�,u� �I_�t�0�mWOv�~���4EKm�/F�%>y�ٸl	?���W��.�,�y�M�ջ�^�TЉ#�ڵ6�LÂ{���]Lֽ+&}�nJ��K��n�=�h>�a��L��/��f��f�Fh}>�_�G�5X�#��� ��N`�������{Z������$���9L�q�2qM�dy���S_��3��s���l/_N'O���u~H_��ī+����c�?y�m����M�����&����@V���������������+	@^!�lCS��K82s�r���+���κ���3�b���2����Y#9Rs����T�^]���9M���Ⱥ��g�������>6����g��#�CG]���)k+.�����v҂2K��ܖm�MWH	��ɸ(�Ғ�5n�7�HU��A���4���aB�.|�P��O���F����/-��抱1;j�,w��<�93�_�wurGWn"����7��lr�+�RA®���ß������5�1�Z0���3ty��|6�g����T���_RJE�a��z~7dN
��m�*�@=��u}�ꇩ�{�11�rn�&9چF�{�-����b�K����$|����hOg#_��rD�;F|sM�YA��	���g����餤�}�tS���x��Ӌ�����3dH�^�8Ѵ��_�j�N!MNL��a ���K�o_=W�Æo�]��n� ��)'l�hi�����I���P��X�AF٪a�Z���d\[K2�ߝ�+�2���S��]�[tU��}L|ds�I��Æ ߡZL�Ժ?Gr��BD�w,��.o%:L��,�����ƿ�b��7��|0�uP��A/���y�ds���J��=��a�=�K�`��L�U�	X&L�h\����L��K>n!���"(���@G��]Î\�Zzwm�f�& X%1�q�.�<*U�̓mt^f�Xb��ykl�rYVFa�����?t{0�ơ%���ˊI�뺠>���k��d�E��6;t�)f'~���W��m�'L��1+|!�ah*��B?�U��0�s<�"�����t�B��5Y��+A�v�5�v(k��f�a�6f�vsm/ōM��<Y8��#�׷ΑE�ڕ+)�`�ۚ0�E��8�+�g���Zx�җ��2X'���[�}8�1Y��Ӵ��wj��UTS��;Ni7���˗�5ٕ�e��e���]�6�1�:��9H#�
�M��k�m�r_&��#�M�;�����cw��h�+#s+�M�^��}@�${�O������'T	��I��CS���dXDK�e��ݮJ��~���d����	�+��?��Le2x����������9���+X�D�z�(���y�Nrw�;���������}lu���� rݽ��b��M�#�dc�L��1:���佹@�7�C��8Z�hw���3K=Aw�o��=�V�����-�C�O7��
 &R�6�������	�-���Q��2�F΍�l��=����u�y��&�����8�)���9��ir�.@��˸)zS�����@�>-w��r��;׆%]�eگ�L�/��y��MD��~����z���8f[�4�L�@=��8���:>kN�;Ϣ�k�3Y�cX���g�����7���R������]nQ���uS�C#=��s����ϼ�Ƚ13��@� ҘJ��J�!�o"Us_NI��}��o��U� b����:cN2�`�Sɒ�X �!��5K�s]��F�8iR�^�-����p�N��g$(D#��X@�O�wT~�ԉ�b�&��d�PDF8{�!މ�X������1�B�,8i����5�\Į,*����V�l6J.t5��<�j����)ki��%����,̆�U{�O��t���V�ߞ�v�+?l��ˀh��]LT+��:��/ܽ��ꗝ0E#.	��T/�a޾Pa>׽V�= !��T?z�8�!�1�ӏ�23+Z���o-ɉ	?x�qN�5�N�\�Ї~���lWF�1�w�á���=Ɩ�J!aG���&�;fJ!sy�F��ŀ�h��
F�I33���J��*����\."Ϧ��vw�t̑����c9���/�R���/�LY�����B��Ҹi��(�r���imUOBh���Kr񥾂��I��
C��f�vK�
�� K��&�~���Q>:�G��m��|�`�LF��nmH�0@C��c�f�cXIϒq111��콑������f�"F��-��P���]�w����X#u��VT�1uLZj��6�+�ů^��<kXn1X�+o���,Z�~��V�y����G�!l��^�W�ab-�L�t���z�����ڴE���snD�#��{x�ʝ�w$t9`i��s��=jѪP�f�^$R;�0���9h�\�R ���>�0�1�T�P1_�k]�5��~h4�����j��k�T#�1i4 @��}�c>H��\��G���x=�j
XA�*��h7!wg�j���ߪ�0�7�cK/C��=���lo�r��d+�2�? ��.�U��_:l��se�-=�0-y��������uݒ��)�I�rI-�.Vh6	��=�BRd3c��&�^�\���_��FR�9Í��'EZP]�����k�{n״K-u����5k#�6��u���Lԏ%%6���k���PGġU���d�3��P���㡪�7�N�A�D�*�J/�oK��7��!\�~
����TX�[w��j��`p�Do�t?�FC��z��/+�w�U�^��)\;��8΃��'�B�k�����	�z_�݋�b�9F�!>���CU_+X��}0l��D �>ZI( Ako��N���s2o��̋�ϣ争I�k�'��f�o=<����ņ��]<�!��7.ˡ�pY�
�!0�Vt#	Õ�D*��(1��L�f��Zs���`^���6�liD�v�*[4��[�J���#�u�S�h\O�w�m���uZח�%=|Ay�m�ث	�&>�ߝ�;+��̣w��}E�e���eJ ����ӂ�o�}v���}A;4n�~�IU>S��#��	6�9ݡzGQ�x�#U��'&�HN��|o�2�>ޥK����+oLq#�
�*F��kf˩�!�jMu��jk�F�b��^K�(��W(��
�2_�;3?�X�SY}�4#_V����4D|X]����5��09s�4oh�NL	K����㚦ebe�s��_T2mj�>��/��Gt�۞�-,��0Z3�d�ξԃ�`j�(��̥����~�X����w2�_r@ϛVM�=��m�؝�=���a7�p=�"n5^���NSS<�q*���Y�ﮥR+��$S�fDdƱ&�4٫3pd���/���
��h�t���REu���K)�~ڙ���(B~:�K�xv���~v깚�[�}���J��h��MDP������)�+ŏ=f�������!�(nT��{ #�yé�*��Ċ��E;� M4͏U[b=-��d���L��Й?5�
��9��L��.ϋ�zjc�،?h?�ͺ�*���|��^�.#�ۂ��j��"�((v2�,���9�!�ē�x�����ga��ƹҙ�d���KMıq�#�%W@-��gzK��F����$|�!}Z��ι��q ��/~�0�,�O%��{�d"V�w���֓*U~9�5p٤�l���i5��y��FW�ՀW^��A}���jj�+3m��:����D�v�!�.��`���C��"C��E�S���-�c����T.�&��qLM�>O�H_�<,{e�d�}�t��K�z����<�{9f<�iq��lTu'D;���� �b=�agT��$N��Q���ˏ3�N�U��,i2�d��J�v�C--����������oڏ�G����8Q)��\e(ki@�8��=t���AFL�R�*��(��H�3Buo'G�*������z����*dΨ�|��U$��{�!x/��f��$`y8��V�F�׹��˷�#w�R���(JcpX��O�����t��e�n�<~�nb�\@�,��e�.�c@�iLW����>Z5�1NHV�ps�gPf�ї����w��5x�\"����b��ZE<�ů&K!�J��8��v������^��L�)�Y�o�cy*�E�g��?F?g�Z�U[Cf�Y@>�쥠 @��m�4R7k������	&�O��_`�]r6I�Sֈ�_�<�!-����~��~Hvk��ͦ�c)�=Oמ�nz��P�,R54�?��IXPI�I�vX�"��V����ee2y���h������R.���������M/Ue�ݵ+6藍!v*R�ƀ��%b5e���ő&���/����Øڛ{B�uϞ4ZQw����<�p�}Ȯ4��}��5v�E�����|DlN�JՐ��� ��1\a�ӽy��b���N�7Y��Z���~�Ϛ%����k�'���	�;~|(��O7�w��`�\�N}�OY���h)9w?*��TWM�eO�XŴܒY-}v�ܖt]K}�8JY�v���I
���ZQ߂�Lk޴�ς9�Ƿ)k���̩�HT(�������[M);�.����3IX����8�Y�u�\r����|1@�'�c
ab1K��i�N�� �2��j���LM���h�wS�o{�۴�d9���(�}�h��l��o�j/0�Nh�7e��נ�E̾�ҀdWB�JC= ��Ê/����T����d�#�-f�A�z�8�
՚���ʞ��m�(72��!,���O%i��̥G`���/���9n����%�?B�|��6z��v�z�]8�yq'��v�.� 8�/�I�J�������AJ�T==a�۶lM�xF?���.��!5&�-�k��3����WaJ٤��yfd�Q78�����{-����.��[�z�!�v6�+o5����p��y��枺M�:~�
�3��0�K��K���Uߥ!�Sŵά��oJb10w�Q�b0�
oS�>>�J'�^�<�+f��3���UhXA�~��'BLC�(6��l��Z#3� �*�5�����:�!#��Q����lMd����?xgC�h��:u>i����k�fb��Ћ�Q�����s��W��fӫ�CS�s�����[z����8��8E���%������پN���#^M~7��6��o�?3oP�ۅB�����`׽&V6�����?Z�=�����#`���ϴVt�����SPX�x��ܤ)_����ʬEZ���7eŉa��b�tB��kߏ8B��
��tϝ��?�y<e��T$h6�{]�mi�
���X�Q!�J�[�w��9���A�M�!�,��R#��I��z��Y�{�]`�VN@�P�xv�Tc����yA���Փ��W��;�'���[�%NX��@�IrM���5�}kӁqjp�s��xNfl�7&f�oi�4���M|�Eǩ!օ���,f��1��%=L)&8�Yl�x��5a�����t���!��w�ɓ��@��?龻{��RI�����jÂ��U���{-���Ú"-r��J�5����@ɶ��<�^'W�e)F6i#{�s���#sk�}bǩ4�4����f�c��.�su-�'��݄y���&~$Fӏ	Atu��6��m(�d˙�^V(�j��ؑ�zE�����٠�BD��=�G�����4.���oa��-tI�=|B���3c�yM\�jy@x^,�����$Q���ЀG���R��Û6x<k=��}�䆧ԣ�.�~N=��.Q��]-d�+z	���if4�{W�/x~H V"ˬ��
ic�����K��/�� �;�qq�TTr���
	��Z\�@~3����hk��ok�U�JsCE%���OEq��u�j�ܹ��E�����Gp���O�LD���D �L��}�r9��w����O�g���~���(��%")�~�>~��s;�8l*�%��ЧYYg�ʎ�����uq�0p�� 54��,�q��>۽M��2�Kko������:.�y��iiii���Z��AQA�n�.i�XBEZ�إ���Yj�������?��]��3g��5ל��گ�2z��si<\R�Ipٲ�{;sV�>Q_:�qr_Bd�#�`t�˯�ˎ�Ը���&;9��� �Ǔ�l�R�~�i�[��0�޽��Ž(�HS�iIU�a��>ҎH�!������3�+5��>%w�?�u�Ah�Em��C��՚�կ@
d����q���-ug���p���S�!�O;�{}%���+W2� ���U���J`��"�����?!�3U�'�o�F�:�����q���]I��,���4z�3�o���&c�Å��i�3on����	��7���r6�ȃZ ��R��ño/.�ūR�t���DX�N.8cz�}��K�upac�:��쐖�ΩT]-���=	)iP�m{lJq���X���j���T���d{uNee����I�[�
���A"j8�7&�Ǣ�	]k����m]j�	��j�yf�pl��B�j�ʜV);o=�P���		r|Z1����H��7y2JZQ/D+�_3�]�c�|�	�Z�r�q�w�(lnp��)FU.��hɤ|�U�H=��N{g}�y�{�ΫU���g]�3�?{��?������JO�T=3����Xi��5���X�.��V�8�w�w��rx��濐�AL%)�L�e��<����i�ӤQ��������J,8|x��dV�j̈́B���ao��;N�� d���q��^Z�<~�,d�yη�=�#��������O����LK�r�a��~���@;_NPh�0���/���G`nǯ���o+.�վ�bwQl��	�A�Wm�lw�����w�N��^��,GRfx~5	��}Qq^�K�*�խ[5�p������<�a1����&=�G�ߺ���W|O�D��
�4��5��|| ���`��e�3�I�>E�|Tb��7P�z���L'�;���<>��FF��+���;U��s�4\�z�й�v�/�Uu�T^2���ۗ4��e���45��-���I�a�h����Aw��hӷL�E`�c�	3���f���#7���C��'3t�h�E���A�3��Ju��p��Fff|�!h�:�t8sQ�@6���Do��mڠ����/��x����񂩡�
o~��G����2�w��y����η�(cF�����Ԁ����u������(??Pê�(�e�znk8�~����8h���E�S,��ţO.����P�
���PqR�0��-�� ���:D�O���wN����S��у�g��1gGeĉˋ��'�E4�*��O�g�ɿ�	���7�P��o>�A��⻊8��9ˬ���-����ԙ���[,�/2x�+z�w���ʑ
���
�[�I8&蒵��Tۃ=�����9��r�{���2;:�j窴o�����S�*6�|�\-�Ho�[�A*�$�d�Q��I%
�����z����:��om�c�!�R��B�Ӵj�����tߴ�éO�z/��9��vs�a���A�j�Hc���nH�a�����Rs��U��|��Xoh~�r��I��s��0�}�2��(S� �A��yo�T7�����=t1f<�Ϗ�b��`Yƻ�h���F8���졏���g�_�-[�x�m7-��ք�7ڥE�@˴��2�` ߎ���O^�I#AI���Y�Q�@�곐�y/5���[�o\n�2Q@��k���3�e#�����U��"�g�Y�v6:+*�gI�F��7?9�(#�	*k�hWhUn	u���$���>Ji]ڋo��� J�oΓ)����:��69�Q�m=���h�7��["��{=Q�\�Z�.�*X���<=���L���Zk��B_a����}�T�}H[��.'L�L&�����2}���Ƙ�L~�ylf�E/�mkP
����M0�4MP���y	�G�^	)�F�z_�Ð�I"p�e�s��P�_�.�;MC�!\l�ǡ���������S�wn^Wv�֗WCN�PD>�x�O�#��O ����SG��7�։B�;�g���w�u=�?��Z�hK����=�򾙙��^.`-��������/D�88�f��8���7.����❶z�ځ� �}�c�Z��X���s�mD���@@�iQ;��F,�;2��͢�<�{���굜����Ǎ���ߊ���*9J�غ˷�&+=z�kΈi&��2`52�+�y��|��������0�Dk2T�]-��\��V�C$��O2�o�����@���ږ�OJ�9��|���zM��x��Z3�+��� �xH�^����}��ί�iGcj��3�d�7�Aj�R�ߵ���pf�fO�mͳ�%�R�]�X�C�d�@aO̹�UIv�,LE��"�c!�q���/�M��a�ψUj�#-}��԰^�l���@,���B����`��X���9�s# |v�m+l�|ߝO�a��ð��Y������_γ@�f�7,��<8\�c���kH���'s��yCѢSr��D��M�[�:�+`��u��/6=(�X�AbB�7�GD���Sr�M�`������״��*�/(Gt44��{���s�z���2���Y�&/�EƼV���˔��1�¦M���	��-�:.9*�!�]�
f���jij�U�s�u�s >�*���))���st{:�8S����	������&��Zܹ�T���[�
��D���qo�8S���N/��:;�cF�2^��!S��۫W3⍱4�ls�-Z��&�,����Cm�%������\���r�_3 |���.y�����y�*y��� �*/�w�������4)�!�O&o=0m���+ǆ\����:/^��P௦%CQ���TH`���D��oin��N󩡕v���W����z�;��D��tF��
�SQ���R%U��>L)t��>��HGWc�4ßz�8��I�⸳� ��O�#�q?�g[э��QM����<e�g����͉�+dAڼS�T��L֎;�4��������30`9�����#����{7(}�2������M&*W��x��BÌ,����&����O��.,�XJFE� ��;��+'�w�(��Ի��c/?����Q����\�w�/A����
f#�1أL��ظ+n<K{�7"�<���K��2.*r^񻻄쿛�)t֪��`���v2�"���U�5#��,�.q�6�-P�+�**��_?��<6�l�
��K��+E�S@�;�=܏|�J�r7��J��W���U������Y�.fJ֖�R�ܥ?��Pz��E��*���l$ �t�-@���ǨEj��(/����y{22�����Q?�mK|X��\'sQޟ�`�?�S����>z�q��D_��&z��z�_�.�G�o<��֜u4�Ǒ-�Gb��hV��9+�(;GK|p��7�� �9�C3�7���.��-��p�|��t���f�<)�4'�8�]�jqb����D���C��0��%�4n���4��O���#�9�$Y��6��N$���S�Ve{М�<2%��&��v�\�˓�Y�"3�j�S��?���L�p��	����:��{�%ΖI��e0{���x���I	%ķ�;p�|8i��f���VwBG�����QQ��4y�S\�{̦���ֺW$7J����N���4i��i�9�!3Y���&�� �E��q���yX���H����>� L.%T��Wϛ�Pd4b�oX�_z� ��Ðm�����r�*�m������\�h���� TO?�����S!�cGٛ�u�٘����4��q�lw�>�4�W.վZ�\��)(��f�vZT=�R������C��N�m��T��Mf[���K�`Z��q�]���Ch�*�,���r�j9R���4��(d�Ho]~;ѝ��2bQ�M�Tՙ�JyS���u"�?	��b�ђY&���^V��f@�Cixtc���M�0;�����ZD�sWg����j�{x��^�(.�ei���?�������Ǿl?�R�:́�'X�>˂=�)~�i�{�\�^�X�>3|�AIQɲ��/L"go�\Q!�� V��������:���,.����J�


!�9�m-sz�FV^/�憖i�ЊR�ߴ�=�2#��d�?����� ��� \p���Ħ/�8����I%�s >���ǳ�a�ue竀"��m�ɳ_���U��,+�8`���X����k���č�[�rLr'�:/[�)G���h�3�/7�%�����g�5��?�쿼?�?�����M��8;V�S�*���*`�^�4��<N`o��R1�����rAG�����&_ݏ%]����C�%�_��(���z��)ѭ<J�Wll��w��2MSnb�±1��Ɵ�o��0Kk���E�Wv���FQ�e���>z����Y�0���� Wz��8�ښ?-�8=��tF���k-'�8���!��	q��V]t<�&�u�4���-�g��^������=�ۣ�����
E�۴�����e���LP `��r3��^eIgk̀����L54��|;���������.oݓIH\-�4i�6DU�i1~`����ƍ����,��	x?��[�Q�[��6�Ƈ��]X__8�WFn��+	d'9�XX ݴ.JA��Q��Cy��i�@
�;���N����b�asDcW�U�N��z����/q��:V�X�tj�(ک􇢑�_FPm$��qu#+nT�
�ޞb�	�J��|�Ţ����a�/o��K�ϛ)�Pc㎏�=�0�gt�$HG����%1q���?�����;��V��k�b�2���K�n��DU��S)dr�ySտ�D>4�pW�ߨU6o�sY>[�*������g-�lq`�n�"mE=�=9渢�A4U�l�.�|7};�=S����`�=���L]��呐@��)�������Uo_���uR�:�P���|y�Z8UU�o��3�Vd���{�7ب���6��,��-S���(�i�ҋb�nqUNٛV�u�:�kpK�4l2���{�[A���Ӭ���k�Q��KE�Q̑���:N�VRWqs�:��U��h6_�Q�	x�G�0�V��롡�/b$#(a�mn�� kI�gR�bmC+E�u�*��i�2��t#R�	�[),��\b�l��B��?���I��9/���h�K�!!V�ʱ���W�ATG��B�?p%i�
�F-�(�*�H҅Je&8�� �5���07���t0���c��&�EY��<g��N����"�_�<ٝF�VV�hՖ��������?�k�ywl|� �<��1ʸ8V�	ĕ��i�+zi��&%�QO������#w��G��@�ΎJF tF�L�TrpP��B�C�z�7��[���ŵ��-�~�lR��Ɍ����<Xf���BAAy��65�H��{GtC�+=C��Mǽk*Q��L�땅�[q,u� gh��d!5�Q����$��w/��I5=u���i����$���H�[H��r�q�
��F3�}�h䯳َдQNr��.��e��Ph�l1���8��q'��
�uD����l̆�M����	�ˮn>��ET��D�A��)#~ڵ�y��z&�>ݢ˛2b%�L��6�q'�����癝y�O��_ˮ��wH�5G?�Jܽj�v�B�5J&W��2��a�R��0��,q�XF��y�
��`e�X��G�O��Ú����y�ӧ�x�<"�b_E�X��#.̆��Z,g_]�PH�����U�~.�;��/��,:��S#'R�&�WH�%��؋e�Y,�1�$�aŹ\�Je( �p���3��������X��w���}=u7�ׂ�ǃL��rO��mMG߇[j�2JeĊ
3NBo��
���~Qnv�<��W���ˏMA{��Hu,)���n:h,ޘȟA<$��8=ߨ�+ܬՓ��ֻ:9��0$�R=��@��X_��ʏ�<G��������Օ���g��t�����hE�㮖p	��y��Q����Ɔ��	ݹ�:�����tA�Ck}���['��u��;�%�e��N�����4@8�8G�Ռ�ޅ@ ����˯fXc�6���@7�ӳD������H{;o�I�h��<�hg/1k�Z����ΰ83�V�O�F��áK|�	ࣧ��L0kX�r�H�����t�nfZE��(;g���lvq��X��v���x��v�'�?TQx��HGE�2���h�[g��Rb]sz"�����@XT���-�y���Xl:\�;�4�l���'�#�j�v�\Q|���b_"��a����"�9]#�?F���NR�וm�����io��7u�u�`��_�0������� n�"��W���u��T?�H,��گ�惣RҎF9e�~�L�P�-���rXi�j�R=�� ^�V�����pH&���N�'P׀����=�)(��w����vC�S���el>>�ph�;�+y
�q��V0�]GsXⱨY���m����Y���U�U���������t�Bͳ�� }�+�O?g���d}Oz������@�L
2��E�E���g_�]�,�O���f��+�8���
u��+�邪˛��#�ʢX�I�lΰ��d�F��{��Ԟ7P��.�D���9I[� L
��m�`�X��#�7H�K�8�$��2
䮣�����,k�g�ⷣ��T������$A��p�\�Z������Ŧ��bv���`�sy�&�y\���^X�Q?[Br��/�	��g��&��}���&[(HεAN�iTq�-S��aw�.+��^a9D�_~��L�p�����:J�<jq��A> n�f"n��X0�,	��5Cl�1�P1N1��]H+���?�U)�K��1������9�s��X5SLė�|Q��g����Y�3����%0�%�~�z�E7;~��<D8���?-U%�V9��s�����_3@K&�����u�%�Rʆ�UP��<��Fq��;�oUڏ�N�����ٮ�tm��������C��ʽ:�}&�T%m�; o�Э��KT��JqD�ܾ@�b�[t
#I�)?�sq)AF��)�D|o��S���]`P��+LK�,�1]�FF2@�I�q��fv4<��41]Yc��F=(�@ξ�,"��t�ڬvM�5�وᝥ�T�S�3f�;�W���;7_~6�[aBo��%�?Q���L/N21��f>��.w��#��-R�E���?K�o���� �������o�/�Z�z9s��}2R)���{��9{`� �]H{U�p&��zN��,V����o��(I�#���_9	2�v@�rv�2����^���	�:��b��i��Α��0~�?����]���D	�����A�Ԃͅ��[�$�t�X]}��7��%l��P��pXЪ��w��Fo��8pIE��:0�$:��n�̣�d�OL� La�y6u�`��Q���ƬRbbd��8��[��DoM�Ċ�E5=D;������.:��ʘy��΍�Y�=s]R�zk��dT��.P"dן��h�+aX�
PMv��r�&��TzmP�5'^qc1�����	5&e��j��W�ƛG���;��c(\�CPm�t�i�Qӡ�W�kM;;�R5N�7<v=k#�@��t)M{�R"S�\/�����J���f�z��܈4�-_jh8:{���љ�f�x�/�D.���ܳ�� ^�i�z����~�B���'h&�kq��7r�������Qm�*]\�u�Kvp��Z�����cS�ݮ�5�v}�o�c����rY���@�������J������R�d��Z�$����H��6~uqi���"���t9�B:I�3f/���� }�W��q��H�,��FՓ�n͖�&}W�[X$�*�+/�N�.���M�Ǚٸz��<�~���b]|6U]K��m�� � k�QIK�u���29h�M�LK;Z�/Q�Zh��|�:�ȳ6MG2u�h��o�>#��<g56f�:�rݨ�c;�~��͜q��a�����z/��]��6��6�L>bӌ��FB� ���Fw�wv����ã�������/�2}�yF7�5W>PR^���r��I�
qtO�zv��4�ڨ��0�X��p9pko�X����.$'�L���x���g���*Hݏ%Б��|�I�>9�;���K��bو�@hBm���V�?ۗ{0����ҫ�84�LUpӋD�+�2ρ�w����~$��1��k^p.=�˼���ϙ�����+o�FS����۬��z9Ѱ놖^bRm����p2�ʁ�����#�с嫫��'n�z�a0��]4����p0��w3mu��4!�ƪ+���	���	���~#���Z~�WV���� �U��҄m�IRq�W��� �=>�:�e"�=�Y-b1�w%��; ���A��ہ���6P�6��(�M?Í�m-n�h�Z4���O���,���n!�釤��l�o>#OЛ��`���%��Rx���CK^.�6]F5V��0�\	-�d�On ��	=�,F/g���a/DlZ����Ӷu��M���E����|H�M�zB��#���+��Fo�ԯ�gMr�nN��-G%�cv�1`)��&���.���;!r+��ɽ޵_;v��1����p������z:����bo?��f�,�`�^�T�ׁ�W4Ue�
�4�=��
�u�#�cs���((<�Å�v�a���t���8ǈ*SI� �F��8�ԇ�����FS�����m�vFVo������UW:|�����{&ǵ��ݰ��6�-�yZ�=Ű���#+�߰d�F;r[�)��v=��M�H'�=	��
{�ظ��g S\\� ��P�A�-2]4���B�MU�1�;1n*�!����f&J��^�N��1�E��֮��!�����"�� {����qz�S��!�oY)�>�{H���o&��&�S!%����2إp>'!km]��?"�_���g���:��sG��'2ω��W
����Y���C8�E�l��>��)�i���O���,\#Y3*Q��U4�c��kE}^~����מ���(�)�1�vLק���n.��==Y��Ԋ���675��d��(b��|�?�a'0� �(,3��2�'���I<F�%�d׶f�-d#m=~��`F��q�xIh�D�����)🪼�J�̉����;Tuy��y�\3g�"R�2In��%5aI�+f½ޢl�t��Y���ڽ#ʛ2��Ŋ��2��A<*��I8��eD��$��J�q�Z��pjM!�LA3�K�-���y���0�V��F�$T ���h�H�HW^��N�\kĹG��^Gz��:�~�ac�����LM�CI*��zߐX!Ϛ`F �N�[�N�+�^�	��;�x��a�������q�w�c�Ʃd ��ew�,/��[��䷌.�ar:B�u�� �># �mA����&�������.��៯}>����CQZ��O�^��[[}��0���g�kY���ǆ׼���*��*�|�ɰ;8�j��׬�?��Ĩ;�����H�xsjD��ɵn�`�-dў���kg�2�{l�U����L��{���:��b8�hsB_9_���'�M-��MM�9^6 �.j�H�D�D���61\HM�����vv4�uM�%\6�}��V���Í�<?�rS�Nғ���px~��H��~�u�L���u���� ���U�h�{�%��yl�!{߻��YNGҐ�4�w��M<����d��*��lle�d�`��D�7�Ɲ㢜f��WB���J�����O,z)�}9躌�`�k��o���>U�g{6�@H���1��o����#�<��Ŏ�Ђ�!��^*-�-��������hL�8��w\�޴��t�cJ���{~|�W�	���x�+}��C]��8�w����uz�Q��D�̇����������J�љ
�qP?H��2N���9	��o��ut6�)(�h�2��Q�\���v5�徆�y)9�th|����ȷ�B�D�j��ğ؊!M�R�U�^S�7`�����Z|��N��<�����p���u�3-S�0X�Ne���gj,���r����0c��MU���/�j-�EP\����E�X�WKS	������ ����LrXCDq��[�8k��/D2��$����m�< �Wz����Zn��JI��d��棶����6�o��;��U|@$�����t^{_`ڧ�}��Ua�)��� NU�1�j�Y�7��P:�/�S%�t]5q�6���E�Z��b�&R����DCRuUOT�i0AL�C�x=I��.X�s;�����Xt�ǂBQ�c�T/3�.j�'oWk�o V��W���:{�n�~ƈ����e���-_`ܭ��p��Ci��b�n��ݷ��w��o�#�3�A7�N��,ŕ���3�uc�s���T� ���q=��2�7��/�1m�kOؼhhQ�0��F��Q-����O4H��s���~Y��~�Y^Z��&y~aw�6�)˾y�6��m��`����_�����m���y�e��70F��y�˙�UXR�_���ym@/�c;�&⣪>�LM��x#�������Z89���.�
 c./��O���iڟ���έ�� ����1����� j��$Z��-|�*�-63���L�g���:�P�G�a��n�w>��-x��i#���Y���Px;�)���nIy���y��7h��C�\�L���3�a0Q=�-$�d`��,D�WX�W7��ì���{���?)/�(H8��>"b�K����'�ט;�W�G�"SL�E�R	 ۼ 0
Ў�>I�ڔM������ӥ�;��i�սt�Sjtr�6x:���a���D�k9��?�{���7�o|�XgE�?�B��3�BL���������m��;���WQu�N[?���o-K,}/�1G��AK�6r��ʮ�ۃt�K4*l� �]i�w�����8�w~m�:�� ��ra�j���_Y��[����v���eΊ�¤��I�NTq(Y�����Ǥ�	ٙ\�/>t���&u��*�c��;�@���Թ���D��]!v�3�4�LO�~��p��Wh���lB��e~]";};a`<8�޳B@���(S�1�0Xߗ���;C�๽/\��L���ؑ�bb�2$y��Z�"�-�t�[�-���i[V�c�bV�Ox��1�{�׀Q�&��g�rbSD<�R�;_�j�bt��|�5a	��o[D����'�Gg�F�o}os��K�W�~rd) 8!���z?/:cV�����;?�ؘ"{��`nU�0�I"?��=,�!i��]��L����Ӄ2���J�=5! w�A�%�HQ�/�����km�,^����jZ�P�nt�S���n!63ÿ���?LO���	\l�O@�R�����)h�&AM�5��.��*O��~���k��B�XV���1�y������Ʊl�������*�G���������;�y9�f ��|��E_s�������O��˒���8�w@�3�ƻq=�\��&������,�uyiR8��A�8|m�v��I��wC�_��mI�,60�]��W�0��� S�3�`z�թ�h/�P5�ԥ��'��;;��a�>����4�����5:�8�m�O4�����v�Lg�y: �	J���?<�`3��Ȝ�8ɹ!U�zսa���܀���X�1����D���|#�G�YT�{E߮�f�o�f(� -�����NDX�c���Bp�Xܯ�qK��OM�0S>��1qI�@ �:��REB� ���s�)�r��/���*
�'��#ɹ��=?�E�&�{I���9�y�P+*�*z>�X������a�{���?�5�1�	fC��4�wR��ԉ%��į�FW64|�мK������!��p��gj3/�b�,�r��'?���'xZ��`W�
:=�у�y^�����1T���nQ��i�1b��rx��Pf����?Q�Ȝ��fs�OwN���VG�[��'1���T�!����6얿�n����Y�uGYY�3t��0���ݪ���r2�ӭ�,�Ǜ�.�#��Ӵ���8����� i:�茞�iJ�3O�z�č�e�Ԛ����OVw��fL�tT�k����=y���jd�;	v�UI�s?dZH��T?�.��x��b]��`�i���y6�g���;���׳ W�Z�h��SW�$Ժ���>5�K��1axw�20�R8�C�T�Ծ�v�5�e`�pa2�.���X�J;!0!�h=�Hm�Zr=�,5LQ��LEv[����xm}1ѵ���a���Z��2���ؒ�{�0�� um�«�4���'�}dk鞐؞xv<i��sJ�ݬa��J��F^��-[�<ŋPQ
��8�~�]�@E%�S���NL�t��ܧg�.��/e�?U��~�qH_Q��O�F�S�#N`4mA'���}I��F�=G���B^�Q򗺔�L�cQ�<�U*��(ں�qK�q���^���m����6c���� �ȍ"�{��)}������XR\S�yɄm8��`�o��<�؋S���I>���X�i�}�b���Bz�e�&�,[]�~Ɠ\���T2`=�(�O�I=W�(�~8.�V�"n��R����4z���~��T9�Z�In����f�E�/���h1�2z	ZC&2��=���L�����t������U����w�,t&���tz����{��mlU�T�l��>�c;ޛ�Q�u�;<�.�=NNM�sV�����-�׈�<�+�t�C�h���2�I�h��U�G��	��~OL�B��3�IJ�h����{�yQڤ�&��l�J������ܨئ��dhi�OW���z�y�uE˟Y��moo_|cJ`�~�s=�*�S�#�M�����q�@^6�څ�~���xi���.�k6s��gG�3>z�*��+�8�v;�|���g5��N��ݭ~��(6ARo����3��A���l���"x���AJ������-�2����"ûw] ��Ú��y�'��4�A��o(d}\��!���93�<҂ꨱV����M�%A;J��1�����������fW��v� >#��x��#,s`ذ�N�X^�Y�:���4%>Û��;�JuY��r�h�����L�%	4b�/�fL��t�*#�n2�?�&���p����+�q��sX�F��;%$Xw�]g�;Ꞝy���ļ���C�nq'i(�����3�R��r8X4h�r=�Wɍ��8�
}C�q*�CE��Fc4�p���,r��v	H ^�g|�az�O�k��M���,��`�Fj����S��>?%�� $4�A
�x�Ĝѻ�������@ Ս=ÄÝ��]��� ��ύ�5QH1���1�cń�GQ@@>Z�A��N:��>PJ�80�n�P4JZ��R\>�s�>�j4����=��ϯD�h��!O��btC�w�����΋������vz앤+��/�������n�{���<m���s����3�Y��?���˳p�e�����Q�r{����r��u���6׏B&�zy`z��;+&��ɶ'�s���� `�l-���)*@�8(�Mo�Y)Π�Q�Гǿ��0L��Ks�D�� �	
�Os��^��1����1�1�� jvG2��������3)�h�A��V�F+司�gd��ߟ���aN%3���h�߫��!o!��
�������K\1���s�A_�%N�8���^��S�/$m8�u<�Ӏo?��lOR2�Q����	��B�m紐z�j[�W�D�<3[g�o�N\z����:»}z�J��(V��s0�L..͛Ԕ���{���w���幨��Tw�����VSII���H�im���m� H�Ԣ������sN��ȕ�[�Ȭ�E�d��_�!\��4 �����Q�F�W�&R�ё�9:��p"GC6�8{��uT3{���s�_73;�����<ڲ*�#6��&#&%��,��9k��Gh��J��[;*+/ϺU7�r�<�!5�z���*w��ɏ�JX��dqY�Uֵ���.�P�b����(�dX�i_���*鋪[y1;g�_�_���>S�Rë�������:�b�w�ѵz�=Ձ��;�I�-�����s�&�?�Kj�{'���P]V��tb��X	Awص�*l���:�X��_�9)�����x'����츒�;z��� �������+����Ԛ�|E-hm�uyVBw��>��7XYO������=�}t�c�J_�7���5�	��� Sڟyb�4^G$�<���:,�'���g��o�< �]:�Jh7�����d��cD���Fި&���aŦ8cF�5e�B����Y���ڪ��;�Ν���w��C/�o�����N ����a��*)����4���)������t`� �@�R�H�"?�߳Ga�Q��V����V�����?B��&�6t-Uð�S-�a���b��=f��]��V�-m�T���~x8#��u��¥�^���KA>�����nͶ2yz�⠚�,O���:� (e�g���N��q邶>)� s���/PF��adrF�h��t���za&90_��=2e�N�4V�7��h�l�SS��%�?���U��-�*��<��}ձ`���d��ʀ���Kvm��$	��~0@� o���]�(�d3�R%ެђޜ����_kcdݣ���w�[��)j���29�r"������X�=" 
�'�
 ��ݘ���72("\Ec��H��
���˺{�����r`�8��j���r/��NB@O���۸-�{�[Y\�
����-J�4#1��=l��ž���@N�o�8��y�6'�������*H������7��������%�ކ���J	�Y`�����6
?������0&�<�q�9�=)���Cr}xe������1,:���E�����m���P�cI�0�����a�nI��驖E!S�B�����L[!�y��wj�	��P]4�'�\�?D�J� C_�������k����k�l :���v���j��\D �9ڙL���m�S�+g��W�� al�����N��M��%��{V�'�Nz:�h"R}�|�ި�:���-O�>ŀ�#Ex��OC����g�;5fO�,��Q&���.qN"<�D���
~���<�閤��D����,|+�)�sM&r�s�rNm������~����]✧���{y�����R懅@(�!��W�	�#���~�kZ
�Ӑ���l���_�G�Mp�>F�ptS\++緆4~������\� w֔��n��?j�""WF�L�Z�B�7�G�A��_�h�s���Ua���dz�^"O
w�?��_Z')��7�������]g�y�-��qY9��V4�W̎�=�p �­Z�M�A-�*��"�+������:�-}j9;�R��s� C�\h����46�o�3��B3=|�B�5lD��i�5��`��5��Մ?��߲��>ݹ����J>H�yt9O= �	�-���������J���1�Q��1��R cڲw��μ!:g��^!,j}�A����g���K4�i��eb�Y�y��'A��4������� au8�2�mE�v:J��o/u5z�{���oĻwn�{~45q^��|�,�&�_�%	uo�F�{�i��fE���`��D2�6c�,��8�K��梈W�Q�(c���"B�<aG0�SW��#w���c�Q񦑂���T��e��=��̓��M���TnjJ��c������?����4�j�"�a�ϞȞX]q�7���E��K���M]�b��m�Ҏ'�o��|��6`�mfl68����	�턮��Z��������v׻���x)���u�����Ǧ�U���je��,���f�N�%,�?�`B��ܗ�n�H-]ݦ��
^ދ�B�{�]�Phpj����\��49M��P��Q�-/�����!#B�oe�U�(��D�NT����c>2��i�N䜵e�W��O���p��H�|���GQ.'q�MA=�]�5vm<� `���l|�}������T��~���{��A���J�b�Y�v�I8/q�3��Q����x����2�gՐ�X�G��`�Lh��!M�����S��v�Wٽ�����N�j������>�/C��R]�\"('LCB�=��=��׽�B��e̐M����ۧm<�����]|��u��m����}�����?pqׂ�F��"�g=��E��v�we-{��E �g�YŴ����}���!���x���{KbM�8��oGUf�x:�7�JKX2O�<'�X�c� ^��8����Փ�w�c��F�q��&��>��Xv��[�����
5�����_�Wm�����Á|*RhSi=M��\B�)� y9eUе3�-d|����̟+Ii���hG���V��"ӫI�yO�1��I��m�t^n'�����:Ϙ8]�/A�׎F�(T�9�,v��퟉�K��>%���?�Pc= m?�G� ���z�<T<Ll������� ��c� xӥA慄��p����=�!�����,���^���˳ӱ���0 -����fڣ�uġ�U�8@sN��s�f���@�t��uP����Z����H8��=��Z���ከV���v��#����Ώ�N>��:���#��	��*���7�S4��X,��P�R������o-�"M�陸��M!Sg|���g.�|"SJ�����{̣�o<���01@!�_G���A���rG�����W�5�5�ߌ�����A��ng��nz8�߇��ޞ�����D�7B����k=�!K1Ւ�����G[�����(q���*nV�r��Lq,]^z�:��b��U�Ou��OK%��̊(B��J��^]�=.½r͆���{�˵�����ƽds�{��.��������#�z�s���x��9�Xၗ�q�d��O��hCN������$�U�pU{�~�O__T�/F,�O�1O��\�r8������������e-��[��U��K�g��+p���o����@h;D|�����y�=�QVT��`~�[q��x�U�Nk�����@��F��T��K#@0��|7��c>^�i��sV�؈7���x�s��a�����ms��F������Z�a����ue{&%�jk����jC1��}m�eu�φ�ϱ�pwƛ�;4~Gڟ|��h_;V��<l�j�.���q�:���0����s<�oӰGf.Yŕ��e$������_EfoZ����֮�TS�T�⡎�\pQe��)�H���9y���Z�z#�ț���G�̦;�I}��(V�%S�:g�&5�	F�M����-}y06�6�?�E%���H*�d��_50�%?��2z����I�T�1+S���Tѥgѫkz^P����=��*@m$
�y�UP���Q%����,=~�X�Q�J�Cmߒ�����/֊ѭ��x����N�E]��@�N��z�l}��R�9.E�K����O���$�m�
q�I���T�}J��J������@,)��R�.�[&vq ��V�ðbp|��EK�r5Vr�9��}p���G�dQ磌þlx��C�A�
P��+/��G2_�dXX�'����w� %��S�F�S��#�3O�~��za[;A�؛��.�6��P��َ�{��y�Of 8�&���EO�_��L͈fM�/�N��l�UA��8���b��mI�Cᄾ����r���q���S��.4�&�l76�;�4y4�E
%' g�C�� �����nBR}%A���ˎC�T��-�7<Tq�|�L"��?Τ�.?RXW��*:QQ(q��O��&��-{Ќ�&W�h��̃�F$��}�K��W��l!�P����$�2�ܡ��#�ϰ�������G��Qf� ZI�~
IK�=�(_������
v�6%�a��(?�:�I�-&,5u���l�K�tI�U`���Owp�|�NK�i�M���a&,���l}��^�<Nɭӽ,+�ƹ'/,FK�M>��\z7Əc�p�taܸ�VP&�B�OWZ{'{a|#�D�չqC~�<��޷s���� �.{9���T�Y���J�!r5'm�����ȥ9.��XhN�1	x���g}W���/>ICii���'8ܵ�<B��i������v�:��xp ��x���1������a�m:f�v)BEB���{|��O�	c�~lJL�?G��9��^��<�R`���k_aL'ka��t)1�Ȅ�%���8���`D�ŠԷ��\�I�9R�	ժ�񬙮�\�jU�*w�$ٰ�QUޜ�ո�F��}�$g3��>8ף}��V�4K�Kes��'=^�*�T[p�����Q�I�Ӥ�e!�S=J�`���50�=L�`��$j��7V�)He�1�KM>F�>2+�9<���.�c�v�� ʁZq|\��[[�n.�����%QQs��\�N�M��QKK"��"�r�'��������NL��Y��^���x�;���I���a��*���Iyff���uM!Tg�ew�G։�§#���M"������ �QW��)~�\N��q�Z��9խ�?9n
����ɾx1��S{G_S @+]�X����`��Y�h!q
���C���^�D�.}_�p�#G2�]aTU�h�i�l�������'��["c���3f[s�=_���4����N�����[h��T,��f �4��s=��r.�fIZ�:��~\������C����~I9�^��N�^��xP��q�ظ]��Ա�L(8q[S��y��Pw�i�)������r�w#dS\����oB�>4�'7E�$gO�o�y�dZ�}�s��m�\m2)��7�;Mɻ������7_8騠��>	�C�І#��wh?�Qv>mu���^\�#�*�������Ċ_P.yqݳ� &곟A/+����ؕ`�uX�������d�B�~�1�dV��c�}rV�.}{��.`|x��(+Ro{�
�\~��^9ldW�Ə�"��|��n��M������*U�|,���ۊ$N��9��*,{������`��4�V!�c՗��4���_�5��Yu��\�1k�\�7�i"@�[]�n3&_W��5�i��2��`͚���\�^��
\�]){2n~Y����MW\���NNsH��S��f�\yŵ_���n�&�L����;y�,���2/.��u�{�k��c��`��`]B{p��VB}��=�esCo[. ��ql��'�!� $��l,&�Rř#sv���n��Y��#<�;F��]k��� *�z�i)�I��o�Y��`����#�̎N�|���t����E=8@����q��H(��Я���KǊGtƓ��<\�Sp�x�Kúi�$��=
%��4�(�� ��6VD�I��o�*�6L���Z��nmѭ�d6ޞF�!u��R��G�r:�Y�'{�B>�`"�W�Rḩ�>"�P�����p��h�����&,GTq��}F�s�< �<b�,o���14=k�o_r�<UI��!%©^�� �?�R�=�g˼�rp5ZӲ�]��Γ�!�U0cc}9��S�v���i�M�rTԲ#������;ibu�AS���Dx�����[J��d!�g�����e.��N}8v@ ���>�o�"�=� g:��{�&>��E���iݏj�^��^�t���)�jh�P􄉞�kx�O�1�8��Q�ޞIm][P��ƍV�	j+��I]>�eOYQ+�zajs]�x[$8sn�C� �؃{و�p������Z���cn�L&�(�5������~�cQ���kG�[b�g��}�T�{��/�.��ͥ���m�*ƺ�_}]C�k�.��G\�Y���kF7K���z�]j0v�T��Xr�̭�]����1G���-BF��b��Ԏ֎�~�Vr:���c���f� c"��Y����߮
��Y��������іvKn��:��[���䫚�h����wFY�}�ǟ�ӲF_�����4L�!�^&�����_����+�'��fWސ�]�ַ��4�B�A�����ʵ����|�k�ۧ�{z��=%���*2`*eS�|3c�>E�j1/���'l��X�^��1�o�o,z	���'V�m�֕N�/��� �����A���}YZ-輳��-tl���_�l�^�t�8�l|�d��c� 3	J�����U�������Fd-���ɗixDZ� ��m��RA#�R&v����a��~X�����.�D/���n~V32��?eU���(��2Q޴���]�>�9��j��>P_1��� �Aյ�I�[��ph�su�Z��1���Ҭ������"5�0p�d?u�<]
jɔ�:!i��GNqZ\z�:�6���������Kn�F�����J���p�����F$F��:j�8��em��0�b���+"�O+��IB����s;A���ݽ���9f~V�곊�2��F����A�D n5����y����7Uc<K����y{KY+9��Y<.��"�A����X)�9y�k ��:j���)�������:W�x�nU����Dl�h������NЈ��>=HӲ����N��y�s�����"�.��������km]D��#���9/TO�ƺ���F*�S78ؘ�^��2w���'�N�?	�υ�FR3C���)��O�z;�T�ׅ��,=�
�P�攜�;W�K�m�)������������ތK�i��$!���Ŭ�D��~�;6�q�,��뜺�U+�q�/S�]���E�x�8��/;~y$r��E��?I��}{�cX���Vea^0�	Rz�cS!�&�>��C�\����ڗ��u����~1�JSH�5�ܔu���0����v�XP��	r�-������/���uHNQ�yhaۍ�+V�bι��U�m7��NF��� ܝ��x��5B�o�s�Ӣܷ�! �G]�m�^\��'&�@Ta��p�?mE�8jQ��dH~�ɷc�4 �õZ�,B��4���5�Q)o�Ld1Y�l���������oKdk�.cJҚv����^Y+u�ԫa�l�X5��H(��
kƄBI�_�/��Y�����bAV����Co��/���6�0� B��2�:�n�䦮�>bjm/��op��P��v��1�(L�:�ݘۉ��Ұf�Q�d4Ã�k:q��ɞ%����Yx�]�j��]�`���tr!?w�E��Ԥ&zkmDʘ��p;>&�H'�^YFBi�{�&V�|K���(|��Q��߰O��e���PQ�C�6oԦ��]����|S�j���a������V�F��b�O�&���qE�r�B��"{�T�C޹�Q���Ԏ]�Ժ��e�R�����W�0���������ϔ�"I�<u��:ĺ�%���#>^��c�V����X���Y�2��ad��*���/��-������ �s`^��NB=q�o7�79ʽdH���"��v'�i���l�KI�e��2����MZ���?�P�]ߖk:9ř�X;��!o�p��X���nA�U���C�mR
7���I�~3��HU�E�����A_i��W&,��l�ߠ�o���lt�B��ia\�L���}&h��a�� �	���Oh��$D6�3�2ƴ�4��7�;�3�,��tu[��G+9����eZ�o�����>}��Ԓ�$�Տ��#����'�d���oK@o-������zi�����i+n���`K�Q�I�WGՃC�>�O�ڍL���Յ��	����8-�[obC�$��)�'�r���1ﯞ��2�Z�FՂ���uN+��y�x�Bi�nH&P�y�T,���m^Ndg���c�uXI�Ze 0�ҽ�5�Qsz��ɐ�8/o<!�h�*�I$z}#����"��[��С�b�F�5���b�M���\���K�O*�ª���d�r�n|�I�n�^���8ZZ�@7u��z�>��}�FR�,l����%�����Kd/P�fe��>��r�=i2@�Ε<���E�?b�m��#FLs2���؃Ͳ'uo��\#s�������O�Z�0��WY�Ǒ��k�f����4�u6�����gŰ��ˆ�tP�O�P�U13�D3���/Oz�-�Ӻ��.��[��B�L5b�.�7'X|!�V�����j/}fU��9�;��# �3�\�c���3.��+�����q�M���m��:x��e�xn�;��r�hN��o΢��4"�ն�`wґJ�o~�Mp[�C��U�8@w�Y��a+��w�����s0����%�e�8Z1,���V��w?#��G*�Q|}�������9BJ`�I[]���a�c 3��u)���*�`�h
�e�W���Q��iսu�权�z%��]ڋ�a6N ��˿��2g+��,]����Ue�wN�A7���疚�b�o�}X%�:��VeA���м��m	$�E�����!�nݐ�˔t��=���Z��F�艊�2ZT�-�(����wK���?ͧ>%�F�	�DHl�VSŌ�J^��Y:���;Bk}�-������ȥgY4�c����O
%�B�N�H���Ƹ|��#����e���t�%�wΆ1rUJκn;��}1�i��
�S�� F�EL1��"�qV���aA�I��!R3+���V�����	�^��x��=��&9�҈�8숺����<���C�v�)�e�'!2�m�R�'yt�˴����\Ѱ�0��\�U����\���A�����#@�V���68�M�l}�t����9k�Sp��*�u![RRjl	;y<a��g:�2䍤��fS��g���7I��}��FOՈl�$�r`���[lL/�}YzV=
�����[6���}>t�R��ޮm�^�)�-���s�}��H}_��gQ���H��T� Gr�b1���Y�	���u��9~7/�.)7��4}xH�-2�w�3�r�Z�[��d��9�zN���� :%���1`H���&;u.�MM�� ��6���3'_�<�Wl����H���ԧ}�J���\�`Yנ"%8��9񘼊f�c#�ӟ]�`n@��or����)j�l�J�e��>b[5��W�g03,.��q�eJ��D�ݢ��F���8�<h������������=������x��e�9���qEvr�г$B�����]�="���m{��G5Я�_0z�ܗ)�P'�%�g�Ǐ#�m)�c1ߠ�)����Df/�v'g��=��+���
O������4��6�9��]��^�������h7V��L�k����.Pu-�OGKZ-ސ�H~&�Nk����g�{��4�3�ubAGA'�K�++?������d}���g�4��|^*$柭W��@�Q�����񒼰\+�X���;S ��Æ�0#�C�����e�L|��[<����g�N"�"nQ<��_�3uhV�G7̲��cbl�s�_щ�7mV�Jd�5���]JtŠP��77���ƥ�E�f)��{�^�KF�iG 0`$G�9e�m:L��������a������޺���e�X�|�,zXc:�yԓ�a����#;�)�Y^��ۚd�q��*�����h�����kT������9Q�����M>��R[-�R��z�j��#$�Kg��9Bo�֬��lV��j���٧6����yiZ�7����o�㲊��y' g�펁��e=~��ٹ�QY�����r��r��!��oW�#$%ꠄ'��ѻ���+s���H��yA���_L!�����(��,Q�҃ �g.�>1���\���4�Gjǿ�]�&訆Y��,'�@5���+��{L������eX�SM���|�#C�����޼��^���qY�;S롐��R�ց�q[������

H~��.aR��c"Rc������t�Em����a�����li�����F�+ڱ���ϧ{��E�����Ẩ+I�}z.��Pl_���1(�V��k���5"C���1͔���=��?�?��V�uY޼ruy��c}B�`D�+i�^|o*��r��_��g*��K�lu����o���ij�4���ډ����񥓁Ub�kχf�M�Qc�7n�kͺ����T�j%FztH���]e�0L�j�
�|nV�G�n���g���YN)�Z��v/T��qFkz4^�_����s�/��w����XOPBo�Q�瞿�)�qtu����\+����D�R3�����];��f�7�$�u��O5�dfT�"��|�hp~71n�����CC"A}c���ƾ��(J�G	��ج��{wtZ �A�
�����NnB�Xe��b{��O���O����I�W�,r�i�AV�g��^9��������&�k
.蕧L�p���1��{}�K�E���~��P�P!k�_�g�lQ3�Å��=����(P�U����\��~�dt�3�CBd�ab���PɃ�ǯCW�C[� �k̞���Ip,\�U=kg���3��kТ�Kr{�!��1��|E�����v{���u����E���ϗ�GO���xgS	�H(na��#�d�?Ar�i:r�@���]�;��������pL����d���Wkq.-r��]�#�Ⱦ�����}�����1�FmZ_~3�|T�9���?(�"�Lr��v꓋��9�)�l&b�;����G��mo��0�Eu��G����_{M����i~zSm�x	8�������g��XSo��ٺ����uE��(�O�6�^5����v�$��!��FX<�]�x���+ χ��Z�n����1�5x9�E����,�z� F�Ÿ�e� _r����6��\�ƿm۵�:��528C�np��b�v�g��I�*����)�pKFv��t���
�7Э�����b���S�~��J�n�/���U��/�P�|e�� ?:�6d�Oɘ�o.��uvμ�W�4�"�$m}L�+��&�^q����Nܥ�2��'×�͠�q�$���2'A�r�l�^{���'�/���C����E؃�%�6�d~	���z���jZ��ߴ��,?��{~Y��{V�J}�Oq��э_ܴǹ�5x�ӳ����X!r��{���i�]���>����q[�6���'#Y�$0ť�-�^�Yyq=l�t�r0��K�Hu������׫���V2�ӝx�лc'��7cD�M%Y���1�aEu+:��+^e�WPv�X�[����UT.M<���::-Weg�����=�O�l��w�\�O��cf�W�	p'�7O�f���G��`t��?|3,��N����I��l�������ֽ"%ZO����O���X:r���"sB�=aVA��|Y�	;���'i�K��6[��rH]�������U�V�j�}�
���EV�j5MW��.#�琀��G�F�؅n6�?��aE�`�s`�P�^��Go��33%�R�fȷ�gH�������~7�K�m��)��}~=7
��M�ֈ��][�j��n֌��ņ2��Q���`���g�*$�|�)>��/�Y� �̷�����}��Amg�7�\�}�k�a=8]ۤ�XR�{l?c����˪9;[�����3��+�i�$�V�;�_!\Fi 	���^A���ޫ��G���}�{?�@�O��7�k][]|��;�3�j�V���p�T<�u[ٯ�"�nM�@�_�r��!��cN����`����`H��w��Z��k�^�L����:.������r񷺜�གྷ������ ����Z j�j��(�jJ�w�CQ?V���л`�fJ j��A���W����]1�E1��%"����x#<��iɽo��7����_�SS��Z��U+	�4�jh���k����{���<e/���|�HJ�O�)�cObe]����qJ�:�:���j7� �NS�>c�V���׻��i���z%RlM�FY���Q�20hG���܁�S&���I���No�C��[��e�%N�*�'�	����MM����4>�� T$P���ʶs���5<J�d��w��J
�-Z[B2_¾����Z�Rﻂ�m���}�,���?�1��(�K
�o�;\,"�|Fe�$�'z��Á�t5`���qo���:�`��QK�DW+��g2��?��0���(�� h�뗜*!C����愅%���Q6�$�P�a�#��&I. �C�.��̥J�ɣ���G����E��_�/a��KS-�G8�s���ɺ};to5���r�+�n�^�:2�s�W�6��l�L�wY���+�e�:���-e*����/T8�Yb� ڇ��Ǫ������g.`j�,�s8�Z�ĵc�74ir�'9M�F��v6�h
�*\Z��~-��c��W�jD�x��+���W��^�������m�^B�RYt{e��(Hhb�Vi�B_����$�X����Q��| �����W8Σ�P�p�����tjg��N0zV���&S�B��aY,|�J��v���#�$7p`>V��_P��fS���k�8o��>�0[��a�bR��N<��W}�)J�*[�Y��%��� �{c�m��)�7m�@+��7���,|��4r=Na���h�̼�*vwbC�Umc�	����ӏ�iE?���p�V��D��YD��P�a�+���n���i����[�q�uuX>��'- MR�>���u��>���N����j����fkM=_
�y� ~b���݋��Oܽ{�m�	%�.�Y��u=2��?�J�h�?	���ŦH{]�R�|^�!0�6zĨfp��α���u�5�&;�8Kof�����8�\W�`j?sN�3�X��?�?`"���W$�S1>�#2�׵�����9 л�"�F�U�/�Y�[[�P;��H��>n�j~js�P�p����N|�V��0�Ȇ����N���h&#�(Oِ2�`7\�g����x�Dp'z/D��#�����d���`K�m�N�%/�����pFg=PT	�	;�զ�٨X���Nn���M��kr���|86�o.���;�5T@N?�~��#5'x���/�����O�?�S�iX��&᳸�B��76�O�Ғ%ɟl��Q��s_
���,P�"�Z�dh�X��o�׾gk�>��� ��{��K4��孰�Ş�1d���\O^�P,.�Ɉ_�������O�K^�
��4O�83i�h�z��O7��⦦2M6ݚ	���hz�s/�r�m�#w>t<5��M�)��T_+&�ݏ��}�*ak�{Y�.�@�t�����g�^� a���2�1�şK��'�����U�0���ᢸj
�i����˦C�r�i�����|��cfw�ߝgm����3�o�<���l��3�_-Wf�jM�b$-dx=�W�4;r=Q��4��&�t��ş6�
E�?'W}�����s��v�}=p+%����ƍ�����@&�h��?�TA- �+[$��4��!�A�	�+���Ł�jմT>�x(����+���^ݠ�U�:���M��_�4�*��$�_֗��<��t�\����Ί�2ݹ�������߿����f��J�?{�R���_���,�0M~��)�?�x�߸Ѫ�>Y5�܄b�CI�L��SEI�:\�E.��}��5f��?��ix!}0}ڪ��Υk���d�j-�>t�i��ػ;w��|o~�s��/��w���N~su�s�Ud-tn��Oc`9������8x&_)��E��T ��@Ξ�9���֊���NW��PV���!xy���Iշg�ۡ�o�<> g�P�E�2:����޶��H���?GY?tl݅�v��!ο��#�@�����S8ߖ8���Ǒ'Ʋ����<��D������#dh��B8d��Kz�n�o"ŎA�n}v��A�w�l�	e��ҟ��פ"�n�3����Z9�n�9fN켄^���/(�.�8���Q��Wt��]��4����c"nQr+������*(J����WL�+Y�Hsث��I�ӽp6�FD؅��B4��)�mf|��H�w-S��H����׌��t%��z�"�\ ��Y|���>�ѐ��;d���"y4�H�j���.z"ބ�;^�ZE��ɵ��>�?��L���:sOo5m������ݵu��3=��C�������
i��˵�MV��$FL�{�uߗ	D��#�{��ga�L�.��RJ�e���.3�{C���8oH�Ϯ��lzY�:��O�8Q]q<�+1�������g���]Ɨ9��b�7��,k�=F:l��?��u��ﶏ& �^����?bt)��"�C�|���9����wP�֜���I`C��=Y��6&*U��ȮZ�E�/,"��R�\[Z�^�QO_[+�����i��C�晃P��_H!z���)�����y����t��*M�0{$A�����p^29-�G�sz��e�4��k�!��͍��R�]P�0
鈊��������.�����k+UI�NF��찗�L�S��t%��O<�O��t�i�Wچ�� ǋ��,���%e5���p!_]��/��ܽ~�	�ʜ��2��c�wx�����of�'Z|����o�	����:ꊫ��j Lf��eeC��8�6k~w��a{
�@�О�6��^`�L(9hgH�D�/J�x�~��Ү������Xh���=��ӑ�'WAO'���ʓ����8y#O�D���{6]��~8J�j�R�>K������
p���F����-�ʃ��ì��4�U�������"��g�?Ɯ�m�r�U�� u��|�[/X����d����Rppz��P�o5�S��!��ǻXT��<�Qّ�ֹ�&Z�g�}p�:8���AY�V�TK�&)K�Խv
�ss.3��ɔJ܊���(�"&�M�-J�W���Ix~J�?��~�M���li�	�s.0˯�a�ۤ�-��{MK��|�~Y�5���K8����;�Õ�qY���G]h&���>�0e���lK��%��.��i���{."m�K��ګ�y�@/�boO���� ��?;��o��>�t�����H�$ӥ�Adì���L����/���.ڐ|c#�B��"��������~��3$�+��M�B���N?}���^�F.�4���H��K�� 'LM��������0X�8z�/M�&�!v��Z�g���%�˚{�w�ؓ�b��3p�#	q;_�D�伵͗��~;
�n-w�����ْ����u��૶�1�_z�R���H,q�;N���
4>�Ar�P?of)yt�=L�P����nt��/Ŀ�_����l�įρe�Wް����̖�V5�\Ҟ4YxK���3����uo5Uj���"���{=�8l��9�u��h���u�K�╡ȼ��b�RerP�iWf�)v2�U�<U�u�@M+��n|IK��	YH����S*���5��%�����\Z<����(&l�=+�\.b��A����;_h�%j@���E/(m�2����Y.�5S̗Eʺ��L�����8d������6�Ҳ������R?�{����i�*��cz�P�ZX���twXn(����	d5����:��?�u��a�����}w���~ZS���5?aD@�<J>��3�^B�o@�W,������/1�� 0�UM?A	�)��i�2GVQ��jߍ�Ru���dl�~z}9���<j��k]��y-KV���+v������x��XS�ī[hZ�<�I;��oF�����_�=���MP=nqiK5FT ��,���1�-���au�{lqӗ/Ln�o��T�h�S�j$�|y�6�[S�xX��vz���դ�SD�<����P�v$�b�-��ں 5Ybb.��6�����lf]P��,8�x����c�
&("��M��"vF���2�O�X�w��I&�wv&�6��˨��_b�*Gkg)�\a�{�}�B7ې�`���ৣJ��$���x��Zvl�A>����h.7X���@�O,����o���s���(���M,d;��E��d_�U��'!��<�
���6y�I1N��º����19
�<�8�����'����&��V��g$E��@Q���}י�wG�&5�i��jd�1A�OA:�`��[��e?�yn��D�0x�����n��&�ZO�W[���a3��C�=���&�y��Fˈ�w�6,f�,j�!"��.գK[_{V�msR��S�U]�:�A�%�,#�!j��	��ڑf�Z��2 p��4G����>���"{=��H_pqý&l��*&��-h/��gd,O�w���+��e��ly[; ~�����S�H�Q@��seD�t3�V\,�ͭ��m?��n-�H��ʌ�}y�@\7
2��� gl��Y��9�)Lx�rĺ^��c�{%c�������C����jr���p�j�֥����ɡם�,���+��w]|�i�?��j�9� eo��m:�A�=�U��	����߯pH�1@�]jg���A������W����VP�ٟ� \{��%�=��u|�XV��8�18qo��s'Ywu�Qk��H����.$��lX��c*�l�ᴏ�&�ȍ
'�t������Y~Y��������6O�D�:5Ǟ�✁c����*�#�>�V���N��xV��?�pܬ���>��B}<bC��$�F�ʁ�?��Q�ʽ�[N�4�:w����>��B���f����9G8�OqP{{؈�@D�F�UR헻Wʀ~Ul�Dr7���F���9�$��0��#�%��nnm���b؎L@���$�(���5{�Y�������$�66=��]�t2��7��q�������?>櫋�R��a� �f�|#hs���N�o?�Y�sc�\XaN�-ϰ�t8d�����^�%nP�d138�W�HLcp 4�@�ۋS�qC{��/���k��V)��ڦ�� �E�ъg\j�j&�T\D<!��oc6T���@&j�q
�d���nD<�OeUƈ�K��?��������X+�p�Z�i�Im�I���͢�њM�u����K��%�&r�Ŕ����E��i!��x$����u�<���gzP�U��mO�
j���[�E^C�C򽭫�Yd� ~�G��+9hV>57��n3�����G�G6��z�A�W�0�e���۟{��~ǧ�uRdx�������M}Cle����έj2}�����q�T�'��νI"L5AA�ouҸe���X*���N.Y�ypBj����2��GG���mΉN���/z����@n���T7� ���1Ԫ��4�*
p�Ch&�>!��42�����J�6\�����Cw�{ּ�hS�/o"#�/V$Nڼ%�wJ7+������E�3� �~N��WwW�WVR{}�&PX#��'�q��b���T��,�V���U�4���M�xx�JF^�nb�t��=��=KĊ������r�L��oh���O�c���m���u�D�<�I~�$����t3�����p��/$	�vʜ<ƈV{���~7:V ]hP�Ԩ�`VL+9g��.5���/����u�ϥ	����E@;F�#�0��}�w;- 4F���KX֏O��B�fJn�m�ae�şO�ȍ��l_-��\o�J+�n��n{zܑ�k�n��#�W��H��1��:�?���"Z_ͻn�����P �zo�|W�Ŕ��ł�e~Y��@NKkx�]�S4<y��p��X�OA�w^}��U %"h���) �cCJ�uk�˩m��0[��y:B���B�E��ͨ��o�qDl�e�������$�A��3Ka�O�Ƅy��?7����A��7�P>����b�ŁW&W�0�ߘ�犬�h:��]��
�]C<��R��:�ܛ��<��Ϝ|�$�KE,`7��N��/:��#� j���j:zo
4�t�~�˽����JX:3��o)ڇ0��coO�����nɮ������+&�j:6"-�M=o*�LJ"T����f�U̍r�ޕ��(��,�A(P�-�#/L���|t��)�"6`_)p�^����)p�fj,��S�N�^�EI�ۇTq��CʂG!D��l�۔�Zy�˂���#�`m��"�S��IcI�k`EHJ��̓��=�����,��Z��9<�t��`��,�^6��)3(��������	��l5j��2y�A_̓T��K���&»�:�T��t!Wŏj�{�e�A�#Z����v�(;mE��sR�C��F�>��oK=���AH���Fv7��@]���;��o&cubO��6fEA�/�����*����$�yEY��uj�cɇ��!�"��"�+��{�A'x�eY�Y�3��#���U3w�L}���엙���Y��ԊK�N���m��>�?W�TBK��7{��jiiB>%�>�_��;Cs3c������G�ʞU`(cO��;�:tK+Ti�/�ϖ{�<��r�m��[�d����b�YL�����A�uw�֮H�����rbrR�K�\?��ca��3�B����o�Nzs���߾@�i>P���>w*@t@�#�Z#۔�����SҰ���R�_���U¯�vE:��p���Xb�ߥV{6@:�g���i����fn�m�j��XG�r7v���թ�O��5��9&��]�	
�2s�"���<�����Du���
���t��5�|;��OFŮ�/Z�ĴpD���a�{v�ݖ�L��S�	�ה�Ψb�@�K�3h���[��>FR�,�����W
�j��G{�����,\{;���拭����K�Ys��ւ����#ec�\C�Y�$`Q��4�}���KțU�ԧ�v̾<J������ZY��Ye�X�"W�.t��h_2��F�>e� ��0\�#�y�8�(��u�p8j���Ԡ�B�Xt&�EN�	z����顣b���K�s/R���u�LR��Iw9��ρ��lիt�<�J���g.:�yV�gL����'?>Uۥc��2V*���3H�7w�ʉF��e��q�z���f����^�U�28�V���J�����*��\ؘ߫��M�������$?I����U�|��d��$��⁩t����>s�����M��H�EIa������[�Oj����ZcUT2��/�l��B #�p�v�����Ȯ�.��GBq��� A&f�#�W��YS%͔Y�L�\�+p���V���(S�'�ə�a;� 
*�i��2�����_*iA	5Ŝ"�\R*/���0��s%E���q�^`��./s	^~�UGE�k�c�Yq�^���8��8Z�7/�r��i8�� �пt�{C;R��>��,ԉ��e�aWK�w1�
�۩�7�b���˝�杜��-tY)����IYj��R1A{�|w:j���b ୞>�@�%s�hݵ��-��#�M@
�6ԵL���;%���kxD��Z"Wc/��ho�V��m�x�O��F����u�V||��M_�����r�#wrC4G;�l�,!~�f\��{/Q<R�)�R s���"���G�Xd� o��x�`*�����J˃:6��u��icϿ�d>�D	T��{��{�+~�����N+�57���V��e65	�r��J?�?��;��&���"*"JU��Ҥ�h" ]@@E:�ׄ"6�7�M�t�B	��P�HBo	$��@B���=�绮��������7s�޻nc�����,z9oT��L�yZ\����/I��+�X�B�y��G+lS��
�jo�&�PV���[O۱�xM�և�W�7xtg��5�(g�=BT��ɲ�s�՛�G���C�P����/��������;]�.
�� ����qng�0ڥdɁ/(�r��|s��	��d���b%EE� ��:���{:�Z<�;hv+8���ui/�b�%6����R��Cs��OMpZ���9]��C�b�wZ.���0��S�9*��x����΢<��M�B,��*h�C߇n�+���]]�?3da*q��T��9����0���6�A���\}�P1_\�ёK����#�k���2���6J�AVU���ދ���K�\��aL`ƈ��N���s�I0]�@� ����-W��o1󟆡���H�ֽ/���97�ծ�������6pA��)�ݷߜ��u���Ǩ0��D�t�'m�bl���W'��D�W��A�����s��� �W������x��m�����nE�û����Z���,�\�?N)������rճO7�=���IBm����W#S��������]\;��OƄ�/Q�(�����%A�.���>�������wX�1�(�����P��u��Y~��&�]2��:E\Z��w\�O`���Ѯ�톊ruL����
����k�wA[���K�1K����U��x;���g�Dx�i#p�$�8c��CX��n����;&���h>����Y6l%���%[����N�~�}�a����-&���R?�v퀯��>@������yF��6-�ʢ���g0��� @���~��Z�����~?��h�2°H�2�b���I�.�x̑j�E��k%;���2�M�6.��O�W�6����|�OH.����PW�sp^,�K��b�#�&�[���v�1\��$�j����C��R$�����y��V�2��_��ji9؀��(ϴ���Φ���@�\a���R��G��\��9b�'m�2��З�}g﮾�(��?�?���;�Цf�$;� ��fc���?�d����o��̀�]	�Vʸ.f�s�iLڼo)�*���?{t�� f�*��`��Ѡ��]��X�Hu0yS�CT�Ry6�H��.�~I��.��ؓp�~������B�!����w�*��~,&J�y96 HH��ݵ����*/��&O��aY�S��O��n�02RV�,
h-_g��o(�Ze9=�hW�(�ٸ�.�Tۮ(s���ӽ~�T��u?����ix*�I�ׂ�I�������� Ne�U�Y���ʫ�Ѷ�'��}�sH�N�5����>Q��j�$��V��q�+��}��p4�T��8�xLx��6�*c{��K�RHļ�ܲޯ���X}��@�8�^2W���P[��牢���9��Ak�ǻhK�\咚Ԭ}�ǳk%E7��X>p6"��z�qgΉr������o�y���E|�8�	���e�T���s�)^������2��� ��M���w�&[�a���=ϸ�b⸷����/W��&L������Gu������s�%�M Dj1N��jNw�KZhZ�?��K�p�k�1<,��� �"��<���29�����5wG�����g�K����.��?;NL�T�&����Qk���_�iy���9�Q_o�(]��ll�����?�D`������"W�J`��Y��mG�dy��k�#���Ȩ;�>�I�91�N�E����xb����x��yoT��5^չN��|x�V�66���J���������DbT$$��).�_��[�a��~^���*�X|૘ ��ɡ]�GZ:W_�3v��z���ΜCn�t&zMHE�"~�j���a�/��zse��Z.���Jܷi����>J��z4�
��k�w$�k)
W�F��܄����o�m�o-��b���S��t���JK3W���
�z�S�W��S��a"IJ�r��+��ǒ���0� �$�m,�U�ލ�]�Ռw��[F��m�����ۛ2v�w4=�<��O�
]4���%=zF�y��-[����������#$ҫ�^h29@��=���۳7�<.�Ҍ�����(5�9��v`�zb���y����	��
�����4��fW�
4����Kxl��"]�7���+��o��9����	ĵ�Ct0��MQ
���k�沕͖y37���I�<�F��1>Cs�M���q1Q��H^6П���2E�-�8G�ef�9d���/�A�Ͻv�ہ�=gI�������t��I���?(�s�2� ���E��Z�+3�\�Ф�e�uθc�K����~���i��\|5ǎq�����_��(�R�Ka'4r�6_s<��{1*-}n_FF������7���74���	��:��iw����D��Nb�]\�����p]S�Tnpp���E���W�����ij3a�-���~�<�0�s�σ�]��ӛ6Z���W|_3p���d��{����Mjf獼����klG�%Q)�'�@����w��+��7�K��|=L�1��R��k-v�˿߯)o��i�R�������6�ˌp$h	\�=ZQ>Z�{\�ҟ>�c��E�羭�ϣ�o��bN)G/�Às�0��cD�`����V�	e!���	�ָ��2owƄ����l���O�lzDL}Q����^�
G�iq�g��
nͭ	�;�U������3�i+�� ��1�����]��p�;[�j��J��}?�	�=M�Wh��%�02��nէo�������mW��Y
h6θ�t/8�]��|�^�F�	3�<y6�{a��[�@��P�t�Ux�0eb"����'F@3i-d-���,��x���+��h(�6z
�1l+yӹRv|�U;uk?hE%JOU��*Z��V4q�h����������Ap����M髬��.h��B��&+Q�"�;Hqv�q��$[9,ؙE�������xK�5��x ����d�\M2���*�B:�'�E\��_��l��H-l������j%6��eѸ�BF��Z\2��m�f��T�<̡,�ƫ?�P���V�����Uܜ��9���c_�;�P��G+짼��*�7����5�������Dx2����J���M��.��X&�n%�Z����x�!�a
/V��}��Z�K��(~�Ь��'g9dŕ�S��� ��}�SyD,��`3>���*�YJ�DG��o-sM���p� Rn����������~n*!�[�������a�9��cZ�N������I���9f6wp�L= zr���������n�B�2�lV��	� �9��>�e6�Vo�s�߮|3���w\Xl5٭.>���B}������2y%{+����x���^��2��T��Y]���W�զ}�u��_>��oo�8�ȃ����^I��<{V��2NQ+E�6����^n;�G0%︬��ͤLߘ�e��|���R�8�?�f��C�"��sai���$�u���}8�3�˥޺��d��6�o����~�U߲M�
�O�Q�v3pu`�s���������|<+��S��L� ��w~�����jϦQ�ㅻt��)���hR�
J�Rv�å���m9-q������ԎƵ���#0b��_�
������~h4�Rvs��s�LP����!ؑs2ؾL�(^�/j5^�����|(���y�H��.:/��R�Y�|����C��~88t����&���=�ցb�����ԩRo27����mw;����fa*���~�����J(E|�Ѵ��(�����!�T=�����6f&t�����B��}�O���
�����T���!����0�po=0����J�Q��{{��^�qU��a_vn�2�(��׸�^H(��k�}���( ���Z�V:z`��Ķ8Z�Jヤ��.�9催Z��6uȴђ9W��Ϳ�=q�y��h1��U�  a���C^��z���3�PS`�]����XV�Fdid����c�b��h��S7�B��ս��T8~~?�n��!w��g���p]���D̅�6��G�!V	�����M|��,+�* �<8blsE3�م6i�2.�i^���2��ښz�sS��/.��ѽߪ؊�py��G���޼�L�x.FSj�^翑�9�^�c9VՆ���ۭy�]����|�'/����m�]���5����RN>#.��O���R�5h��J�O����9��dh����}<C�)�j���-6��Vi"?C���V?}��"
HZ�U��˅�58F#+c��Rg�9����q���,�0H�C1�t������Ʉ��h�
��'(nO�%��q�UX�����H���{����׷���Ȩ&N2��'al�X̍q��a�5���k��&1�p9m�[��ᯐ�^�����a���M��o�d��`�s$�����u�ߓV+��,��~XJj^�/��K��=��s�ϝ�Wg�,����C�%F`ὭdVP*�d�+�\�����<��}c>��gyt���4�!b�ț�E]͛����'�T����Y̚;���n�p�{�F|�ɊN��wT��o/XQ�\� ���'��ɁBrݩ���9���\�����-{�:�3y�*���ĺ?�adZ�|)��Y������B+�� s-u�y4ӁaAfJ��[���A���fv�k恤)d��@Q�~"h/��[
�������[��i��y����K�%����*;?#��ݱ�'�g7�}�Ô������/�@�?=]Pc�
�MYB偃�衟0�|�q(�SFXt���)m�i�%F��^����AOi����O8����߃��	�8��$>]193��h_���B�3H|��R�~�+�=�S���̜}�:&t�+0^B޽�J�����W>B��U��.�S/��><�I�Ο��H�9=�'����h6���`��1gQ�з��J$���㙮�����N(���r�`m���ܟ��� \��q��+��2�i)L���Tj���G���RMlV���	�������`�C���aeK��;�e���:���H���E=�u?�p@�����J<"�%+���Z�1s�r5������E����iN[oؚW����<��x�L���Cq�`'W�����U��O��Q'o�T�e�f ���H;e��R��=\u�B;�	=3e~������n�"{�h{���H�����׺���Ƞ�K�X���\Y��+��q˹��ֆ�v����sQc���D5"���B@������,�2�,8kN�%��e�ty�/?/z��4z�ӛW{�0Y��031�dհ���@�1b�5��[�M�ZfN�@j1 x&1I vv��E�kq��"���j`��Ii�E�A
%xG�A���ۃ���3Iϩ�ٟ>�;Ȗ�#�wc�'��4��k�y�}񌀑�<u�aMda�LX(� �?tq���u��Ô�Gj�u2)�fW�؍i���P<�������[��l߻�D�jEy*n���3@/J��j\I�'iJ]ϓ�F��zv��M�ES�4�/X{q�]��l\SS���G�0���ź�#�>DF�J%����E�]��C���n5������i��{8H�\lu�����wE?<п�|�b<�3_�K�a^^G�������hꏶ��	.BOðO�7X?;����s��c+�h���fA����彥X����{�5��	�+��m;!�Y��3�b��W�wt���o=�՟�f�}`���x7�R��&o=0��Ԑ��[��$M ��[�9��~j��"*�D��8[�t�^�8ob��~����T�z�K������QD�N �r��ŭ�?��A�ࠛZO��]���S*W��="2�ue~��T�G5|$s���U;9k+~[���ٯ�[D� �<K�sۅB+ȋ^/q�&?g�V����2�M��R�Gc-X�<���?f1�R��Y�S��8�5��.�
	6��ˣ�E�%�����ߡ�1�w���{�_$醼�J◖�ȯI&�T��ep�Wo>[��b!�|e1y������� ��,�2n ��`oN�E��%�$/�G��G��7���:c�M	}2���v4)��髛e�@?�a��}/�=<���cؠi0T�R]���X٢��λ����ja�Hн&���Q4�����Ac�$Đ���P�.-%[W� ���=�D�M�����Zm��_3��Z������DR��Ԣ$�G�1s�����p�t���]w��~0Q:�9��8�h��e|���6Z�|1�!��wl�M����;A_Ը��[�)(|Y^~#�-��1���~g� R�V7� 0kv{��ܪ'=vzܵu�Ubmo���T~����Di��2:���i�>aԢ�$\hހ�?p��c�����n�z���A����V��a����oL�
��	�>i��:���T��7Em0`֒�kr��)u��G��z�	�L��Ӂ�f_����0E�V���X��J|5tޥ�����ܪVTXt��
{�v�SB{�O��<���C�.p�i�#�F
�[P�Y��;dE�뽱B������PN��9�����u���(A^�p���xQ@���FUB�]���6G��v����^1�&o���l��ZW���2� !�-�����0ʫ�v{G,讇��{��7�8�n�DI�^໑���aa��Ëp���|��Y+�P�8��(׵�2��3���K���3_�0�s��j�D��3Р�M���X�"݉��N���}��I�
KR{uFf��>r:�����u�_��y�����d-��[sb�ʹ��������J�^���U�,T��3k}����B0��]F�'g/���8
��j7���x<@.�v~̠ۘ�3M(F�� �Ol1�v�,o�9��NC�PT�kƮ%�
�����$��-��K���W�JI��{Ɂ��u��T�]N��z��Y����hRb�;�\ )�M*�}w��>��2� �p��]z���:��F�g�.���� �mq�?�^���8<��sŭ���p��ҁ���P�ƅ�%�����II�>����<`�E���T��O�p}/����';qǔ���1���=�2��C(����9���C�o/]je�S��V�Pcc3k��~#�x��K�*|`<>��̖-Ԟՙ��Gf#'�	L��u^��q����1e�T�D��in���2�w��w;���w025���M4����[N*�b���H���N�}���W�g6u�������i���QQq�T2y�i�����Jŏ�a�^K1�(�DH��S`8���%}�G��.7x����{��� ,�H-.V '�J�Zr"��gG���G��k���dL��f~ޓV��B�����4v�������	[�=�%�}y�hr��ً�'�=T�XB�OP��Q��3��'y^?�&�u���)r�����J/����b��v��Jj����{����Ԋ"ݭX�VL�N^�Vqsc'�� �hX�g��5���c�܎"<�
��{�}�r����v-�����\����=��^��y��t@��v�*w����/����z��76��n��ۘ��������M0~�2����t�o��͐$�}8n4yE������io���]�^$y�7���"�&��.�j�h&�OXb��Tox����3=�M�qj>#���{�M��-��7�:Ν�ww�H����ё�� {Us�Otn��ѳ��*z/C��&�Y)?���%K0@�_	Z۱���]���)���`Z��o���dQ��ƺ������'Y2��NO�<!D(($W�!,��ek�"}Yca��C\��\Dh
R#	�Zr��}�J��5���>��|���$s��j��n�z�����km}Y?0�K����sPs<JD5�d+C'�����'P��k�M��	Nl�����SEepyA��&�x��3�����|�1 �l71x�@+G�˼d@ps���zSBe���'O���QZ��MK��{�#��	/~WFg��<��H���%����T|�LU���"�5C���x���2�S���J�'�-8�W�8�6�v�>Gt]j>��PJpoB99PG��9�*.���<�V��	��@��\}ܹ�U�k��Ǜ�柙 �1+����[2������{'�Q��wʬ��/_9�M�w����?'�Ը��W_3�4�P�ٴ12��܁�e��\���`����=�0�99�4\g>�8��Q���X0���4��S�O�T�ܜ����@��.��V�H�ugV�OT�wO~�"O�X�]��P��J�"�'�C��Ŋ��/���g�I���YG�A��� 
������Q8h���S.���񷑽�Št`�v�'W��k��g�A�7���K�טҼun^�U�˞�ףּ�{��7�G�5�*�.<�>DY��Y�x��I�)�ђ��5v�~m���P>���oY���@_��;t���$Ez+'&�r��0�9L�f�@Lq�6U��V�{!��������G:ܲ�$m���w���%_4��l�8y$?B����k{n��C�+`[c�{�;+����j/u���
���TU��ɾ���W��w����"���5�}�#u.���f���cIr���g*)T\LV��ݓM-qn���j}K`vd��:;�i�N����x������65��:DWy���`�)#�^�+��:��b�N�@�r2;��%��T�����x��O2�d�����
�2A�gVG�c�h�5����� �zh�� b@Q����}��;���vO�v��4B��`�k�B�4c�i2/�FZL���,�]����m�&&�j��}}��ՍJY���B��^��0^��j��Wf��C�Pb��: ��f�
ܺ�,Q7��aC$	|��i�.������*ԩ< )�����ؒ`�X��S�껒�_~�k^7c� ���B��ٜ� ٥҇�a�4�N ��Tw�8Q�ƥ^�
~,�U������m
�f�g�%���}����g`S^Ql�F���H\���8ʹ�5��Ї#Yr�^Op�D�J�{�E�m�~<�0K���Wa6�pO���u_W�>u�x-N�r�Ӗ�NܼE��,���ߵ=ta.e�q��!�O����@�qG2�蹮RDu��A+�x��\1ƛ���g68�n�H�:\�����%��<+k��=����4-KQ�=Δ$�r�K��x�Q-y�p+(Hp��@]�eMO���Tn)"�0����z�F��7n~��ly:�H`W<������o�FE6!��M&��\���0���F:�rq�6���jRO�hl������@�k�Oٓ�R���ۙ�s�^�e��.�~(퓽R�&����p;h&��D�wU�TX0�e���.���>�[�ǳ5sw��%Ȳm.w�lFG��}nQl-���+^ס�������N��H�oj&F�yӟ�� � �S�3{��d�1���4e�����gw;Q��n5��}�!7��X2��b:(��cј�߷�[���L;:�V�a?aXx�̼a���j����������������|%�`��%���,��քK0��H�P��o�6��R�`2��A�7�����k�>��V�P�������-��-g����q��v�����4���~�i�Ⱥ,�Mp���O�� �(�8<��e�鍏gn�>B�Jt媠��*��z�vC'Z��|VJ���
��TX�CIR�i�V o1ֺ2q�i�.�Bе��������>Z�ty�H���U�|(5��pQ�L�� �SB����~���[��I�j���������"u~x��DX��@����/Z	�ө�(+��we%di�"�B�Vd 5���A���&����k|'������Q�9�5�Lf"�&�V<�&�e�b��>�]��$%&�$�!Z��^Z��/�2婝��܁��7��� �yC�G��	~�����}���鵮�V�-��^�s��Z�)~�vlx��+����x�=so��l�A-?�^�{t^	�^���~�S�^�=O48�㙯n,�ĸ}�Fa/7lkd�ǡ�������Q��#.M3��B�e�2<�T�uRW^E��FJ��7���ۦ��D��!8�Ǭ��M�i,��	:�b_��q��ͅ�%�[ߵO�L7]=VW7�h�6ϪK�فis����ָJ�����J!e:DC@������,�<բ�D��)��Fo���k��>��|+�{T��Wf|�Vv޽��d՗�(�{�����pGGRg�L���GAD��]gq�Z/�c+�Y�b��ͣ����ۀ���Wz((�2Ի�2�am��i���S/�e�$
�@�K�w35v�,hY��1Q|'v�x{�T��wPQ$[��Y�Ak��N5�&�Q�:�ׁK�O�P��D(���%�������eFK�"�7S�A�&�
?XSn@,�����e���3�[�Qysff��5�K��jg���q胜v�P�=r��_.1#�����Qҍ��2��t�Q�|�iRB��QŉLv@tB�w��_�Zm�@�'f΁����B4���SR�O畽q�i�^�yb�c�`npII���N��w�P�Pޠ~L��+��H1�E�o2'6�Wo���$�F����	�N�!� ���kg�F�η�[ ������[�2+1�#9m��K�6ǻ��6�)ms��/�t���*W�|������Jb�6��f��Qb����PN�ʸ�u��o�Q����439W�ļD@`�b��:����W��`m�V4���*+M���m|�+�y����m�pz���s��Rw����ɀ�ۖ�Kir��(�L�a�x�{�����'�j=�:%��?8�@�p�ho{�BU��yv^��弴Q�`���)��e��s�;�XmLo[�~v`����v��r�ڛ��zu�1f���y�XQP>_ao��cE��Ta'x��²��pdO���Q��%\�']h�iƪ�Qj}|cb]����} b9��'�� ��������sMTjl���H�~��С���$b�$���̱½��O=h��'�q�����^��J+,�8dڝ����K!���U�d\��#y�ˍMq��K/���y����O7�ݚ�eg���Bd�N����+ƕ��
��j��6G�)��_0��^���������pޏ���s�.Gmo��q��
�����/G���A��.�i��w*Z��k^�o�Qưf�SeY��H�A(�Ӝ�0����>mf4�ذ��.��Y�դ�e%͛���]���f��]�dc�_cM?|�~�b�2mhG�?T�^��������ˡ{�̽[t��*�Y.X�&z/&]5�~�}*��� ׎�Ï2��Uw�Ռ��i*�F��� �5s�ƍhڝ����J_'{��V,�S����<��bS�诽��F=w�b�K��ѽy~-�ڿ00���Q5'���I�g�zM�����������[OZ&%��i47H�%ϴ��-�s����,f�a��J�-���X�v��J�ϥ3�d��l��N����๗���m@��t�zG�̪�Wz�?^��<��3�o?]?�@p�vj�w��4�P��(��G�a0���[1CRe\�F���O�Q�!8ֆ�y����F�B:�#|v����е�h�E�/Rz)���m&�2��0��#��VQf�p��" �(<�(љ�X�^0/������x��E���D%k���E˘Sv�������*=IC�/��|�����s<�R@C*	�0���.�Q��jR�JS�V�o3�K�R�{0�䈡�gEw�ꇼ(΄��c���!g���1x�JAKݐLL�f-��ř��,��$@:��P0��P�U�c!�U��ʺs���K����ì��񂉟oRMc�������ݸ�r?e�gx)��\�2�� ��x|c>I/����k�l�z��p�ə���U�l�s�t�������!���s�fko�0<G��[ռ����?ϝ�*l\����Ȅ{���άɗ���H/�)ɻ�N���U�h�7�'R�*��d;�>�qA-c2�%{�H�(���U�L�oL��?F-b�l�@r̠H�D��8/%�pn7/��G>�7(���S���=���d�EC@���a�j�J�j�xW~A���b�g����b�ֱs�3i���k��1Q�%T/�m�M��j�.�vC�j���׽*����g�d�C�~y�t����P!gK	�ӗ�#���X�ʟ�u�J�1@ۺ���iJe���u��_pyo����'�&7�Z<Q�Bi���{��NYЊх_Yq�&�5�YY��x�D;:��-W*��G�R"!g��2Z�J�z7�Y]�[�|������b;��{�>�%���t+�V+���d�T���`偪��cg�+�+DP�*��8���h�7w�!	d'�"�3���+SL�V �]����A-c:�h�DmqP���@�&�mlg`�=2K�6�Js�4�䉑rN���!݃���l����NxC���6�6��=�����̼��Yy{8ƥE���o�w�U��M%m���Ɇ�8=e��w��>h5H����I�����Ҋ���
갫��gTky���\}����G6�!M������gD�P�V�{��y���������z���[�/��Y�ܨ�}�I����'��12�i�|���=�!%��Ӈ)��^�|����M�_���ɾã����e J��"�X[<�<�]{H�����,��Ї0��{��f3]�J@�!�	��ԍ�/�{�W���M|������>�ݴ� �6��X��`�&��FL�u3R��v�=B�k�S7=�4��F/��M,����ǐ'EL:�z��MY�f�n��I?uQ��*�u
�;م3�< �@�"e(<�&�/_nm	��h��=�H�0�Jn�-�:��/�`"m�	h=��y��N��tp�M"m�;:z���^MwY����d�}|���1��w�f���{�(1�ﻎ�P���L���"e1e�Ѷ��c,w�	c`�ؒ����]���'�l����s���J��=Mϕfv#�rZkwDxs�������۳���l#P�e�=�	�A\�a�HO���|Ľ�@&�>�D�E�g�7X[�z�̄���;P���Fr��ш�� }m���3���9Cj�QWʚ���֨��_��~ǷЗ� 3U7� y�s��]9�y��n�O��ma�߫RH�ڔi���o9G��W�\s��@.�U�C��&VP�/+A����LxL0�mB��Q�L���������R��KG�bF�.�΁>;�p"�PZ�T��6�1�z���b�X}v���tb�/�%b�nrO�f�;-23��5T�٧�L֗� �|U����K��ֽ����M|x^B#{~��q3�� ���z�o���5j$,�`{z�9�~*C�!\1jѫ�'�_U��!����Č�GJ�{O�,6?/����� e���*{A���{�&'��v �*�FĐǾ��m�kIᇮ�(����^�tF�\
��M)��|w� K�(?u��?+�,8G��y�ͩ6o3��R��Q�sG�s����v�@�M<��<^c�q1,%+�V���qk(����Q������>{��=�z�uOي�d1E�RUe�;���XA��V�'��o坫���?ި�|�x��%�szzP�x�����0%���4��R�y����C/��kg��K�mfm��Fw(��닜�y�mőR!����$��#�RE�%�N۩<��I&�]j��K��|��v���z9������ *���k�R��L���Tz��@��R�0���3w�����h���B�x�8��24������3k��kI&��ĳ"��,�`�.3~���T( ��Tc���hպG����/lXFe?+B)A��2�Br����e��НNݛ:~tM��ԟ��j�/~1�)Ȝ��ZC"X+���j�cZ�YҢzi�I�Xq�B.�8�6a����תԉ�V:p�7v�� �d� ���*��l�=T8���P��J�Ba�AG�`6ҙ�5�lb$%m�q�^���%�O��]����&���e�k�Kd��ݷ`v�losˬ``}�Ds���V�hDY��x�ӛ���:��}��&Iy;2��8������c�wd{c�-��:>�0����K�V��7�С�p�dqI��D�C��97�(nw�C@��S'+-V���]�t�˩'+3c�u�|e��\Jen�斉V���n��jb6���rX �T{"2۲�)�魦�\�M�0) ���7�a�Ҧ]��;x��݌pv���]��	�
Û���G��W�?�D�[Fq�ޘ"���{|8��?���y��Rƪ��Vm;>VO��2�|蹁�Ӓ�a_�LD*)-PH���y�֪�ܚ�2>w3},E���̽<�_�v8��Ӫ�^�~\�&ei�����ͳ� �x���EvD��kT��<V̅]tx�����k`��Kc�[g��ǥ��=������3Z���r�Ik�Z4�ғV瞇���ب�])e�R�a�2ؤn%vaU*,UA�۴6i�!�����J���Le��8���A&�<[4.m.;�؂���������K_s5��]��ɜ8��R�-F#�ջ�ߣZ$]��C��v�?�`��I������Ɏ�+�-�64�q���\���WL�b��M8���R��W���@�@�\���[����q�F�V���V�B�%N}C̲�ֳ����g^������^j_}�	.�"z��J]���6�\�,#�f�A��8�-��Q��¬���ew���D{�>r��.��f��t�^�f�����8���Ϋ,��@ɷV���rO�K�����v��]W�[W����hk�{g�m�������) ���a��ʬ�Z�.10��B� xM֤[�"N)�y�]?0Q;��V���@�|��,v�&��L/b��A>̚�"Ƴ2�'�Y/^k;ٔ��m�4�;c|���V��ŵ&6�]8��@3����X�^�E�w^�׏Q��f��h0|�a!E��<V���Q����P5;B��mi�V#�ƌ ��E.��E�V����)I�QW䚄\(@��o]\�rB�5m�}ޛ���ew��o��e �������$:^�7\��,�˂�7��N��E�ߚʝ�,wMϞ�:#����4,��^'�U=$�⥔���4����j���㛯��ޛ��9���U�ڥ�J]h%-��3����mI�]@G���|������@,�{zY�<�3i�<RV*�LC�#e$.���Md����Aty�����vL����8(7���������3��W����&�zG'jc�D��j`�_X>M���spG���]=�C��tq���K.�9zyP-�;�k���6Ri/�{�0ikۡ�Q�NBUJAԒ��-�������m"����!�3�":�?=#j'�QT�D���?��3᥺���	##�S��T�	K>.�^���	{g�#+*� �{���ο��x�<��.6e�%wP_/.�w�vV�5�1C��mR���e�;������&F*���J�a$$)E�����a�j�t����|?���2����n��;Cdw���a<pu����p}����b�ۘ�e�ޤw֏r�ٚ|:�r���c?Q�������v&ƣ�8���MA�����k�I��� ��C��K�5MZ����MH-"�g�v�IK��3�f�$w�����Y'�x�g���!�'P�����Ҩ���V�wr�e�������׸��Nf�B���.�h�8��_�'���^1k)�J�s:_�������T;,�RH����X]��*�5�q�1 ���d���pM��#iJfQ�Ff4�Ff�+U0/�=8kȂK1��Z+�����̋�YP���%$ߞbU����{��B��+[�~��`l��G[��؆�� �(<{q�mʡ7�����ߕ.�x!TLq:�M�+�ʯ��%����wt":���Z����T*����]�k��N��Lu0�f�:�o9��@]�������Ύ�3�i��k�I9�l{����q�,w{򰀫[�{xf��'-*9WChU�ڌ���s�����S#Y|F8��n�|V��Y,,P��+��+�u��[�n�Q�V��E����X�T�kT0�~��r��TRE��2рI/���
>��V����g���鯧�$���X9.i/�[ۻG�(oŊ
�%��ae]�� ���;�&āD��'Dn�#3�Vd�˼�`h�ޛT��)/��g�}�M�r�*x��"�yr�0<�q��HM���E���=�`n�����52���r���~�����+w�AU#O��5s��Bx#&H���c�i}���
�8�����f+ii����Ⱥw�ii�w?�O�R�%|)a�/±{RuE�|��g�ħoE��?����D�ǾT�`6A�:+�uS)��cb�Z�0��W���B0��y�'F�'�j�{��������$t]�p�]v��B��n�Hi���M�පF�^�y�6j�c\Ԉl�IY)\��L�@J��Ş��l�/���8<��������n��g�D�m���-���ܴ/�Ȗ�U�
���X�L1��Y�Տm�K�u-��iMG�����ƿ<Y.����d���c�'Y8�����?����[k-��d��C���s��.%T�R��MW�|�\���xE�n ��N��`�.�Uo�������8,�!@�IO�xF�W�ش!������P~o�Z�X*��"{����,	�CH�ƾ����}˞}'��%��ub�!�c�a��}>���iy�^�?f�s�s]�y_��9�}��{�'�a9�"a�m9R�P��;����q_m'=�H�3U���!�^Jc���L��Qwm����M$d�6OrJ�n�w����h�^��߶�o���^��J{�"���U���C풼���]@����r05��"�	3�^��ަ<?w�ϸ-�����Q�����8��1�ŵ)�#Ϻxu��'�{�5�۳��!�� n����x��E���q-qWe�$ɼ��)��|9��!hXЏ�)?C��� ��K{�_+]����,x�H��R��\Tm�)<�Ձ��f
8��!����й�T��$�ηM&�g�:���]�:��),2�(��4�(�<���l�0a/��ggNY��ԓ�Z 3�KdDAC 1GĝR�%y�a3��.��0�FK®�rzRJ%�*��6��K:��r2���r���JԊ����T[�hїuѣ��X�SE7�-����^x_�6���U.s!����οm(O2�xy�2�-jm�9���(�jи�ղN룊$�����g��J�(`�o3E�=8���y���6����z6�4l�;��� s��2�?��d)�s����.�~�X��8�dz�&&�&��}dȀ���p���ހ�����8 <U�\Y\w�2.���KZ%�9���zT o}����2Fk�ǨF��1�OP���m*��ZE���������8"4}˼�$������zTb~;5U;��n	�-\E��.��D�p�ɢq�����~��Р9���%^����m.���*e=u3�"7��;n���/�6:���*�S�Ŏ�&�}�|��Kjh�p�1����]+B*%axݛ����[��k$4[ك�PN��g����־W��69/�%\�k�(y��&���2]��LY�}ѓ���1���/��"�<���sz��ܓP-	���9��g`⚽�����xiX/J�k~{����Cy�;pV^j�n�M"���#�j��-�`�)�dk�"�=�Q��TZ7UxG��'Jb�!@~�Z0�[j���s.���m�s��^L���Gއ�����j�&�u	="U�7��;�����J�;a|f�7�� ��f��P�ur������f"��9�;"L�_R�봥>t���)
(����0~��?���<�a��X�Y�_X辴��Q�{��W���?Xy�QO˲8lil8���E[��VD�Y���I��5[n�d�|�Z�v"F��,�CV@C�=�3�Э����7$b��uɫ/C}N�c#�ɱU����a�b/���Y���7�F��I��Fe�|������Zo�^)�����nʁ��\�2�ʻ���z5bF�Fp�u�*��`���u��Jy�۟�zܣLK�_��T�k	陔LW�SٳN�ɧ��Pm�%h���Cw	9���Hؠz3^;%�}<��s?l�3��>�W�7�[�[��������ݖ�ӫ����먔*�:�zh�q��P~���(ȞM#G��"�����k�u����[�d����5�/����œ�ip���?F����*G
'��r�x+|�f>?L��2�i��g��:���\g/�8�a�d~Y�8�g�Y龙[䀾�X��5;�u���O3��O����"Tȭ������̪�ڦ�5���g]��㘯�0֛qd|��� �=�y�s ���D>���Z�mH�6��\�ɻk����J�F�F9�e������U�Y'|{�B�2OSff���o�tE �c�j���j:x�";��������֙��r����!oH��*3så�I,�xb5���1�"�![�z�9���`�n+�o�*{sj���iy�u[���,���G��<�'�R2�V?�y���>�to����XH��OXG0����e�P�؟�&%ת�Ld{�z24�(�#�9��l%�'��@g��ո *��ɴR�$��k�l����Zp����n_�FV3���T��KH��G/�G�!�C������@�H�8�D5��Η�y����2��A�Eԑ:�����D����֠��a����T�7�$?��1H>&T_j���10 �w���h��Sa7�yp��T{]G\��I����"��x�/�e� �~"^��x��S�u(L59�?{sg��^���ݝr�I"��8D� �$��������j�P�ɀ�?حO����~鯙�*zW�<z)1�.����5�s��'����ca1��*O\+�U &��U�����)/�o���O�Ǔ&���C��`�7YN�⼂�`Ҝ$�"*SG���h�V��4Z���H����ST@�!�r%<�$+=
�_,�V�B�g�,"c��E��� �0��1���	�r�g�?�۸|b�%B{�|�JdX*��C�/����*a:�scƞ�0���������UQt4�㊗�?<Y�T�8���� ��{�?B�M��7�C!��W�DYȫZ��
��1�͜F����/a_�$���b���k]+$܌��O���ۗ��I��d�X�o�H	�`y6�|/������[����9e�K/qCҍ�b�ţY�&CK(�Y�m�پ�ɢ��gV�DDr���O���Z��o�d��3�61�}��HP�k�`�7���pN%��5���Nk��N͆������$dC�S-Ue=Ge��k���G��l�S��?�<�<X�_���c+;����gk��~z\�D;�(��Q�|����똅ϟڑ���	d!�6�	�XZ1\����i$!�8����ǎ��F������=��?�4k�\�������L_�2�y�����Z�]���tUv}��eC�%}-:)"�}Hz�QË�A
�^��iWnU�~�I�2:ʤ�tF�/�jUo識t7�I�v��SG *=�z�co,z��F��T�R!<����D��W�>\�������J��Dֺ9�W˞{�H!��"aa��Ź�)����ޮ:h�^4 &���u)�s[�Nh�)�_ ����d�@󘪭��C8���ͮ�j�D�;}LΨ��p:�D�Uj^�O�+%�Tҳ�x��{�uϓ�)�멡��b�g�4�4��O�wm�(&�b�jq��:�5m�@�,2)W�]�S������r@�'I�8l؞.WU2PϾ�;IoN_��^6X6��ݧKb�@{c~n'͇,>w�X�[�)=�������;zz��M�Z�P��s�{V�;Z=�X��3��X�.��\�Z%���DW�X�z������'����J��$��:.���ݦ�כ�d��{�S�M�e�*U��?���r��@�[����������
a'.�2�K�O� �JW5�y5A�GD�+¨�*��$��J�Tm9 O�O���ޟ�[;��H̹���s���1ڐ"�&�ݝI��C�wk�ߏ��6�˿�k�d�Ni:A6�����n�)扴�s�[c:�`+��;�1(c�����"2ȹ0Ҵ���I{'奥5&��l�7˵>ݬ,�}�oZ��\Ԗ��qQt@�
�ϡ8�"�Gw���,6�6f�Ѫ���_��x0o��D�cgC�������YG15���k$��
K��r���8��'4H��(���z���d��mzL�:��<��=\bf5󭦆���ؤ�z���0�ҠN&W��!L!����;�x����}�F;�ηl�ߙWx�f���d`SJ���w���|����F�钡s�Ҡ�I�����^r�!�S�\�:;�@P����B��N?8G�������Hm�;��lP�N���>���f��k��OÐA�hD[�g�f�����e��)��Q���B�<6�ĄI7��P]���y}����8�K���
_t4�c�����=��*}alqL��K�>�B�oM��m���'G�A������dD��vW����t&a|��"T�o�����߳��aV@j�*�w��0C#8\f��|,��U��u����ȯ��`&��ˍ
�0�K9�X�d����xY���N��!���
�of��&�լÊdr��fd�5��%Z�}	;�}�&����zߵ��R��r���-�q�/U� �ŻŇ�,6A��=m�\߉<-5��dWQ�^�(�+��h3��c�����/��f��wvc�U%8<$��Y> �M����>��vw��
�6��C}YeI���]��}!�,Y�����y��T��Xb�'��z|��z��G���}�!x�$����l��n�+�y����n�*�'vjx���$�x��\��L<Zl�������m:�qIw'6`�q�j:[y�O^� -����z����mi��ɷѼ�����gY$ �����9�?��zd�>�$���Eǲ�_�Yr�Qغ���8�+�p�tCq�>���"ɬ9Pz�)��c����;r6�l5��wҜ5�E�a�u8t����� \�Q���'^��JCwC(�TN�)�8r�(c�E3�����OX��j�����[	�o �D �\i�����W�n�P)MȠ�%�n�&���BO/��Z�׽2͛}j��KN?\�����pG�CѤ��
w��0�3�R
���^��>�>]ug
.毖���*!���"C�!���b�25�:V ԋP�*W�vv.�Lt�$ۣ
�	p�+&�?Z�\�6�@��L,�%A�1�/ �%r6o	v����`�#V����ӭ�w��CH�ia��B�#�B��屡֝oNzPGA����y\��[dā"�o�=��8你j���Ͼ6'��ilm�8��QI���ۼq�vP�������8yO��� �`��J��%m��,�!D���3T�Ν�7;��3$�⊝"z�F����]�=���9dE�/-�/�F֔$������8��r�A����/y�^)SE��N���-�Pe���;�7V�?7e�߱C� _5������_6�R��Lk�uX?pXA/���ihn��M���h�'��	zX��ù�0��i:�q�Գ�H�3������×>r�yRn],	:��Zq��rLC������h6vQ�;]��r�[{a�'�˺�􈏎�;ZWI��%F_��a������c՜����2noK�N`8XB�m�$rc���a�,lr�p%�T����2�JX:G��n[�〤z��%��U�q�t��A���/�Ug	S��K����g���c+L�r���!Hf	���U'��k����{�D.Q�)��*�Lc�����I)�+�ŘQ���%XU��ݍK�!I�������ɔ�SN��!{5U>@Lm#l �׸�;��Y���=��q���7�_�ˣ��l�e�xRZY�{�c~M�(��7-���O�%X��)[�&P���{���j=q$��
9IO�'�A������G�?�^�
�4G�S���'���A��B�5o���V���#��!I����A�;�wR���ud�xҋ5�^9��A��H�T�]��=#)��A��'ft�7FI$�uӲ^ي�-�TX$��gN�3U�������s����jZ�N&wӞm���^,��� �B��g�ψ�\���++"23���0��4��Vng����V��64��_��"��H�@;Kɵ��A��3��,?�aT1C�<x8c���ҹ'���R[���\w�E�+�v�G�4����0s�r7Ο�]fv�ʡ\|y�}�pXkcL�qQ��ՔWmɰ$��I1�����P�cf��'m^�t�B�=�3�	���m����"3���vq*V�L3�l���D��.[�r1+�)f5�p��VF���@�鶁b��m�~�\��>�������5��҃u��R;����,�} W�����Y ��d�X��1���ڈ<l����*��DS����SF�ߜ��sn�?��0�(y�s~�����3� ���iYt�����������,츔Y������F�;�c�a�׉3��ٙ
��ܯ#39�cu}v[�b����öZ=�\b.{���кk���h�43���h&�_�@}?����q��!u�j~t>%�7U���d^�9+db7���HG���q6&�%$ɏ���9S�ɿ����6��hש�%Sf��G,���6�p�`.��S��3�ajb�m���o���JK=��ɟ��`�r�I�1L�y�,�LH�]B����NM��6s��o�aUv)C���g���I���E��`�窖�3ś����c�V�f�zJ2S��ƚ�O*{
����n�n2��<�Tz�� -�c�K�rkk��%_-��������>hn�sE����v��v��@��#�^|�E�s��n��J����}����[��Fu�Ź��[��G0�cU�چ�Y_��p*�����W4�vn�#��s�����_��v��í���9` �� ։ˈ�8�+�=ѱզ�kYo=e!��1{-�Gw�ߒp���|�y�uJV�	r�|��$���z�e����n�_�����������r�9�RM���HQ�~�{�s1��k�+���� 3H���x�_$
�E'TScK��!��^�Ӆ�N{���O��ϼpFԟ[�"����z�u���G�5Y9*��{3���t���w<g���6��#*�P	��2Mi�|"��N@9uw��V��\ٯ��H���Ӌ&^]����B�RQ���UWY�s�g�hkh�դn'�/���	2�n�
��2B��5���s�P�Sr��Єo�U`DV%x�d�DA�~܎����@S�A�m����M��A����~%��[���i�(���C�����*��6R��o�=
��b'���������0;7�Ǵd�2� |7<�3��s�M�ѕ���"]SG[4���/�:1����܉�$���LNP=@^�a��}<��X����X���kh^P60�2 ����%��]����A�5GϿ��s8������=y�*�/.N ��z�'�Lٍk����wa�ƅh��\����ҫ���;�ƞ�1��Ӷ|��=\%ص��k�m�u:����>�@W��f�� �����������7&����>J�㊻��b�ߢ����4�޶s�*bw�qr�哊��04;{F�T�~���/D��9_��ٿĞu�ѓ�����[�7�i�(�A�a������35�g���j�hZ���W�>�y�Co��ޚ�~q��_4�����v��,���Ѱjj�_Y���K��墰�?j��8l�겣T���\��A�����F�����6v�,"�osd��_%���ߟI��my����E�S�������dl�3!�"ؕ�n�	�Р��������ח�b��[�'�m��yW����m7f��`�?R�PV��Q�悧}���2�w!H��	g�EB\qs��,B�����!�U "h/�`�ܖ?��4�R�:&����\�R����_Օ�}��3Cxqd\wRh�r���^S��m7w������2fB��� �.��1 ��P��B���W����$g���斏��3L�o#�!��ȹ�FpS^�妴�v��՝e��;�ffڕ�T�}�7�B��K�<���unN/R���ë����5�+ (�BM܊���?���7��?����)�A�������_w�Φ�5�K9��x�U&v��K�Y kr�a�$*��UϠ3���{�ĉ����.3�4��SR&ھ�4:D�ov(j_�k��[1����Z��B�-&��.�Ðw��Y��z��V�6�̞o#v���U�[�;�앉�.��%��V��D�&����\��(���j�Y~��/���kˠ�z��a��K�F �^�$K��á���3N)�G
��V�d8�uZ�ؖў�Jy���I���!a9F*��m#���!�����]j~�e��n���ʁ�)���Ȼ��F�x]ժ�H}<�����d)��kӁ*ݾ4Ht�pn�+z�`�k?� �:���g�v}�$N���NFϤ���=��&��f�������}����u0V/�w�����i��o� |��j���!�c�-���8䞢����]L��[L�ze����M�ON�f7�DEr]������A^x�b'�H~=w���ZRĤ���z1��ŵ�fn���qf:]˶T�� �����!�$�3	�3�Z��e�u/w�~��]�3�D~�QV��H&������T�l���ڷ��h����=~ձ��Xre �W��Q�a�ǵ��=�M��J0L������"ߺ$4[������Obw$ �Ƥ��Uf�a�Wֺ9����k=���?�wٱ�Q�[����[�|v����.H����R"���W8<��l]�3��~��hh��щ�ڇ�86L�>�Zj��G�r�Y��crQRd�=枏sQ7ϩ��N��ƿj��/��]�%�ǎ9H�*���$^�ջ��s�ǘ4pŉy��mlM��oh��ߢ�tf���љV$�Ez:E#�ohXp�`����ﮉֈ]��K��JJ;x<�������-|`o�]CZF]٪�0_�w�w�,Y`�^�^��&�hf�&�L����6e:��F����GcW�4�� ���(G䚪W��?{��>���n�[��ajz3���/e���,7QghE�ʖ,�����P�^��s�����/�Į����a����T�U��3a:7
�Ǆܸ��F�	��$3�ի
���X� ���k=�{%{z���BXm��i^8h���n&}R�7c�B�v��r�W&�}�+��	4�$
�7���|��Rs�o��ќ�:���z�Q�����ᷣ�P7h=��q��:���ϲ�<r�Qr�&��'�r��nUv����Qz�\I���'��A^kk���m^!}U�=D� �&?�7�a>oe��P�~��W�5�Z������S�p.3�q���K�E�"���z�.q֥�R)��X�K��b����Z���0D��p{��07ە�a])[��+5�TjxJJ��X�������[	t8BUA�8V!���^���;� Lī�v��ܳ����^���;;�o�u}�����e���h� K��h���T��*��)C_K�)"8.~7G$$��9z��+�V3��3Ӻ�\'�vC�IC�;�}O ��P��:����o������N�$�v��:d��È����U2#Fb��ʲ[S���~���n�(��έ�������2[�
)63�E��'.^+2��_�=C�~qm1��X�:낟���53��C����F�?��G�c@�[J(	�h��l���JU�8����y�^�nA� �Q|IU}�z�<Ӆ�yb��(ns1qr��������'�r��"6?N/r�O��P0#2�Y�M�O�����i�
AC�%m8�xXBxx�vh��;R��k��?��rdD���~���},��q��(�}���_�Ow�E�>(��8B
���/	�/�>a��B��˼W�gPk�Oy3�/�f�vqŞ�����=�#a��_�X�����j�[�����K�}3���c����o�T�'��l�T�I�욄K�8t5l��`9@��{SKico��ߟ���\���z��^�V�}Ҡ�Į��B{�q���=4�>���CgG�Ç��>ճ6?��cY8�8���U���/Ͼ���� Ll��"9ެ�6�����<�HrVw�Lx;�?]-p�b�
�R���j� WRWU8f݄|�}/��؃����O�z|򤾻�����L�7r�N}�7/J�Y
0\������¸��t�ϔb�o�/uU�X^�~"�˧/��؆f�)��'g� �D 1�͓��V��[}�IE^�j���jn�~{��a�h{<K�m�(��m�i����]�~�.��N!j#���'�B`׬��1b`�r�p�>%C��ޗ�Ւ 窨����]α���"�h����d��ػ��[Ţ���:�E;�,�=?���lӍpY�~w';	Q^X��2:(��|JE���O��83	��
+a?��0�����Pg�xu��
�m�©w�A)�iw��P���c0!�����v+�#�~׍�+�h��� �
D�ɓ�Age��=6�g]
��t��d������*�[E.u"M����urŦ�����-����
�#|�d�o��e�Gmu��r�55
 dL����B8���pc�₰�"����#�c��W�h3�je��\�y���7�s_�+%�=ӛjU^�X��b^$�1^!M�q�u�.E��4Cy�g�$�z#�Q�+ƃ��K�ki����	TT��ih�;�Q�0�a�x[e?ƾ)Ǜ ѽ�r��U�m��O�%�9r{I��:���%HS�?�VQ?�>�����_tw�|o�8>OGƴ��9�e��{඿����@Au���f	x�	�^=��,M�ز��б�*�F���aB��K�S��$��"�5��wrD�K��Jm_��7�����{�cK������ ��?Ti=o�8��Ye� ��{:���m���hM�\o�~���t�2��Q�v�@u)Oee|emw޺���#wy��uϘ�D�H	Z近�^][{#� ���"ĝ�O �:Rz��i!!Y�����*7>����*�w|?��O���D6tU
��,.�<j9��e�L���I�ǉ�]�ϥ�:��'MV�R��9m�"��_b�T���$"��կq�J�"h!]-{aɕ�ė	6�a��[��h�sԦ5�)����T��I��N5�e�a��m��Z��8�=͖MF\='UZ����1�0�C�EWԥ��P8`�rP��Ho\�Q�Y�# ��M����TkmSS,C�bF���^��B���
� �TA����= )к�d�]�!����� �>!a�\�����@ev���,30�EN�S�8��M@��ܤ{���7W��W�c_EF�V�vz6!�>��:?��G 3~Ӑ�pm�,��m��b�7��k�V���L!��0�c��ۏ���u�߆��Q�/��ˍ��v�A�B[#��Ml�F��� =4/�N�?w�_���N�Y�{ �+�Hj�N�ރ���^+$�hUɹ�C�����}����[`�߸���+�w7+�� �5���p��F��^��5�a����xx�r۫�T��p�N!�v�=1���e��#���o���+����Jwqձ'���6E�-G��R���RX"F/�W �=�qt{�@k4�T-��t��,w���ɮ�!��k��DGi	�����!?NpW�;�~�~$:�ᴗ�&�&��v�ʑ�	�'" 3�2N>3��1),4p��k������=}!�W��c��1~?YX��Qg��VG��d?�<�>� �>Z|��1'��T�1����d�!��L�=�����"��
��!	�ʂ����{k��u���փ,��$�+)��+�Ȓ3� 4�)�o��p|`U��s�n=�>|�xc�߯
�W���d��Z`X	�U(�&kD7g̺ `&��%7���e���E;4u��7o�L�R�����{�`��;��|y����Ω����-���~����Ʌw�a2S�}����N����|R���^� m=�n�Z�,VV!��%	��!��m�|�En7
��v�gǛ6�SM�ߛ���p�8����|����xgdf&�`�[��w#��^E]ٯ_O`����ݺ�pt��� �J!�C��9��Nn&���`��m��@g8~`ӏP�7	Ɖ���Y�-/�<O��G���������GI��Ԍ�Z5�7O���}sL _a���y��?����Y� F��Ef�0p�^��@F�y�DC�n�,g��>z�w��w�����i��4�P
�P\��X����b��t�B�1`^?���S/���)����?�o�Q²Lշ�����V�_�bb6G�z��>��<S'j��~U�3x&?��rJ�8SH�Dz�5�Xroقg�5,����!��9� �(��V�^6/��\��h>̷���ۆ_X�':P�#o��S0:�[dg�(�����Zё��`�2Z��.��[M�eF�_r`Ō�η�R|�wa0�#r��ߊ,g�2���4��U�Pt>#�mƛ�+��/��ß_э�u�2-iܘ�1�~��{DLQUB�;�������>���O`,X�� g%o;�(k�u����G��Q.�1�٩�e@�ސ��Xv E89Q��ԅ́sQ�u��y:'\"���ť8\A�C��5�sOڑ{�c&�I��#���*W���8[�d7�Ւ��аo���9<`O��0[����uU� 5ƽ5h��V̫�7�Z�z�Q6l��+'��g���o'��b��?�m|�#��|?W��>�����3c2q�OF�k����ɗ�8���L�3�R��VS�>T)� [�ii��2���S�����"�y�B��_,�����Ac�}Y�����d)��-�oD�G8�I��ޞecJ/�'�K٥�X|���]:���E��}����׊��)�%qx�%�����i>vaKk��d��R���bg�ƚ��g٭ ���dЫ�yE�]*�A^Hu���_v�6�^�+�#2�w��� 5!q��측�ٵcVab��\��N��lo@/�\��/2��W�ݟj̞���g쓐�]�?ބ ��U�M�yē�>�>g��ӗry�X��/�vG۞�\P��SD�`����+_�6Qm��]©�
t���T�Xx�����ؙ���L굋�l���>���IW�z8�x�Ճ���i�v��������h@�^�ȉ��[ ���Ou�S��(E8i�9(n4| �<�*vM:)�ܨq�g��WR�8rG]A�C�ݕ̖q��y �&)4!ؔ=L�f�x�����������V�W�@�U��j�.U|_Z,��QbcEf�E~!Je�ށ�u����|�c<��_�t�o�\7C},��wBoS���͡��_�8J%fm�$�/^g1,:k{%;�<�r��q�B����8�cU��_p0<��.��0O����O�'N#�S�@,o��H=Z� pB2�Ln Y�6<c�7�%MA:j�) 6ꏶ}�	�	�����]S�����z����-u���:_��,T��t ��P�u;6������GD�rG��$�8,���xj��+�ng����\��y��O��A��^i�W)~�*$�L#�@����p��vcv�mSNy.�H��;�U#���ܢ"c�8c�5�C��;�% :JV�Msy��O�6��"�`�%�����u���kv�%5H� ]8�`��9:42QD����*��O�����>�A]�\K�1�[��|������O�'��ǕG�W/:�u�Z8\�y�L��[ۼ��Y���/M
P^\���b�jw#a[��@��> �[�j�!�_ ��8��= r�6+1���vgCw5,�v�*6'��۶h]0��25�Illh�[�y�*����joE��/��lNq������br4�����JP2����˪Ff��������5�� �� ը���b:����w !8UiՓϯG]�g��Qw�Hӈ�a�.J�#�=YMڼ��E2��S�	[Q�fW3D�W_��P��	��@�paI��gT��O�$�g���f�}�Jw|��Ŧgq���c>����l�����+%p�*Z�����ZZ�ُ�G�%�sNׯm��\]0�{L�L�� �0��S����w���A���L�"��W��?�Yļa����θW��8�Ƭ�~���b��E�8#�ȧy�������>�ys	YO�LK�D�lW�`��]�罢��b�D9򊇉��No�����#�ڝ�c�`�X�����6�\��ّ��Bv���ɤ{ȑ��[�����C�u��CE5������㳹���V�[7�;+�����fϕ25)	�}��K���^�΋�]$��")t���X~h��  {r{�,�bC�
sz?�"�pc.l�!7�޾qu)�?e��T�܇!Ȟ�^j�d��Jc��:g���6m����ƙ��L�J�������,�4�b�_��Xi������'4^��K�iloYY0��}�?�^�-3X����C;�Q�b�v$=��	�j����{��bfVV�6��5����,��@<�(�%Ls������� ��W�` �����O�$9�׏xV�5� �������I���9��?���.�;��m`���D�wg��3J�~��IQPg�<���b`�p	����Y�8�C�����3�%qH�	�"�p�I�UG*k,5����/��}����ެ�q��`XYl���@ |���dc����#RF�7|�V&�������f�^R?Ըo
*���ظogH>s "�zX�I��� �-i�D"TޮQ�?�n9a�˗K\mƳ־�^���j�z�uY��c����S�>�Zf�����~�-�L��v�������P����!'	4�M]\�y�g��Z2੣�V<�n�~>��z!�V�-�V�bWb����wJ
�{�q;m��-w��7j�ipɞ�uo+��"�Ӯ/>�N�}��R)g����G�_l.�T�VKq�������W_�H ��t:6.��1C.N�[&%��-̍C//ns�x�xY�- �6V3}���/뛯���yo	�~�ɑ����#�S/�[��|bb��O��ǎ��C7v�x��M�+��4ze�$RߝrT�������>�
}r����N�^�dwTGӦ�
�ގ���Y[�/�u�ǟ���i.�q}�O��B�ѧ���� �������.)�&	���G�(��|H1$Ma�mD�	������F���z � �H�՞��o ��{+;��ʙ��{X�(Vr!���phwx�r�u�=�vT��X �y���άĤ0G�ON�&8!/%'I�������`Wd�����p dǿ��Փ�0�=@+��.���H$�@�LMkQ�?�k���"�6��>�)'�E��=�v�2�R`j�����VI�I�������oV�S��O֩F�"�L�i���/0�Otҹ�Z���+����(Ŗ���X�����1�������^���:�˥���v�&�Ҹ3��E���=ϩMw�>c�{�q��~��^Nθ#7�^�r�j~��)h�]=	��r����W���/>�G�.�7�`i��>���w�]~�o-\�6]����L��1�z=��u�T�gd)�`�s��n��S_��i0����i<�±�P�����F< =��\����/��we�}�s��!��P��/�a'��.��D<��5��آu�Î^���������QEU5��QX#ԟ�G_c@`ph�V��Y���׉��ܽV����Iƚ�����v��js$��禇G��ָ���hbr���1Ru�1-&�=@�\���x����y�UVŅq��>L;w�'��5.�7F���V�5.J���yI�#7�!�/������e㓿<�pW0Q�����7Ѱ�Y�J��S���A U���0��"eJ��}�~�Ү�z7���É�j�'A4�	v-+S��R���4,I���+?0_9 ��]k[�G�jVAW6en ���3��o�"�D���X߾��=1HK~"ԜE�����لIp�F�?�3�[yV�������N����4*e3��CZ�w�=�t��	��g�ф�l�����-�Dp�æh3�ed�{F�@�S�~�o��yfvLЃ��KNXH��W����a'��IL=Aq�C�,Mm��>��"��G>�"��+�+(���I�.E��4�̮м���K�>mGn�
R�r�q�!�i"� �tt	N!�z�Sd��f@���9<��[m�Q�D���p��?I�iH��D��p��1/���da�Ǳ������mz�8��'{�%Xuq���]�?BT]�J��ݥ�����"+_>��_�����P�N�`�o�%�pCɖJ\�N��9GZr��#A�}3N_��SD�u���j�D���u:����)&�N�j�t!݃����Z>O�+���^�����_��J/��cڢv�*�>�c\f�=6��ж������v�(�7v{�v���{�)�ԡ��/�*[U=ās%��XУ���ئ=Q�Q�[����_ކ��r5���U��5y�Ƀ���oڡ��*�5 �b��q��B�z'u�!������W�Z�vv����"�r�dn�(�M�s�(�_bt��to����7�7�L�Ct*[�a�����j�_�ٗ%zH����=P2f�v��7u"̠��`���ݫ��wYͻF`��h��o:�P�x��P���y��n��yʌeǵ�Ȉx^Z��L[W�:|��kѷ�6v�_�C�\�m�1��޵?:w����M�x�����y�"SË�@��=���/��Gm�,Y�����(ٓ	���UHW�6�%��&���r�[E���͞����8�RS��w��U٪eT�^�A.n\r����A&���K]b��ZQ&��y��<	\Q\���*=b���x�"��q�p����&�z�Ja��ts�v.)��s���R��ݲ�ꐸ�m/p�N1���5%!_����l�H�2h�6��Ƽ���4_H<ts��@zp�C5z���׭��+�����'6\���K��}j��Џ*�T��gmx�dI`��{��(����&��%�]�+�:�#_lq_�|Ǥ9n"y=���]0��Y>Kp~�q���9=�Wc	<%�n�b��<>Vo���B��״�ʩ'�Y�:��#IQs��|��JH��R��RS�3I�>d2�d�t��-�`�U����-�|���Բ׾��Qs���]����p��B�ų�
 P�2��M5��~{�Nz�<�Ґ�kc�Z΅Lͭ�����t���<��e�p��r�Q���'@-B�rsN�B�X�5�7k� �k$/�e:&s�3 �m,/�'ߺq�C�b؃8����}Q$�x��u�����"}��rĞ���q���*��e_||��!���c�:��ڢ-6�*R�7� �&�w�Mz	!H�޻�@BQ�B�H�I�����3>�3�7*�ܳ��k��}VҿB>�M�H���l��-�ݱ�Ǡ�Yy_���Mղ�w���HWQ|<S9َ�C��	�ɿ$^�+!���~�>�G���?G���Q��k�ҵ�b��$�ޟA��2��EmҘ:��~;n���?� :���[��e7ɮ,��u��RJX̷�&�7@`���p$ftr�(�{*B���X� lV1�V���/N�����<�U��mk����U������?ʔ�,�S'J�>`Y�V��q��n>(��o<*�iW��!�Q�Ǭbp��9�����4(�����W�C�ʪ��s�0c�j<U�������d�v��5�N�C*X�{�O���37�I�0S �I�$�t��&J�^��C��q`�2���!s9@{ǂ7��P3��z�|ː�P�o���4�𰽑6@^WNܮ4�ꊂ{A۳a�f��C<H�L��d��=]�R��0��4����]\o �O��T~����܏mϳ�3::8��O%q��x�M&��r>�%S֏L�Ǵ�Hu>���&���*Ȕ��E�����C�y`o�xh��^*�8�r2���F�8�a��|yVue+@UT,%�^DR?E�?U�U��[y�w �A����o��|��Eq�[�����-�F�$q�������I���lBZ���c�2�H���$�P��1ś�ψ��؉7h�+�6/���M��o�6�"?b�	8;��P���U����>��B�涖&����M҃�XQ���D�^�l��И��+��Y�4���3k�P�\3�g �:ܿnb��> �)���@����@o���>�K�����㾛��n^9��>�<�R��>�������G$f4�����6} fHž���ɗ��s��?#��K�� �釟)�}�h��q�)A���Rڳ����e*E.����b�ߝ��Y�IN����oE*Pr���1j�	�Nr-XF؏0�����˗�G�a>����+�N=p�/i��~3i�/�O$PE�2�. e�;Mء~��_LQ ���yW-U�VA(���ϵ�ԇ�u 8����J�鋁3��4�U!�F��=:ϥ�<E�\l����0+�b��ST��9B)�I	���So�I1�)�˖Y��)P�?p*�}~�Le7C�(@&�A��p���`���v:�`��Dڿ;�/��I�a{x��He�M?�|P0�[����v��hw���#e~&�?,rXrKd�繝O&�����������!]a)�������͵s[�~&~e��s#<E�JU�-35���G;l�Z���:R�N�g2��=�P}�-<U��?D�bI���(nk;���߳N�;K}f�
�=�Rd��웖*� ����
��Z��/ܚ�a��[�����t�Kb�
LѣB8hH��Te@��.�>�=��&=��c5Yo������[՚c~���&�L���s{u�b�v�n�ƍ��Ҽ�3&��U[�G��;p��G"7����^h�+h��cg���=u�:�!��+ �{G����0���_��E�ZqX���B��t��&�-����MY9���c$%�����ms|�-���pԮ9m�N�����O�ٞ��lu.`���]@��,�F+@oe�πs��^Q�2<�kl��\V0j@�D˽b�A�]�C�ē;(��.�� \៬^���#�Y Y�=�IY`I�0�8D��Q(�Wk(vy-��gcS��c��ǿ���	�n͖a@��Vx�4���_.��r{wa�G
�9Tg���Ӕ{;�]kg�Ⱦ�#Ok��]�?�H��/n_��z�)�A)M�e/Y�� �W_~� b�#E��Br���^���iC�ۋ�����K�*��#�5�e
Ũ�y;�+Z�>�;{�}
��\�ض|U沜��/A[��O7��:��ˍo"�?řIvx|\��8�sp���ӂw{r��h��y/k�F�u�-#+������?���]��`���l��(@���qk�-�/�f��>N3��C����P5��m��$��(d��&�_v_�6>�-Qx�#?Ӈ"� f��2?��@������R�O����-6��G�Ҏz<囒[S�Ml�P)-l�y﭅
�x���5���5����ӴE��`��P�3�fQ���tZ3)�{�?j�5��:=2�ۗ�����$���"���Qmɏ���Hqg�'xz�o�!���p{T������㹗�*i0�cR�����B~F�/b�j&B��
�1s�l6K%/���{/��.�˵���ޡ�Hma�cw=�䠹-�o�`�������[4���)6�r�v��U&G�����d�w��Ӷ=��L��������P�ǫ��^孖�����捪��B��!�!��)�3#e���$����)�����	�@���EE��l��U�����J��.��ɏY�5���H�xv$q��s���	G���/
z~u:�v8�N�6g_��O���:����S��|��.�3�G���ƿ�鉦,�P)Ga����v�75�b�0�.���/��T��?F�f������I�]L���pt��Tr�VRO�i���^���'9ps�Fzd���Vuv�`t���I �ǐ;`&�]�+�m�*<��ɝpL���)��1r��ք�9��T1�������w-^F1�:v5�}W� .�������Ԅ-Ǻ DK�w|-;�d��������L�w["���$XP����b��NT�l�u����f-W����<)waa�-�����r�����oG����͡�ѹ�8�Jc���O�Ʌ�>\3��WEpy#���u<�VV�Z֐+yu�L�d��\f[�5�����{7�(L�[eΧ�����) *f&Z4��c	����a� �Z��]��_5��+�m譸�eU��x��jU�mN��t�G6~x?��4�7ذ�-���\���gǦGK]�0J"b58�R�!�e��1��>qJ(�a��+��@n����Yd|����eH���"92��
��M�V��:;8�Gm)�W"}[Gv��Й�Wm�s���R�5��$��?4��4�ɧ��)�7�~��^R��q��^�Ԣ)�~��|KU��\gcz����6� z�����^w�kJ5M̈́��E�T~�$$h�\��M�Rs�2�T��t������b�C��KkP��W�3�r
r؞�Kn��[W���O5����Z@?��1���G�T��T4���Q�Wbrt�S'+<���TN�,�Ww̽�d�z
���{R{�[�ϙ�i=�1l���3(���:�t<*C��z�9�� ]됴B�4fYi��|�J�a�tL�l�nl���HU�����b*O,�:��m%�p���T���6e�iY�������!����*�g�}o~�Ǻg1ec=�'a��K�������f���f�0��+���)iL�.��)42�ɹ��K�o[50�-�Od�fa�:��!^Ƣ���>�Ÿ"8��$T�C;�d�0ʋp�7�|$�^�Ƣ��@V��v��$x�|:��ݼ�Zl�q���L�S�����c'��E�,���, ���Rk�{\b"v�2?^�-/��*��B�:Z�1���6=�R	�6[e_Y�-l5z1���%jNM����x�❪WM���.�Rף���������[Xƃts�Q �YfZ�G�����((D�x�{���[ g1�Ͻ�W�G^XtL-*����G޲�	��k�)�FBBM�`T� ���^�F�B��d2��D"���V�3������Xf��m���sRM�6�Qg(�~�|跢�����`��S�/+���_�g�qz�^�k�6�q��6f�9ڦ?���n�KF�E�����"�V3�M6Ƭ����5 ~@���Ƅ��Lݰ���{/ÜD�n�(����}R�+�<:�:+)���`q�&!A�����lQ��p��4�1���3�G�� ��$�)�#i�������?�^;�.�%�L���C=�Z�KĽz�`��W��������1����"�i&�/��=�;��r�(���Z�r�rD�'��x����ld���֠��0 ^�HJ��І>S!�g􆟇�����kˢ��ֹS.>��}mm5�Ts��q6�	ڪ��e���Y�������B�G�"�ٶ����-�9O�H��8�*;�'��S���c���'[g�^��I��Kޫ<C�]�UW�M׌�t)��p����0��б������ !�J����Mt|f�ӻ1s�r��#�zԜ̖���&�Xo���e�B]�<��21 '�S;Y���e���`�I�_�KV�1v�s8v���,9�0�Gg�[ ��T2���?{'����Ud���S�潭Fi�bI�]�����2KAb184�k���W��0�km	��2~�|��G�ZMl�����+Od��<�1�hj4��� ��C��C�%�!K��.~�1ֹ���5sȷ�>����Syk��i�c��Y�$���\�?�א�����p�&�%����~��㘼����G٧1Ƞ9�� ���<!�17�Ԏb�l����=tQN��5�A޷�?0�X?9ݖ,���|y�޲��P<$�Bsi�GˋG��O���	�����_�w�m<�i��kn���?�I.�:�G�s
�\r|� �"y���J%��C:�j�a���6 qϾ����bk�t�蓲Wt��v�-�ܹ1Q� f6s���8gѰ�@�\�����!�j(�Ԙ�o�쯫k`F�4	p�Z5u2�@��)��c>i>M�q\�薦t@'Ǒ��*��Ӡq�����Ds�1��?)M�>�Ǿ�S�~�u�T�����I��#���T�R4��Nmk뭸���2@�qs��xo����uGM�vY�&�&Ɂ��Aۧf�VР,���D�"��tb��gz*r�QȘ���/;�t�=�^���Y*��/-;Tu�@w~���Z��o�"��j�{��.q�T������Hj�sm���):��y��I�:'q;xQ�gx�6�KBB����j�I@c�AK"q�qmY͸�`)q��w���m���Z��+���E�)����+��l�����D/�����D���{����5;㡜��=j��L��s`x��X����V=-�G�K:��עP��\>��D��o{O�ͥ
�B�sF��uD�������u\��J��j�y4�q����`�!Y�t� ��X`(o@!턄��6�̈ć�9��^\�2�9�;9�JFdަA�W#�$��9��<%�.'QtϘh苞4�����J������vtp��ZZiO����J��D)+Gu��g�>CY�:�apPEm��cW+��*�r�w��ov�MRg�����g��l�]{G���-?,B|Z�}�xWRXj?��d���Z1�7�Z}�f���dΦ��5�� L~+9o�|�*h�:���ţ��F�;E����q���@�Z����ՋШ(���)z����'���X�`��T*F��Q����k������N8/�兼@�S�5�Rs�bL-�����|_�Y���5�	@�j�'���p�'�x̤��'��*й�Ҳ���z�\޾���� �k��d^�c<��jQ+e���Gi����F ���h�|������Xc���n��
N�v���_A�Jʊ��b��z���TY*�!U����o�7�
���,i°{���s��r�7�<�}����σ��Fy}��,޺��P��_'"<�7%�B��d2�:�f�w�Ռ���o���z_���oؕ�\z>+@���C�������ĩ��n�˾λM�+���u�;�C�\�r�'�ҵϰw0�����t4|�Nv�MU�g��o�^La��!yE���$�dJ����3���Q������Ù!W��ufF�W�7bkYd�M��/�?HcȀ�C#����a
.�vc�TS����.�u<A�$E�K�|[�a����t�N�x��D�$�ׯ�m#�r���uV���f�L�Ͻ�Ë4�[� ���Z��fa�s��y���Y�9����R�����c��F��Tc�|Q3כ�vʏP�W��<���JZ�xU^�n� �CC��T��\��v�ja�X������(�\>��C�?U��B�Ϡ�2�ɬq1���8��%�O4�]�B�M���L���TS������8�j#'��G�
K��@@|Hb}=X�"r�<��x����Y��(���B�׎��h����0�����>����P[����:ɹ`�٥�uV�f�S�3���K5�N�������\���[Й�����s�dϟ����{Y�97�C�e8ESQjEz��GC<���Ի1��Q2:�^�j`�����җB�DBJ���9C ������Y��;BB5���H[������Rc�.ǳp۹���튗��I*�����m�/�� �$�$�_�~f�5=3b\�$�!@j�t\��e�}X�<>j���/-hTR��Zk9�3�_k�<¡P�*�A�����W��឵,ܥ��m���	�<g��/l��=v�����&��ǧ�Y2��F#N����cc���z��e�Aj����w�^�1����������H�E~���J��Qfe�c�z'�_
�6n�m�t*�ϕ�"?��7_H��'[��&� 1�1BV+�E��X*�3�1�{�wPg
P�3�ظ����Y��wj�L3���.)k^ 8ܐ��'�d��0)����W�X���~�B=UH�w!`�m�Л��2�����u�E=͏��`���w�?\�!&"���R���=�aX�p`j^����/��=y�i1#�������R�îw�|n��JY��H���B�������;*�%I{��._�F45�H� 3KgB@M<��1������o�,k�F,�'����^ל��uupe�c����z��tE��_W�G�^9*sv]ŗ>��j��ih[%ǈ�AM�?|ȉƟ��/"/�obt�^�G���$� I���k������l���1.� H��~5,@>��\EOl�8hkvђ��Q������rW�����6�~�����"{HU��Ա�_Ǽl��/~�YP|�y�a�.���r�\�8�&7���F��C�b��L�c��B��?Lϼ55u}�7�T������}N�on�w4��U���r5Y��ӕ��y�C��G�]��i��R6�{Rǫ���	 $3�	�>EbF��vc��=I� FYXȞ$jg>">�&�/,ɓ�dz�'�t�6����X!�'�ɁО�c��u�!�۬ ��3Gsʍ'���Igz�ͻ�o�ϟ�7�҅����_�a��ˋ�rp�*������������Az���z��\��W����"�7�w}�]{��]�o�1Zd��ݾw0ފ����Kd��G���a��O�����;E���+y�4�OAE�jW"v��Հ��Ý,P���(�^'�ߙw���/n�x����uե�����TVj{��hW��=#W�J�]�t�H��8jȔ�38��h:W��-%�s�>���w
�k4��M��u�#E#'�Υ��\��p�Y�w��)׼�+>~L��5�|s��{_O��~�����ޔ�`��tv�1�a��"�}dܼܽ�u��<Wީ��D��yw�Q�m�U�H��0I��)�}
̔����$��)����?����V����a�Z��ρ��ЁZ��o��9J�8���P#�=�+e�?�-,���ʼ¿���V��5�8��2����7jtO�u��9w��=�Dw��)K��r��C��|�xX�9dِ<BK�|h���E��S��6��	OW��ٕ�~�,&T>Ǆ���)�nT1h?y��~j<�E�����(84�����'�\{����\z�w=D!���}�S�y��q��9S��:�s:~~�\ܦ�<<����ᗵ��,��qx�K�~��)�mS���ZۤmJ�å��'��7�XZbz�&J�sBH�W�(q�q��:��v�<�{\�qN̯�Ӡg�/�&n��|}�BM�\8
�!���_��i�|���z�V�Lr1ն�U
�@+��|�襻�R�J�UZ8�H~�(+�ԫ����Mq����˝O^�ɝ#�
��<K�C�F�N�R֎�z��͇��[�}-(�X�2�G��8k;�`x�-�X�4�a����"z:��F:覎u�n������x8E�d�r~G��__IB�|��M��¾���}J�#fn
x��hh�*l{��UƑ/,�V2ޞT|�י7���N��.�U�	��K���'+[��SC�kä5��s�H6�99����E�[�#kq�ǀ�ʻ�}�%���+&���/0�`�T���K����g2/�-zuaf�G�p�ɝI�~�D6�&ҧn��=�Dou[%d8�b����A'-Y�����i��O'FF&���1�G�qi��MY>K%ۘ��eb�43�����G;�Դ�) 
��T�Ձ���{f�L�^S3�1�����^ٳ����E]�@v�o�l�����L;U������N�uY�3o�_^��<\��ș�?����-�#a�lB��/����Z;�����-��o!�6Э�����|��G���U�Re��6��Cy��=��~�=����x�.�K=�����7��{ Y��o�`�^`�-s�'��+�h�V�w#s�O����&�t`�]���S%��b&�Y�Hf\*�~��x?L�u���CV��V�ʿ��$�
�|���E�ơ{��^JX�i�����/��j�3�a	�����|Whnƭ��7�^��~�\��l�Ա}:������R��G�yv��sg���\+�⒚�2�{��8�{�5�U1ҵT����Q�g�*�܎���0hϺf��0'�v�j4_f3��߉<#�k��.3Y|x�"<�a^	MS���!�%�!���A���&Ψ ��<ǝ���\<B<3�u&.��5�z}�hUT,�b�[{�����Փ�z	��ƶkt�^�L��R�r�s"`����a����������VkcE�U�ɞT�4��F�4�(�-7��P��ʛɋ��#�����M�N'F�9�b=E����iV���O�'�Whd���Rd|��_��o�?{���z�;O���/_��ys���D�	�c��syq�������	��W�Z�S�����r70��N0�㡉���7.���{ոq.#��Pnaa�o,��O�.�kY�Ǜ�A��;��FF��������K>�?�f���niK�U�0��z��M���'(��!D|�!�rr����;�Sv���5����G/p���)�]�#�טa�O�U�/��{�u�z�A|�T��W�i��_�up_�����I/5܆m,�/��&B�y�)���ng�g
hP=T<�A����tU�ӵZ���R��Uap�Wk0�_�e�prm�!�OQ�(b����D�!���̼���NC���ON�]��w��N��H�� �6Xp�W��%1Q������Gk���k�f쭪Z��}���'���朷�#�Ѩ_�Y�5h��;���c&5��å�j�s/�#z~E���r�}�R���إ��L|���R`�_LJ񅓯�4�1�Mΐj��yt�}����'�����u�qH�@f(�2X��x\�� ÇAnhɾr�&\����@9�?��'�2AwG�u�=i�6/���}^b��v(w�p����)#aCX�K��/��lH�A�z��w�~~.��*�se��a��Ov��%��Y��%��\��yO�;?4�t��F\�;#HH�$܇K�G��l�57��5��Dq�[��]�R\|	\ܹᗡ��R�+UXXh.\P����jt�h"mm�X��O�#��R���Y���Yಷ�4�V�N��7��y����
�HLQ��kÔ�s����<sΩ�]k���@O��t�L|@f^|u��{*�@�|����Û�K"��3I;Z��tnd�]iG�HK�~"vX����Yof�V�`��>ãmö�z�o6�3ԛ���|���kl�m���j (8�Dr���-O�9�\�ş����+�}���"������%4*��w�j·�,�jځdu�ų��ś��A��Ė=�3)eͣ�g�@�ҙ�Q�����*nf7�yi"� �	��	=)�F��c2=��T���.a��ͺ{�֬7���z}��������d
:���N9�kM���y�T!9G�a�v�Z"���l�����s��sV��b�[��e�T����7J�	o"R�Q��q�Ғ�l�L����l���p��9�m��cQW�خE�d�C�ʥXe,�&�����1�[�] ��c�ť���1�.������9�G�5��r��<�S���5Bob��\�������G�*h�ؽ���$E�4|g4�|�_���O����W��ZɎ��v5��I����K�5�nM�,.ܤOXV�-�"M�:��K��^im]���oLk6�OѺ&њ�E^]���v
<�����Q�0���8΢���r_�qy�uP�H�E��a�jQ�M�|�ae����Z�ꚠU�<*�}��P�ꓷ���c�p\6�3��$�T�]��1�
&ϵT�������-���y<��-ɞ���<hC���=��l�}8Ԟ������Ps^@����[�E�a�C�c�)�E����+Q*fhQKI鍔�����R�����7`Xˮ����s�	�%�&���W,?���d	��׹}.�y;�|�ʕ�#6����>2�&.���.]�,v����R984ռ3��Ll�U���^h[ZR�8QgӼW���P��`�aJ܄ Ԝw�>Y\�u�D�K�Jj�<X�6s�(E���1�Q�3?;�$�\~��yO��d�C/F��ؾڧ������R\\|�H���{���ĕ����ə���j��V���p��y��]���skf�P�߄�7�x#tu|¾�J���t޼ɕt������}��v���S��r�S.P,�<p�^nۡ��#"ϔ��-Ҿ�5�q���~��+i��+�y=�5��N�K���.~�|��q���dԣ��W5�\zFjM&}��#�[�Ϝ�>�_�s��A��-�����S�(��d3��!��������	Z���K�$[���z87i�:R{(/�&#u����nPL�u��]<�5l��]D�!�U��;��| �v�M��"Gz���u�lY���"�k,P�Γ�e�����\�K�"b$Eu��Ѓ���>�e�xlB�e���z~���ĆϱY��7�:%z�Q�5�5����0�G��Z��H�W��%닪[;��oY[���b� �r��x:�DM��{K��~��tw����-���v7_}�8Q��Z�u	��� )�S�%i�'����3���n�\�~O����(�1�!�[1���"�p=f =��g)�#�8;{�*Ҡ%b]dѽ�K�&��� 4K�oӅ�o�3�<��ڐ�	ҔJt��c��bi	x���0��i�c�QM@E�Zu��hq��ȣ�-����QN�쯳����'g��{{�Б@�bݴ4R}ass�13��X"�G#����=zNC���-X��.{��޼��J0����E����ľ�x]������������.�=}��YX;�u X�����"�U����r��{��jr{�y@��}��"�M����`�*Ҩd\dz�1�V;}�#���mk��P�"Q�B.z�N_��b��,�z�|�u���{��ɣ��\�`/���:i�1c�D���}d���:��Hޑ�?��)��&m�C����
��%�a�ez�cQ�N=PU���W������I ���8}��.���kbRv)�I�:�J-J߼�x��ƙV���~O��w��^�h����ar����[��]���3��\��-��"o���|t6�K�)+��SNy�;NV�FOX���kdW�^a��嘝��8��h���x֛������4r5�G4{{���0.K}�y0
���Dv:��)��6aE���{^.����O(���7zZ���a�Z�h�̗�w�n=K/ȣ�*);�>������Lh�lx`�6�4<j�f�}��^Ł�{"�Y�����S���)>�V�|�2�Ng-���~�?-�1�j	_}5���z�RC
H-R�����3�H�!������\���5�I�ram�$T.$̻ە�	��=�k����2<"��(�`@����<����s��1��"�fQ�<�=P�;���E��+��>s�����q��Y˙�J�+�,`S�fF���>�z)�o���]M�sa������]�:��v$�W�y���̑���;�e�+WF�-����Aq[[���د��`&��>��Ɂ��r+�fҩ�t �ax�qݨ���ˣ$X
�۹�~��[�.5���nk]�e\�.&���.��ԃ쟞#�����gpš㵦�]�^9��4E�����vv�
��%���(/c��d8'֯o�$B��r�M���o�5����܇��� ��	�2��g�:E\	x�^� ���S��;���ۛR�C�t��o�U&��ڥ�:�y��l��mH���Y��|�_�@��w��g ��PU<�R�!D ���Fh���S�醊2DP���]-A�<�~��T�����d�i5P�b�#�:������\P�u�i:�����T�`��J��{6��Q��/��B,,ު�%�y�2ղNrjN�J���f�����G�wD�Q��pA���4So�`pP�J�8M��U���)��x�)x�1�*ٳR�^��pbW�B;@h]M�~�RӇV�\VnGݩj�7������T�fB���FK%����<m૵�@{<23/�:�����9wpȚn��$g=�d<�)Y��PȖ\�&輇��G�I�\�[���Iz1����u�~O��Ga���_u��\V���#���yT�a��^C��Go���ܘZ||2R����t5�;Ӌ!j}���Iɩu7��j$Δ�����h����ڛ����Pvs�������Ռ���Od��l�h\hx�n�%]�yT�4���f����K
L��.L����J#�{e�5F�2�c� ���x�Q �@;߯��9�6���s����9�܉�Ȍ�9���ɓ	�HA��1.�yKI�*C���4�"m6���(@�Α�ƾ~���[�4��ǫU)��86A��K��q���!�ޓU��L/8�2�f�.��ʮ\�b���fȣ�F�ߦa6Y@°���)d|܌�ٺ��ټ���ȵ��qz \�Ih�|�u��1kve��-�8D��W�M���ApH���j �B#1Aw�mU��:�����lSa �e$�1a測J����{���uK�,5oD\�(�NGR��/���c�Ć���Yb�}��4vG�V_�j)�4�ap�U�6(��(����E��|��z~�ީ�����]֧�Ԩ��T�S�ĮlSĔQEg�Q��
��K���*Q<��_��6�>�w�º��V��#�L��������~U�]4M�ʹ������fc"r�_O�ݢ����c������@�������&'��Y����n�N4�h��G6�_c��Q�1K<�ѣ�v��)Ϟ o�E|ջȈ��DB<"������}�Ѹ�����V;TF落3��n�\����V����|Y��Xʨ�[�mZ�0�N1��C���/RԮ���$��mw����o�,�`�� H�l�J�:�XtV�2R�͔���͢fiIՐ0�$��޻w3�N
~X�E	y �^>'�L�����ּY��Z�2u!�g#{ �|W~��y��N?֤%5*ntZ��I�=�{�J,�����/�Yg���Z������Y�󲃆��0��ZT�3��a��(T�Ns�7 �·}s�o�`�純Í��O�����=nlėEX1���m����j˳��" w44�p�����y�f���#x�B[�_q�H���ȉʗ�yϻ��¿QLv���'�@�E���� �x��P�$�/.������8=�C������n�!{' 3)�e���$^�lC3|� om|�gNę5yN��ȑ�G}�G���+^�_:�xQܺ��r������w��Sn��
�®v�_x|�S#�O[�� m!�~l�#��
;z�: �+�����2m
(|�
E���'>�@Ƴ��� B����n��V���7����[��
>�� uu�	Ⱦ��w��Ś3Q��6Н�Ǐ��k�[p�����!{�P)l��n�=U�Q�'�����6�5���1	����D�\حpFFd��N�D�p{�����YA�s�]tr�-�m狁�(<֬��Yp'"Y�k��E����t�K7��h�m��DSsu`���QrA�� !qb��7e���K^cb�
c�ס��f��8���䚨����y�XO�k�D�^c&�$���9g���F��ό�+���J���%���kU
��+Z��G\NzU
�TׯS�pGW{�xyƮ�ﶉe=8X[�N������c����[�ko2�ʔ+6�/�����ơ��A����������Ts���j]AY��P�����M�����V���BX��{�?Υ4-Ш�F8�T��-X�f���ə�W��T<�gZ�u�w,����o��4����R��$L�q��z��U-��W<��!Z�0d����O���JE�B��	��룙r.�����fb����'< R��5��z ��VK�%x���I�ȴ�C�B9@{��؉Ab)Mѥ<Y�a�n�L4�O��ez�̉"�,��&�R�.�[᝝\=L��?UW�)� O��{ ���
�b�r�\��8=�X�B�wm���*�>�G5�8�\�F�B�e�J��	���W�Zo���M���
�J���hn��-n7�����@e]�t��K2�:�s�|�a�3�߀a4����UY�7�]@̯�Ǔ���e���'@�r����e8��]� ?���a���-��YF�Ts���l�t���seSU�D�)���]D�O��Z����;��Y�;S&��.����P.n�g9df���B��A�]>�%Q�!�.��:~�ĭ$"���$��5��ȿ�����6��=4@�[�J{�c0��1���&�֢�!N��t����Y�2��}^��D��Sd���c��m���I����	��m���T������_�X���s�Q31Y.!�E ���^�6/�n*ve�]�W���::e�1�'B��/Rj>ɑ{Pq�aDR���`�r*������a¤e�� �
Z�C�ܹhȳ4�'rh����cdT��%��� 	��vŰdQǒ%^zn�:���۷�k�P�Bñ��DZ�a�zy�Jqy����̀\:x��|qh�Q�a-~B^pqQ���U�*D��ZB�����]�<A<�u,�|�pE�?^�q+��W|���qD��7ؓ���1�����X����U��~��^(����-�5LSĘ���A��̲�_\"��b�)6,J��^�����m������S�O9`!���gY[�zf��,&˩����+S�ri���wv�h��q%�~�T9Qz�ʕ�]�g��V�7i�um7T�&��R�~���������/h�F�܀���΢ �o�`©��G� ��3c�3��^�S���D­Qp���&�/��x�e��&"f��u	=^Xx@�P��x��-ډ��/�.�������Ve�����d�
^��:�����"��Qin����/G
�X�1��"�	���&)��زo��o�c:F���yq��߿O=�_�c���vC'|.�l��5�.�ދ������xmYD�[��󘘹 �*��K�L�jγy��_�����#q�*����}?�:��g�e�p�$v�A���!^��6��4��Oz"���d�Ix����6��'q���5Va��U�E��Z���\�m�4b��&��˲�&����Ӳ[��z���R�6��1�$3�O>�J \F.75?x��)�ۭR!�D��9bΆ��G@k��G��������˜ �~�⪎;O}}U#�FuX�S��w��kI�26�H��~".�X����ѥ�.�1�/hE�B��
��?O��xd�Z��X�Q%�������!۶m_��n l���f{zĆ���ę/�0 h�xM�.�*���/��c��$j��2�Dap�k�Y�T��J��~=�Dn��d�E�R��b��o�.zC۲Uk,'�J�*�o)\qH%v��C�(����b]s�.��M �p}�+��~��§�=��ɋUV�@�qL6�Y\ Pʌ_�"�CfV�@�k]����]�r'n����~�=�]QVAR�޽��;���	|��������rZؠ���"b��\��݊��5Pm�::��e�p���!�r�+o�����L��m�{#�(�5�A��~��K_�0���AY��,��F *���=��<�0 ��{=��ň<�x�c�W�5k��?�M:K�(�Bg�8@��F$�gέy;z� �	�M_�Lk :�����ΕkRLP@rg@e�rF�	��?T�[�(l���Oqp�@>�M3+�iC����%%�=�o�,�ۖڠ��uӭ���1_��8GiZb~���E�q>U�q�Xݑ�y�ö���ӡ#�f��U�o��AgW���Q�A��9ݰ�ػ��ؑ8�R��+�=�'Z!R�d����!�n����
 1J���F���p��}��<���mD���hf�����_��
(��GO�]�ӿ'-��<l��#�~�VR�p�	���0��N��s�ѠjT+��f�j|���[�<�g�Z�T"b��d��o3�`Kl0��P�Ȉ��q�;�:�p��5t��X�
�������D�lU�m�ʕ��L�咁3��^kŀV�_H�%�����ߗ��=��
�W5��ԧ:T4�#�Rk��|��)���I�z��W�F�e/Eea�;����Ɉ
5���Abު~S�� �![������U`4��a4�~��a��á���aZx*K=��Y��"{�}(�2�}/�E(D���}3B��o���e0��0�{��������Q�!�����:��s�78���XO�� o�k��&�m�L�&%�bx��E@
LO�2��S�>��e��*�`*N�p,g�*���X�	����NWY�|m3x��K�8�:k�Y�2k�W>c��K����Yn.���r�e����_]\- 8g�lZ�l�rY��f��DP�ŗ<�T�!�7�j@��S��?+p��E��4�}�<��c�&��C;�Oޚ�L�w�u�����Ty�d�a<�B�mAD��z���bO��{�dW���75�fDOE��Z�,��S�>*r[R>��G�I�̟-��;6�j�,D��Ƈ�?�kUA���/5N܈ɛI�CyF�4i���W@x������rv�N�DT���S�v��u�?#�?K���˿y��\�c�/�0�mO�{��Ŭ2GhmO؅�xTp��*I�ꪫ�J'�߿-J�x`l�
�y���CR��xT�_���H��2ۑ��w�=]d��VW����5�Ɨp0����������D�.}��:~�;cj�D�jA����!2�4�;z�ZW0�./�����&ݱ,�(��N'
&�Ty�нfr/ h���P�\��u�$���ð�������l ,�k���6rŤ�M�:�A�h���V�&}S2
�Oň�L�~�67�ܙ��&{���&.�k@��A&Z
e�\;W�g��}�M�}�*�O�z�4��'ގ�Y�;�e{O-�x��<�Fl+�;�\�l��q���M֜���rl{q��>��<Ϊ�lm���^���T��x��Z[���сfǇ(�;딡��Q��<����~a����S�녪�_�o���v���QS�>;�c}f �N�_��(<�wQ��2���4��S��gO���4�|6�N�jffS���Ӗ�� j��P������O���H(�aiDۻ^{��'�v)�rax��� ��g;�@<����ɤ�-�ų1��:���D��gӍNdp�2��FP��y����~����{-��t������Ys�
M?Pb�
4%��+Fi���� ������u��S��ޑVD{c<v����RHQe�N~��]�`�Fhh	 �4����W�����"'g�G�T: )M��� ��۞.k\@��z�����˕!G9Xz:��-�����`��P2��8������uۿ3}�;��C/V�;Q0l6�
%m_����4�����i��y�l�_��MY@�O��L%U(jk��f��ƪDH� �E&w���k�τ��y�$	��/e��!��$�;`���ߌi�}h7��bk��2d'�����Degd�M	=u�����~`|l��k��%MsI�:2��^��R���b�]�>��@�{ÿ���*&nyHc�1<�;f�����3�w�p&
G��<��gަ�ol\�#��'o~�[��B����p>�]�WL�觷eU-*��{��V-��8�7q���HĖZ�o�oZ5�1��"��b��·1$� G7����b�S�b��~k=&�fgh����튏�� ��}]*����ae���C��fӸ� ؝ǆG���Uhpp'�udqh���|*��EH2�Jum���n��H+�v�	qf�G^N�]�n�c#�\-�=�/�e���J�x�Ke�t��ŋ�=8['��{����1AP���R���P�F({�\�$ef�B��j�*�֩����n�$>ȟ�y�^��A�����qk:�������N9�7������-AB�]�����o+�mY\�12+s���RGJh��a"{�_�"�5�t�_k|��mQ��м�������"�P���j�>�L��'/_�Q�5�v�����L��t�}�E����`q������p�~�#�T�K0�s�P6�]?i���_�[g�e�m�	|ۍw!ݧD�a0�j��3tc�������+�Ҷ�3RXq��@i?K�����B�;�Kp@ArcżMZ�ٵM5�Li�l״:�M���OI�^M
ˤ�%/�]�6�;���c����h�����U=��k|��|o��Bت �8Y�Q�ȝ�9w9��Ot?�������f���L��=���2���u��WP�C�fs��S�t�	+���4)�A�ȟ=���N���? ��ޯ�đ�|S;XAp`E薝�^��h�����6��6d|z����"��sh�'	�C`<�Ic�z��[���:�J�7�����e�@.���fגʡ'Ul��~n�m�a�T���!��8s����5÷ww�Cl.L���3�~�̍�֝���"����Ɠ)�M��ĝ�}4�g1�ΟB������k+s/l�����,U4+��Г
(;����go\,dC}��JkfϽ�2��x�c0��u�Z!����}��לۑ�q��N�}$�@n��9q��&��f0Wkg4�&�d� Hjʞ̱ޭ�g�:�U���#x�R�b�@R�_�boL;E=3�}_���q��z������a$�k�����;�J�]$h�,�}��/,s������,¡h}��im��h�Q�E��##uzXD�SV�C<� �����{�K�
�B��G�v���pTp�~(vA�~'����V:���� �H�-[�
���K$\RD4]G3��i)���I*�9v^����V&l;eӨ\�P�N���,���W�����̱��w3�ȇ&>�D��Tj�{�_��es���8ʽrLɨ�@����5�7fN����ߧ�Z�c���.���{�YwřW�D�_��z"?x�o|��:k����T�{1�1quU����
�t�t�Ůkw�ô\�2 %�����"G�D(Y|f��\�-x	����L�7�Y#�����nH�}�����7�u�NO�?ɦ���n.�n�GX��|��?�+|CH�.�帕8n5o��#��xaҤ0���h�Z,`NG��6i �~K��ȱk���,���Wp$��[;�if�;�'�㻵y��ˋ��T9�O�n��Uy�\�/I�q�7�7#��~x'-q_� �������� mP��z̀tO�P�a=@�+m��%Q/;E�仚�uG�%)q*a�+�����|�WگAu���V�52�~~,J(����m��Z�8��y�Z��w�%�DD�����`���bP��ڏ^�#��LXS�bC*��(S}�{��Z��-�aPЭ�{<5HV�<���?��YE�l�ՠ�߰������q����p'+�~3��&�u�`��w�y�?�:��M�9��"���g�:�r��2i.���qB��(/kq	>
Zm?G��>S\ e��#ݗ��Q4�����P�H
&/�}W�ﱾm�g�F�}X��� x�+Ic�Ј� q �y�J����M���Џ��1A�C���'�f���@�i�5�{U�I�谥�K�>h��#%��7VP�_���4KͰ�^{�Dܘk�gꬫ��4#��5�/I|-~�pLkn�K�������u;Pt�>�p=q�^Xj���	叙���|���fr}�4X*�w�x/3f��=[�q��ȷ��
��#H�7���������b�[�O�ǩ�/e,�MC�Ǳ2���\�c�ᔂ�����U0 �"��۷�mc�pd�ww��x�O�CΔ9�y�#���⩍1s��B��U��n`ڕ'm��G�����;�ܮ��
3����4������vW�s�Q0�0?}Y�9t~Z� ��
^�	��Zi�PU!��0;�e >������I�s�E���4[���z˟��C��=Ȇ4�|;��t���V���� �=}��X�3"9��X���)x�@�B��'��T��\�e�^w6mfȰI�ӠfJ���ɺ��?@"D��Ġ�����c""FֻC}l;B�7�� �S￀��(�U|��oc(I���1���j���b���-%oqN����sCby���war TJs�f���}�E�wG�wu-��+`�u#6	�p=� SU�.u��Ӱ[�d��=��<GF��矚�8>̿'�Ř~�3����5ϖ_C`33�3�*���b)�c���;��U�ܮ�b@60ݽ�wD,�T̎�nE7r�:����v�v�Дs�ݪ�R}Z3��9Ȇ����t3���E#���&UA�R�F �(z|�7"�$��C#�C��0;?�	K����uo0~�jvwp��$4~ob��u����q_�p#�.7o~9�V�9�8������O2샚Z94�Ld��x�m�L*�C[��.b1㍂P�i���5?SO~����x��u~������D��^a ��}�*zЬ�j$�Tu���C¤��4E����̃���6�-dF7.��p�;�]��0�;uH�xT�	?��Q�j!�EF`��!�5B����aoy�y�5��%o����llk��
���GJ��{�p��lLk�����y���yk�P�JL�CI�2u3��4�k3<���}�({:nn�?��s�+�����v��Ĉ�/9EE:��9�i�ن
wCj�ω�L�t��?��^OHw�z��7��QA�N_�!���k�Ǵ�@���
�24��c�á:�@�$�
����VЀ�3�J�V��\�ez>�gyk�ʊ��h3WT�
�Nb���۲-��
 ��#��tԝ�!�H˫$�U婲���IO4X��Cx��_���jj�@7�
���C���� �.� u1��+��I?ː�;5�,d2��w^���?��P���d��ٽ��L�?��;U�I��Z��5TB�a�Um*�LgU@W��.H�cr�M|��K��"��d���ʸ�^�8۔�l�0Ɗ�'wH��pEuyt�cQ�̙㇯VQ��j:p0UG���3[c�Rd�������H|�ډ��v�g�݇�'��3����!�TE��Hl�������(y�߳��}�� �a<R��ν��&E�!�&>�s���iC�����T�c?ji8��x�S��ϔp��-a�[0�#⯥�&�t�H|�KM�����w%�l��E[!2~�bj χ^��_�x!͐q9�Dߓ�B-�ŋ����r��Պ����^=��\����A�CJ��FW��Ə�P�~�������/V����K,�
0"��]�:/ӻoG]5���Jy=��9y�~�\�v
���)����%dc1@t@��=Z��������oC᫫�z�3Cp���6h"Β���=#�Ʀ���P�;]=±�1y���ݹ͍f�,�n��akF�juP�~n�;���{��T||�"�>�:��:��V�H9�s��גf�oJ�|�޻��^��8���D{u浉���zu!��f��9��r>O��\��fǪ��cSq��V ���*�o1�nN��;@# �v�y�!U��1ШÖE�G���L�9���O|=T,V��(��"Cu���{M�ki��o��I�ܓ�H�ij��K
R��_���U1ij�Zy�N=�7��X:�}��u���C�&��P��ZbMC�a���v�f�{�|������@w���)��$3�������G�P�;rȏ��l��;�����]됤$n��r4XH��p�3 �ENh�S�����5V�N9+!^��u3�=wb���+��3��l$m� �/����f����Mq�M�"T�O�Z+�/�?�T�<d�i���ᤜ��Լ��S �V���lBJ�#�s��"�W�h�,ƹo3Ɔg��/�*�=�$O3��wmV�ZQ��rdo5S��31�����P�H]�n�fE��Ԙ:Pzz!���[�=b+M��+G�c>�
���L���1v+5߽��R�����I�Y���7 ��2Y�g��RU0vw��q�{@�4����IO� %u���90�������k
�9����_��D65X�b=W��~`"z����
�J�-��;wF�D��U<$Wޫ������?~-�r��9�0~,[T��I�>�B����~��ØLy<�v.O��3� м�``�$i?��(�����9a"k$Ƣ��;��/�%���(�2k<�g�!ݽ����$��k8��!.ZI���t_ۼw���Os�]j�爖��ȗ-`K��#��@��83).}lM:ġB ���&���P����+g��jJ_n��y�[�{���XZ�l
vJ���*�^.y���޹�[����}x]FJ
CT��rb�zu�q�tl��X�4����axȯ2�N�{�������2�E~��Q�)��p��e}̼��q`��e��ߚ�AM\)W�՗�%o��B���ڮ�>�E�Q�5��*�&"lt���*����=�����bD�5��襗^!c��a���M�2&�i]�#2��P���}޽�3�8�/�z������P���&Eh�F`h�{��z�;���aQ��v|����͋�t�B�j�����g�*
��5�h͡6w����{�ldRi���Z8����R��C��ۙ���������y��q�U��=�D�[�kg����/��C�M��D���F�@��m�X��T��`I訉�P7�I&��z�ҩNz����4B9M`�s�4r��Ft�w��Q���{w�3M���p���]ٝth�v?���M�#�O}���I����|���B�R��o�<�M�w:y^!��f���`��m�ob������M���(�׿���ļ�.0�sS�l `V���N��R�|tm�v�����xGSh�pA�J�@+
�Bj*b^g퇦�:��T���ψ�;$5ؾ47H4�*�����wm]��X�kl�w�U��{�7�����Yn�E��a�!ԇ�e�З3YM���^��s��-ڶ(θԷ|�,D&gd�K(@�����g$13�-�H˛dQ�>���vm]D�x{�����JV$���/�Nf�!G�:e�FC���p('���W�C'5�Ę��m���+�!Ƚ^=�sa�f���N��a�JSG��80H�QN�.iK���^16=�i�^�F^lye�K��8��Q�n�W�d_W8}���Ő��X��-K�x·'p�^a���0�>�W^om/��k^�����(�������m,��T�LޣG�:+�]��B��v���x.��h�R+8p�E�74c�<�(B��p����&N���F�D�4iH�<���?�q�=^⣝���L��I[qo��<��ՋW�j���j�%�0�d���[u)%S��;�M�l��V���FUA�_�W�!EJ�1Hw̓������K�`ZKӒ��~G~��1R��K�A�X��I[���\V�A�!���Mii�I�K,#�"�����{�!�̒z�o�9�*Z<������.��)sx u5d/�u׹�i���R��yk�9�!���bK>t���>���i 0d>z{���7Lv��W� ;@+�fEpS�tuM�a���
V�o{�|���s.����y�ʅ���w��y@��m|N8�h�~#6�Kj��uA��F�}O��se�)�[������qAu��ZumU;K�'�^����i��fU�a�����W�8�����sf���!	����������>D���46��};�R�rNfK��= R�$"�"( >kw��g؋���^���2-k�Z���ʵ�x�G?vq?X��9�∼aL�r��J���Z�W/��s�Q�	kSy�V��H���ؔ6��4[�?�U��l�۫��a������Tb��x�\/;Jٽѫ�zd�7�p��A�|�E��,���[�V
�W/\(X&�v:�}�,�/j�X�x�r|�X�E~�:r�Io^���[�e�:�^����NU�=��>Z��B<2:�tѝ�M�KL�y���E{V��J�u��HJn�������Eہ�ir}z�7�h�t�q�_�[�VY)ۛ�#Y&Lk�i�D��������U5��;�����4�Ë����Ȩ���]W��e������y�x��njU��N��b�{KD%�Bʌ�u�u>y�����r,�2�;�����t���й��}�������dM�k�zJ��A/����
��ऻ�+�f'�� �(�P�]���`������{}��?�[�|�<H#"���^'?n/I}�����Z2%d*�'oov�{!�v�D���FT�w澳I�����E��@�����ctI����S�y�Fs�&b�>��b������Ԓ���h�h�|�)�B���&���q�=���S���hT5����Oy�&>��ph3w��;�8e�������~c+��B]��������%��s��X�Gk_ȓh&����Q���b���-�<�H�7�ٰ�*�^]0�k��VXp/�XF�p%Q��:�A� 
-��bd������_7��[��F?/��# �856�i�i��R��񣯖���3�?��(�M��~0��טT��9�'���s-���+��q���$��>�qSo@m��yh�Zͤ�����NXӣ���Ub;\R3��|��߮�L��<�踼��U#yO/����U�1�/��	;���Օ��o;�*ήL�h�Ĩ,�$���5B�|*M2�Ɵq�e�pq�RK�L��!=`g�~� �Rp
�z�JP��siJ|h�P�yV7����p.5���N�>�L������h�F�؈K�
��c1����a7 �ow�Ư<s�z�ho�U���z�Ӡ�>6����v�Cm)y�,ŝ2���q�!�G��/l�����;�%��j�|W�d]��Pߙ{�=ڱ �ypu�蹮�k��^9�ZP �h��#�x3O�����AJ��'��m�$�7F���.�����4�7�t�/e��ʽ{F���� ��$k���;M��=No�G�]����i}`�[�I\����{(��qvS`*�
y��Lj��fq�vN��|�����K�m���n������P�:F��� ���c ��G�$� �!��F���=-�5�:��n��A����&��0��,�����>b��s�3���D�!�-&2R�Ág`��%�!T��ind�����Ýka�*�G0��	�U���� a+��N���Ύ�mD#	�*��䉚S�<��B�!�3F}�q���y������p�TF:�����u�N
�B�&�[A�
'U\��2�*{�$�e��������j񎀅M&7��n?[Q�c�p��~:�~n��U�;�q�����'�G���2c��g�?o�X�Aפ�?�[��W�!ȼ�ًkLI*��lݛ��A=��z|��ܔKM7F,�#*��1qcb=�.��ÄDr:�a��>�1١�N���ω��Ճ�L��Y���r��M���!	TU����߸�K��j,�E��9�k�y|A��~PFBΤp?�%ΐ�HC���@��A�}�,��O{6�no�Y�O��)�zF/�d���;���$�Q���d�(-��{z:#k�VxLz��u�HI�K�� �z��J ��\�ϕ��E�nY�t,+\G�cq�F` �.\({/<Zrh0�u��&�H����)C}�G�&s�k�oy;��MM![[̭?ݕ���P�':@㷱��neP ��1*�-�۱}�_~����5naaq4�X�Vٖe"���Q9@�C�
#����8��p2��qY%o��_��Ϯ��ޒ�J������C��5������Ǥ���we���*����Tk�Gc�*�CR����|1�6j�K��&p�7�%h�<�y�̒�+"h���t�|�ke��'^^�!���b��+�x-���r�Ν�Wn@�Cm�p����۶84�^��zw�S�[��̴z�&9v<9`P�����Rؙ�nv��O�����W�B�=�4{�c^��y��gU֙�8��1��y��#J���w�Pլ�h��C'�=�����l�#�u,b�kJr�o�����A�� �֍ז:�[ZzW���3҉�YQ��o��C�!Q�k���~�po�1��|�V#aZPP �qv�����yҍc�~��[^fQ��y\����ů� ~�JPT�3G�0-���H��Y��+%ջq��i��M����]����5����$:0�;k;�ʠ%�������}!�����kwr���m�H�|:�m~���������p�c�̱�w�L�Ҍr����?d\�I*��L������N5'�����MJbq�s��4
�_jT���٦�f������!|���iF����ͷ��D�����D�ND�cSC9OM���	���2�)��]���M�F�Q�d�:��xh���M�+]��9u��`����0]�|�5y�z��� ��bþ�L&�'"nפ�V�d�K�,�MK�m�����D�R���z�ӰI�u�1_}�<;<DHh9�D��x��F�E|�7�k.�ÉrN!�$�X�oQi,j�8x�D��L�g��z0�Ơ��婊4�t�*������Is�ψ�x����E�[Sc 	Cb��������SB�o�`}�J>y�;K�~��\젠Z��AppH:�B�2����*��5�I��K3Z�UnN�?(1��5���,T��aa I�KB�/�UiY����Y �ف)�r�m�b�	��J�`�H�k��߷y=�V��@���=���/�aoY���
Tۥf�w$��.qi�B�Vؕ��R��f�oT����O_|!㦓b�a��=׆�Q>��*��[/���:�ͭ�-y��F���^�5=���M[��@; 7W�X8E���_����I%=��?(��zg7���{Ԧ )�	!��Ǐ�DC��[	�/�,��yt�v��'���5hBlg�����ŖA=!�/��ě� W�E�N�	$��}t�~UY��0o�}aaf�P�j��^�:B�:��rѥ5�/��줎����
_���E�l �G;,��XD�E�W;�
xp�(_3�i�-G�	$�hN�Q� D)���
6-SAw;����� ������Cs�VD�v~~/��})�8���`���贬�{>��5�כ�i���U*P�{�'Y�تI���*�S�$%�^~�/��G�F�G���GӶ�3/����]E#c����Bqݶ���g\R���~_C�;��Υ���`_ A�#w���۸�\C���%X�8_���J���廄@m�#�S�v�q�k@%��RkB\|�{�Q�u,��d˻�>ʍ����7;�
����$��_CauC��m����qE����Jl��լls.����+O�Mۗ6� �@	UtI�L�|� ���BE�P.Ο_�����N8�Q���Ӡl����-�z$?o�Q�ӣEk=�R��x���>;�)~�<~yYzGD�i��>�8J2���w�j?�=��P�q��4;G�M�޹��� �K;�� �m����	��b# ��=N7f�Qr������K �l��~D����_��.Eǅa��c� t_�5�	��x1>}4�[Q	�f�YS��1�v���+�"|�2��)V�
dbq����ؽ��+����uz��v�uُ�z��=��@A���9�����G�S�^�:��[&�H����oCC���c�s2hGy[g�ֶz�����2�(ih��w'�}c��e�3���nv���s܄e .CM�@�4����&]���0�e�6O�=���*����F���ßG��66���U��C#�aЙn}��k,�o�F�ݺJu9"7���]���M��C&@�KGL^ "�uv���d'�9�%&*�N�M����fY}�+�(���8Y�����n��R�X\��V�CCL�Z�~��L��KaӼ�e��g���I�O����
�ZE�'�R�h��,`5RS��*�M�����;@� �VaP<a���[qq$i��u���7O/~���d9�zbM)�&]�Iͤ{�qz/fP�^8\xs֛�ށ���nm���Je|��h�(AI�ʔ�0��ݬ���`#$C�Q�~B�y|<`�!?�xTT0�Z�{23&#N,���ϲR.��( ;�\6��3=�]���~��A�X��=D���Ό�CA���C[D��,�<���S�����.�E�9 ���������u�r�~_\)�ʀ�= �lx���1�_#S[�~�0�|�C��H�����z�?bQ߶�W2m5�nK�{u��.�j����|���.��ʎ<�A!<402�O��آ�����V]v<���O��*���PS��]��ςE{r��[
u'KJ!ם� � x ��Y�<���i<����낄��g��A;�{�G��@UG����;nK޲�d�ֻ4e@z��Wҳ�-���k����D݊�,2����0�/�h�%N2�4k��~g�&����~���v�[��� ��<4tttJ0�F#�,�HYT�W+x�WalPkpo�Ъ����Q��f�x5�f�Sj,��c�eBŵ��"F����&C{S�K��,E��8�ךu��5�4x>k����:�v��K���k_���rc�e0K�ed��w�9Xrt_\�ow���-Y"r�rݞ�]�#�(�y
w=gޣ-
�S@|�hJ�j:�������ꀐ������.\��q�����Ş��+�YΟ}���QlR6��󪣎b�5C�Ǻ����2����z�ed=��4�c�˒yi�M�G��R�g�m_���pI�^1�'���S��^�U^��.s�7�"N)D�j
���
�yr�$�^�L��g�BaD�y,�O����y�d5�f$�RR�̑���<�f�:��C^�V\��0���!��1�Tϻ!�5a�~�I�wM@�G��_M���4��-Й�=
�������7�м�ޫ��!���n����xD�8����=;[��B�?�����'(�b��������
��-.��žL�h�"�Z䰿���d�~�Qkk5�E�|%�v���n�D5��ߋ���\�ݟQ�r
`H3Vof�>O�H����ä�B�I6��]����ژ�mž�Zh��i%� 2Ұy���7��?��͋|��2���e���FX7V�S��oy1���N��s�ԯ8AV�n����4�o�9�BF�9�o�|./���:��z�	<��=3z���|S��hN�����Q�Vm����`U�FHo�U��M��O���	=CC$�:]�*u�D{k;���cJZV�tӘX��U�-�TQSb�	�,4�aa6fۂ7H�=�L5��4�y�t����IVGW�͛�c=(��u�] �иIL6U""ǝ�@�ӭ6���j,2"]����'b��Y��gi�����^�`���-cf�����ɐ��[�d����XN��K�&��F�y��D��[��F�Ai��c��@��`{�DV�{ש
@.�߷x�������Y�M�*�:��/��Kq��@�Wi��^Be�L\jV�WQ�?9�̡�@V�,�ݸo���!�p����'����#^��m�
Y�'Ԉb��0������dOY��x]˚�f8��'.�����.�٥���[����w�M��\���X�A@YgO����,�ʨ�R�tqsE7نC��� �r�xu��5O�s�`�nI�<�l"Y�! ]�"w��������9z'�cQ0/PQ��_��l;��o�q�I��
e�H�/+ǻ����c�p4�lwT+��\�E�W�j)�ظI�nN�Tkm��o����v�އ�m6j�KG�S�g��.��3���T��>���A�y
?���Ϫ0�TC؟�D6<voOEC� j&��`T�ɏu#�29�ؔF��W���/�����_��/�'2���i��?���m�G9�I�.%&�#�7���Q�I�� �c��]B]�[L�6�g�F��-2+u�����z��I_4�1�t樛�R�?Z���2������A�PY�1*�W�{`�Uj^<ꮤt�a��j2ZD���`P�x6
�8ܡY��'��m��6�C���V	X� ��yb�	S C,/᣻�Ӯ��YB��ܪWB��Y��g��V�]�Z�1HU�.5��)z�3�I�r6�]���,���l�aH�R���o��}��n�ph��������L���}�`����Ȥ�-b�j-��w�yX�cM�@R�%� �F�6�,9��)�|�lt�"J;��w�qz	�Z�.��V+5�)�(�`Q����q��7�NI'1���$1�C>ZN�����]�������	
ӊm�{����E�!���g�i��,��\�X�X�l���Pk{�"��i������!��nP��}\���������M��+��S4p=r�c�7����A���7�;'����T���q�!�!�E�L'&���'�&�7b���=��� ���r�"(��;'MkF��i��;�~W�o�,���gQ��S�Hn����M.H,/T?��"���gf�S������v�%��y��J�}z�NU{��K>d��!�ݾ�O����7)]]��L���$OU���[~��C�b��r�Ƅ�f9.��˧:)/���"+K�wR\U=.{��>�&h�F�`�m��{������<��z=0�Z|w�)��s=����G����-���6 �<҄���@����E�R�<����B��W��Qr���K�C�N-��ېe챾)����������k%�Xi/u�T]��O0�_eU��+o�ZqM0�=�z�>��ș�-k:��T9,��R��
���uZ�.�l�:u%U��
Bu��>�<K�pU]�#�S��o7�|�f�S�os���b}�3����~xeT�7D��j�Y} �>#|${޾{g ѕ����IA[�/bT����ڸ��j�յ9�����N�,(gL��w�o8�/������'	����pX�F˛
0�N<�ϰ�N�/K�����;:���o�����-u�MJj�:
�}'��M����`�^�n��Aw�P?KFb�d��8��)�����6��z��~����bfn�8���<� ��&�A��DJ��[4�o��y�6�R�� s�����<�ʷ��]��s$a�S����㍕L�7pm��ɛ�C��ٻ$L-,�D��*O?3��Ԇ����� sq��9&&D{F��w[&�I���3;�g@���.1T���V��}�����h���Sa}�楅1�������ENw��|<]��Q�7L��
AJ�=�ب[�(qO�4�ʋ9\�Z1���r=&�C��/�$N�IΦn��.p��ڱ�*=��w �#�oX1Tc����a�b�՝��C|afS�St:d�-+q�0�o��;-�{�2o�Ov���T���j��Uƿ�5愷�T0+��4�0���Q��/���S�d��;�����[������g��`o��d�Z����n��k�s��i��]����s�n���,�i?M���E�_��=P�OFA�2�P>�ԍ���<m�gd�e�6��ࣽomZk��~W�[]\��{���d�OJ��?�Z|�_뮉��ά��<E��r��{�7����{o�B���K�]z��53��wnݸa0˽+�|g[�sc|�����x��M[�����z.��=άx��ue@�9�/{T���
��k5Em�9E�$b0_���� Z��Y|��2/P����xb,�T@�;[���K]���zi.ΟGZ���<�:F08%8���׺Ό�6�6��T[!�E��/�u*Q��aM���%�6�I��1qӾp~�fS�����/�����H7O|��P�P6���l�Gn���2����E����凧V&S���?%�E��:up��<{��bj������U��%�D�ƍFn�br�l��]�c���[�W��L�eA�L�v���|���;�ګ�:P�����-e�a�0^+_� <����m�r�ù���U6���I�K����U��Q'X12��p��M]�6lQѴ}�0ҝ����]>�FQ1�8����B�4=Y��p~⇊ aPl���o/�e�>g.��_�e�7�rW��n�Mh=#�<)%{6�M�G����D��&h��gs��3�_��(_�^��&�:;0]��mR$x��Ҳ��?j��;�t��?[��Y�4�<0:�L�Ϳ�V��VG->^.�P�H"GE���z����շC��l�p��xJ<@ԝT���w��Sb�W��<I�;<��ň��o���δ�SХM ��k�	��<��:)~��^Z���nK���;ik�
0�7)Y��2�6�J������X��{��2Չ��W�C�utMS�����׹�����o��Y�s��u.p�7"��5R~���k�k.��{w.;,t�OQ��C��5��ѷhxȃJ;8��MNjq�4K5Ť)��̚�=�T��N�w��vF�~X\Ժ�~23mX
��(�L*���-���N���˝S*6q��|������Ȋ�pj-g#��<�q��C	��glP:3魽���w���<�{L���I��{V��?G�O����k�$
0��>sI��1�ʭ�6.�- �s{k?��������y��	�?��#���S�H�]�ަ��P�y6���ϫ``�p��T�c���M!\5#Ęн.e}�|���MH"�t�ğTq(ú��7�.~&6*��4[�Q{pS���]]H]R&���5��kΩc�^���� �}���c��m+Ҟ��������&�b+�m9	��:3��"���X����(	����]S�! ŀ��Q�IOf*=�0��<�}��_u�v"A���L9�5���5�J�	����}�#����& uT����Uؔ֡�ݔcm��\-��p(0���
-�����Rw������%�D��^��y���skZj�t��*�VM�0�8�k	�Ev�RY�C�t�YQp|܎���	6n���l�{��Z�W~��xX��ҳ�}�ze�t�������3�T�O���>N)��'�Ⱗ%9�@���|���4�ũ�N��eVn��UqG�����`|�;�XdLL�>�.�c��*O�r�����<��\�qm��&�
T�t�!Q�8]6Ä4$�Ph\�V�J�>�S��|z0���E�v�r/l�`���o�=� ��bnN|	��ϧ(z�~�2��'	�h���VhH�����^7��B �bP����I�b����+�9�[w�8��7�(��iyg�N*��U\ƚ�'Mi�ʲ�̸����	S�Ǚ,i�laq�%%�-�
_񌲕� �%[_�K���g�Zv���=d
b������y ��%AA:����U���ޕ���umN��N)zZ���^Q-b�����<�Uj֣!��iUUMG� �5ϡ�Y�Xb��H��T�|����~?�?���+�˵�~�Z������_�x5��{Q�S轳����Te�s����gʳ;�@�u�J��\��V�Jx��՚?S<캕�ԙ���UW�/��y;�cOE�t�3���h��U��.~m�ɧ�s�HIYN|h�y_ވ��<�����Р��2+��.�|l+��Ess��6j���M��*�5�z�%e�6��j v$B�[&	c�K�i~0�6n]埠k�	�3�)1��Z$� ]��p���f(����U��A��uri�P�m'�LRy�����Jd7.?��������L��୨��̀�F��c�~�r4¾!�h���|Zl�.	0�Ý�O@rҰos!l�����~���cQ�^�ͮEG�(	�
E��v{n��2�C�M��|��D_���TG�?�F<4��ws v[��2�4�G�,��KHg�m�~o��$J5��Ԛ4 �el�*s�Ǆ��A�$�}|��Nk�~�vҀK�F�؈8��	�����;E���Į�F������݅��X��u��gyJl_�S2���"�Y�R>�#p������#O�;��	p@&+H��ܴ��&�/�����_�ƿ��b�4�w=��Xzc��V��E�k��P2�d��*��A[N�%��Lx��ô܏+���{�$��2���>�������^�p �;�p(g=�����Y���/ ��P.7A$�[���17bQc��9��ףۗ3�h���?cQ�T~7	ʲ����t�0jf[7�����@k�px�N����M��]-��~0?���lCQ�D�����4�S ��Y6u
�f܀��Q\n�Ex�?������v}gj�X|Nt��ޡY����t��6�2�D�ԞT)�&b*"��}�n��*w�L°4�b9���IW�Y��������	pE=�F&����ҋ6	��D��vW{�)5{<ڠ�P������tR�����7wH�P�/����yj�*���Z�#>�LV�j�:��L�������k�'z{�D��3R�$B0�Ğ?��Oh�ع�G����f��9ێ&����V׶����U�MY`�nO�u�*���Uwܾ�^�/��z�?�f�����P{{��ftF��:��"��mԺatY7d.,��u�Q5�G�{�m9A�H}iJ��*޽{���U&?��>��3Z��c�鹋Ρ�v9LwֶU5	e[���(T^p�ߵ�=���z?�B���\<[�!*�P�
�e+K4� �(�|;2'#�>�:"_VS�+3rr�ij?�{}�]q��3~j؟�R9\f�x�]��^�X5ѩ#�H&�\�Y��F��:υI&{�>؛�\��ý?�<�$-���v�N׺�nXF-�Z��J�(X���B$P;�ؔ��!OV�K05��U��7��.�#���w�An��l>f[����`7��Qr#��S�T)z]'t:@�q��<߲�L:ֳ�f���pℂ.0<�}~�+�[TN��I����5l�>e����K�sؿm�;�H� � �����k��ײ��`����)���*d�9;���k��NI�������o.%�~$����|�,���i�7kcnp��=���pڬ>�K��]�%uwM���8��7�{L�鬃4&��t�������bԈ}F��>���Å ƠC�ހx(�䴃��T��1Uq�O� 5j]v;�\v4{��υ���6z���\��蚕�jZ�����O�����p�St=�\.���3�e�?͠���V�<	�����H��-	 �*��F�Ei����\�s�����4SA�3�>��@LL����*g��V1 �+��0#p�K��鉷���~��b5��薿�x.�Ɋ��P!3��U#��π����+��~=?u9�W�����F���u�ȑ�B��BD_<�!1v��>^�63xn䌌]M;��?���,��wd�Q��T�G�z�s��٨~�(M��'�XUP@,�S>�z0g"}d5um���[��E	���6�;�[�5ׂ��A=9X��n�v1��Z�w��{I�˗�>>�^��K_-6��Ȋ�S���Qq�-��G�f��F2l�砿*��HS>)��nOLd�"��a�LV���B�"��q"D<[�8������K�Y�\�.S4���ϧ�8��������e�lҸ~�Aljj����lm�\dro}JI��y�u�l���T�sE..��=�7���h�p؏�����_��������!-��P�W�|#����(��#~ma�bksu�-�*��Ϧ�v~��c�n�y��l&eɕ3<8�d��u����U��.���-�SY��:NQO������ztkPݸ��;\A:��s<�u*�BF��������zt������ݸjd�Sߐ���bqR��Ѽ��?�pV6�5��mߡ�P��}e)�T]^�5�t���z�EG�c�zo�	q�F7��Ҝ�,_�Z��z�z��
�<�� ��[�j ���b~\�6���ٯ���L,^���'����ʣ��{p��k��B�w��bc�j��D}�fRBG�	�-b?XC�6�~���z�Z��$���p���I�O��w�/.~z�k6#��@=
q��%k�ujo��E&E.>���2����Ȧ2w��=3qIb?}5$�╊����<ݾ��׭=�2���A)�n�CX���ʦG%���J�\ǟr�T��8�+���O���&چ߻W��ʣPd�ћ�ҞDP��z��⋵S�dP�R3��Z6���σ��ܼ�[�Ql����*��׌� �_^�쐾�nˆ�i��s��FуX�#L�u�����#B����n�4� �C�*�����u/ߓ�MHQ:�"�%ST�����Cn���
H�Vv���!�����viq9*QM]����{e��g��u�O\�a*"x�@�m@����(��O�y)j��ϛ��9���������X�E��h�Du��gY���;|%�����2���� ��0/���_O�Ӏ�Y�]<��=$u��ҦB��cvg��a��]u�NS�z�|����4�4��&��Q�̜%� ��MZJC��0�!���$��k1���0װt6��)�ݽg�Gժ>%)����y�֪��EE�`�M�y�t�4�m�y"T���#��'����BE���X��9��O'�h�%���a�x��ߞ:d�@���D�����8&���{�ѶA5�N
v�w�;7~j�fթ Pk7�L!+m�#v�I�q*	�ҴO	��o�C�uKjFu���� P�^�qʷ/�����t����3�p|�2�}��R澸�)2�|�����D]���k�x�LN@𨸸8���U�wZ�F�})K�w�S�������-�mr����*G Q�3!��k?���-����'�K�������i�`b� ����B}��y��5
��B͝砆ⵐ*Z�g�޸����%ƀN9&����_��<X7�9r��h�p�/5�F<-n]Z�;`樠�����g{p[{��g{qF|ж�꿰`%Q��Urr+S{Օ�b�D�$�m��b_��x�lJ�p� -�g|s��6 K�������d@;�Z���m�.��FI�n[�vMO�@�7(�0�퐔�S_�5�/���ڶ��^
ǘ���S�>*H���czG��VgW���
�_�*1��ɕ6�����k�~���nJ��M���A�z��F�_�������6���;a��h���M<;'��8�-��*Hp�3R�������L�\�?���0)�F�h-�~�l��"���Qi�N�8pS���62�;۰�&f��f�:_�$�G�����^YZL]���ݧ����t"h����Phm1��5��q�Bd5��h���^ wTZ����*���"���n��g�e��ʡ�	j�bbJS���\>_/��ڹ�۪fJŰ�a�Z�ǇF���%�������:��~q�X���L1�W�u���z�j�-��yǹ�>k����y�B҇sSk�d�o'��Z�,߶�������!�(�-�bdu�@��8���.�m<���D��t�M��ϴ4�J��Y�?g��{Z���8^�Z��ŀ'�y� ���$����z�?oi��̳�}�	:m��/o�e�gN�܃�t\K@\�/5���z`� ���{�[��I7S���͍�7�z��i���,z��\��gh��+�`m�u|М|e�l"�A��S���LK^_�Ϩ���U���\�m�f��a��]�_.qk�]	WK�7�=ó���Эa��UuFk�e4�e^u���1�ה�C	�0�kq��(I�5ЩJ5*�,��5E�$@Y��c)r�vWW��F^���fA������l�~0-P�@�w�=,"G/n���۱���U�ٚq�4
���]����ܐr�<����e)PP_����伱�@�FW��V�/Cű��7's�o�����I_Nb�Z�a�Ag�:oO�T^��Jd�Z��-��׮�o���x�	eu���O;\������а�;�e�F�}�ͤ�0�'�
c0{Ԉu��^�����9�����'����ah�'���V�sr�%6m*\c��e��P���E�C ���H\ y1�</�>>���nwɌ�#8镙���X��ݴ�~�����B��2���A�f%#���\X7�z��Û�]���;.{U���Ӈ���t��E1���;�ce����Y*���&���UH r�RX�[��U�3�q:W�sq�π5���a�V--����l��(�\Z���:v��m�T�#�Ϧ�h���6F����������l��B?�ك�H+u煸����ΪTx{���*�=�O9.wQK�^~ ��q�E�K�d��-s��6޶G�0GU���y{�o���]�_��O_9����G�=�L�^�j����'e~��>�V�'�9�~�}�.��N��UӥE[z��?*�h8��f���������F�9ȟyoZ����c�ѳ�Ř٣/K475�1z�+�"��D��-m���F��#t��vuAH���{���� N�� �����'�n�1w�9�P¯���8�Q��[��?�W��*�_�����S�au�|˛��6���*U�e{���[��'��7����˨���|%�T��5b>�z�T/�JdL�I2[¬*�m��1���QyȢ��cz������As��Ж�ۺ����מ:���aO�9���
1VBf?۾���{�\��|��xy��*q�\m�@q��ʕN��Pm�>7���~�F�[�T��z������'`;J+I%u���Ee]�d7�\�+��&4}U��}?�+"����15��w��m�Ъ��ԝ.7�{�ű>{s��� .�=�Q��h��́������BnN���܋�U����m����[-V��=Tg`p����^9����E�9{�&�bjC����l��҅��Z^�'���ڒR	��"�Fj��o������f�%?����#��Y\��{�Exw�2�ѵT8�E���SP�ٕ�PK��8`�WoZZ:!5+����x���S����	I�U��>~��C	t�N���X�8,��T]��@m��j{1�E�z0�gy�W�%5�{Da���
!sW�^8���׋�O�П�r1�}�c��"�������������O/�b��ۯ��_�������E���_�v��w���w������*z
uF�A� ���7�;���'����?|;��<�V����K7�PK   ��!Y�H<�'  �'  /   images/289c84f5-bee9-42dc-8a56-be82ea7098c8.png�'w؉PNG

   IHDR   d   3   ai�   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  'IDATx��|�Օ�_չ���'稙�4���d,@`ȋ�����bl��[���5޷~k{^v��6�&�,���P	��&��z:�P�ι5-$v���Ӕ�VOW�x�ν��+�-]���}	�å�*L&��/�Y�CQu��+(**D�9�p�
�/�^g�F]�X�^7��\�-1$�:#2"��r���ũ�?���M�^�D0f���A~A�z?bI��8�1���������������|���K`���&�T/
�����D0��ǋ,�k
��"5!��"77������4q����j�"��f�ȶ;�^B��1"�!7��g
#���\�Ԧ��I�+�Q3�;r�q��������R��cn�M��@�[�!3���vy�]�H8�_��5�+��q筋q��/�Q��w����x��N`	�������133��^
Р츶a�nh�x�&�_�%Ņ���n��R�{����rMⱗ�H$X?7~t>��9���9HE��Oڑ�����Ћ�D	������044����z264y��5ؼ�<vy �����E0��x��a��������.Bw� ��,!��p��V\3�mm�~o!�Q|��e����_E@��ҲA|����և�m3 ����cA}5^~����`���wW"�L��\�N�ݠ�ݩ��أ��������$I�bg%��Dz�m܅67ؑU�9,�=���P^�b�OÜ{������>lh4���v�������,��A�[��1<�4T(Xд{=j�۰��^ܶ̌�yw"'�(t�6�Q��MZ�#��k�ȯS��t��T���>|jmrj?[��/�kf�4-���,m��So��#�H��:#	��I�9Ľ7��T�M���!�*5�Ev�]XR׃�m���V��l�21$����;s�2�+������:�K�@Sm��ҏU7K(����i~��XzO��n,�ڢ�!��+b4P�;�F$���*��fŶ��$�?Fsk�L�bHj�o:����h�v`ݚR��M���_bڗF�T��Klش7�����hlZYJ��{P����R��8?�ơm���t��K��᭽øv�'�}"�����*�zkr2Zs��8�7�������$�Y5h,����c��O��9�E���2��m�[0%t��S�8�=���?C�`��y(�t�]}X���Ic��E��q���
1DE��kV�a��q��G�ғ@na��lҨ6̯����c<Ů�$Q���X��;����F��j��˺d���>(�5x�h�0a��	��V�o�Jet����h���"(�(J
�vaӟ�c�D턂^��#ZR��Q�|�S���\;��+B:�F<�{�e�x�#Y]�|�4�#�'�R�N"�NS���<S$~G�.���PQY�g߱��SE=�5�X	���\���#/?���8�P ���T��ߩ M�fh~>�O�k�N�zS��(,,��
�z�CîD�*�_�q�;3E���D�q��4�Nbz��hP�W��4�d��'ڑ��ǳ{$Aϡ�����d1YT8�V����^"��$ɤ%	��-D�l���Q�u�e�D\V/+0�W[7�v��JJKs�^:m�B1��iD3�t0�0R�d*I�VEm�����n4%\L��)�1[�B����w�b��v<^/ȩ��~� ��j��0�%de١��$������m�98�\b�012���C�>F�!��֊90T����|���c��P>��~[Ř�f�mEg������!a�Ѹs��!|�v�:�`$NG�J�D|�����F�-��x=�ɶe���h4�i���R�:i�Gm�&BaQ�xɈDR�*�R�J̔Ĥx��	BK6�i�Äf�1��o��<���k�E���W�LAA
��Yj��G��PI�B�� U.��T�5����2�*��ܢTNՄ�.��B}:I�	Y�$ 	ڔ�T�P�L��㎯XCΟkEaI�IB��b'�:>Aİ@ ��J�見�, �2�PQ�E�7%,#W�O�\C^س$x' �	���3��H�YU���NP��C���Aj+�
"��Z���"������'�p}zz��%����R��x4I�:ю��2fn(�c�2:;;�x��##$d�}vww_���Hv��N�%$�
��X������1Ο?�ƙ�������yd��WI���b�=��J�����8>�ƈ���@5�:�?��gn0�սql��-�)d�	e�8ӕ�M��xuO��`¡�IT�¹���p����ّsIB_��w+ذo<&�"�����n���hkkGMM5IjL�l6a|l�fXbw��)ꭿn��[��Q�$SS�X�h�(��Ӄ&�{���H&j���mQ7��z���K�%��iLze��i8sq��_�Gׯ���2S�s��i�zg^{�M��o].3X��º��e�w��m�+ԁ��x��y���c�����Ļ���b2�B�԰ъ�����!a�Or٪yV�)7R�*��Nm7a��)�.@̔�+��A,u\�ޏ.w�����b��$�F���
�V�x�lLNN
)/-+~��r]�?+))���̙3�a�X�v�:ҦJɯmݲv�����L2����K�Cc�ϱ`�����<�{?U�߾�M"B��H���q��a|�{ߣ�0O>�$j���ފ/�f��f�ꖔ�����;8�Gf%\�.�@�O�MAT�)��t����,.ǯ_W���C?��*������ǫ��+
=+D�L��(;Q��_$����c/$
�`t�N�q�����C
3�&r�Ѥ�+�(͓q�3M�$in"��B+'2��fX�T�!�S����#���O#�薳-�ıfTSY;X3��O��Ts��/֎,3�k�ݾ�pG��� �FmA�ޚ7	����Ghnn�~����?�>~�B�G�]�a[|�7�����������|g�x�3�}�4����[=h�ԋ��Z{�,��7��5���P�GZ�NaIS�T�X�a�ڹ� �&2S�]��l��=tH����<����=y�1�'P�^o ���={�scppH����>1��z����\I72�ʒ���c���<g'����3	�����r!�Z�۷Oԫ���?�Go�r�ҕ9�jQ�bЈz�z�7��g��~�Y�[�/]`�`:;Hb�L�L&.Gh�����iA�X,.|EGG*+*ķ-ۆ�N#����9r���_���ĄE�2&=2V5YIs	lXex�i�/B�{_Cد~|mr�2Z�b�niFǂx�12{2z*�m_�&h�裏b�5K)|p��{� �u@���cW
{����ɕq��!	}#�4�*KPy�ʕ���H�MLkk+�4�<��9d��)Dp��f���5F��DH/�|��7#JS�D�d6�i6u�� ��,01	i���V2�m�Ol@ �6I~H �tZ'�۷4�_����W��4;F�q=}����+�C.�h��W���ݷ����sz�<����>
��8���'��&'� ��7����0I.���ygD��fs�ٰ�>nO���͖�Oߘ�
I>�/?�_�� I�L1���5��♎^N���`�N�h���,��`�;��c���E�%a
�*C�����M���eyC)-�"�8��րz��;�%p��y�gF(��OMM�s���EF���3m�4�\��K�T}���0A��!�ڋ��nF��h\B,��dԣ����b�(�C -�.J����v�CZ
��T#���l�2��.1�_W�!���p�`!�sq1��T"&a
��(��G�d/�$� �IQe1��^Mrr����h���Kv���!�h�(��K�(v1�L簖��9�9o	E�X+M�!��Ѹh�H厽F1 �L�Č*|]�h�3\Dy�a����*k��Z������ȟ����|8t��XX��Rr9+�yv�?�9ോt"M��@X��R��1_#I"�?�B�����{#I�a3bb:��2:�f��c��!���{ȅ`b�m�pd��/ፀ���1
�5�Kwm���e ��E��y+�-GR$�_e��UfH8w~��ݼk�|��.���4�.8�L�,��d��]�,B^!���	�v	"�z�J�'�q>J�*��^5M7 $��p���(|
��$[9&��u�Ւ#��/E>�6�D�Dy
Yv�Z���J�%V�b��Y�I�0)�v&)`L� ���Ե<R\�IS�0�6o��
k�8��L��@0&�2��d�/��"��-&M)���:��R	=�M:�l~��^c~G�!���O
b		�6Bm��!�xU�vZU�
���0Bg���Dff�LzZS]���#�q��?�T�a��q���W�!��)��hX��aN."����d�u���"C��-�K�!��T~6O!��rl$�DdFf�^�ǎ��mG�H��	��T6�IF{{�h''[��>gΏF�_b��߸5n&�� L�!/a�hZ�n2�V���*��bl��Z����z�Zh1iS���0�i��i�3��V�<��0�1Kuy6J
���Pt6t�H;�d��o=N�R1�2�E������I�~�̅U��뗣�Ӏ���x��b�,6tpvy�MAh@qg����NKĄ�m r1�1�pj
��$"e��Ń.�rҢT>�K�FN߳��ȯTV�!7bxx���!Z�Y/��D�\��A&�,�%|��g.�j&H(���R�T���p& �H"�Ȥx&=��wJx0l"���m�M$������,.k�10�`���db�; cb<��R�+e��R0:��#&�9�X��n���Yȝ��ՠ-��`�z뭘"l60��a{�b<#���0#d-��eM(���o*I�/�bx�S� ~��"�Fh6U�Ó��ǩY8t����J�����1"��PQ�#ߥ���bZq��j˥з� E�u��^M�t�ʅ1s?W�!ySbm���o�����8pD�{�����΋d���]3l�t�Ԣ�;�ʥ�q�zTfw��!��em*�g��ǉm�P���/�}]��H�����a�r{	Mu�l�*���Br���L����X8�x9��,-3�z̕�p��m�w�Ó*
�� f�r!c�>��M35��`H�L�/�,����,3��O@0����kVbj�=�]Q�����9}a܏�4��(�j�/�-N�_���6c�'��dBh+.�W70��#b�n�"u���n���1���Z��-~keD�^�iE~��G�$��&� ��4E����2�Tި��$��Q�d?�6f����I�K��,�KW1��i���c�P�������^��9�؉�� �֓IR)XIh�Ȧ�S�}�����B�N������d��4�n�Fqq1V�X�����MO��|B��	�ω���?�O±s!$�s��Q�PpM�G�]�Ԯ~��F�;D.�h���X����q!�P��*
�c���]���d���rƗ}�<~�u	�%B]�%�>9%����
�9����ɐI "\�K�2�'�.&���h&U��dI�V ��\a��	�����إ+�&WĹ*� ח�����@Z���		�Z��"�{�`G�J�i]�	No�+���c.C��� *st"��ۅ�-*<A�#�N*^��~��;)�PPS�mo�����3��D�,�@q�LfS>���^E���{��f�Q^����G�I����i��'vճ�����-.s�ԙ ׭)���v�X�4�����E��8Oyz�n��&Umo f�U�~1}s�}�e��r�����|��
���p�5�3���"�]L�{ǎ���5|H0M�t��L��g{�s��L�$����}�$w���e���bkl�F��]��r�'��"@u:�qg,��12��ט�V��waNyy0-��j_:p��Z0�тCy�!��9[p�|Z�R8zg�$.�:�F����g�!F��x	��% fāf^�O#?Ϲ�k�܈����!^�#�[j�z���d6� �a����TG�%|�/#���]�B�m�p�[vk!��T�ܢZ��<@�%l{���5�o\�s�SD�>�X`��gT�*��O�Zp�99��0N�p��i	��@=]籤NK�KK"h��w�q��̼+���H�g�,�s�Cx�o��{��`���I��O��
��"�9$u�0�'�-(ȵBg��e�8"�aDA����D��#?���3�$F�h�W<M1G��l�d�O���pf�/2�U��"F8J���01˾��"F��h�ef��{2)�~�z���ZD ]8�����W�y��\\�ׯ-Ś���h��׉�FFx��^�>E�����~�$���C݌����
Y���x� Ҫ��b4%�V�����*3n\mG�q'��^vtv�?;�g�
aG�*|Q�bf���y��_��� ī{�^�lY�Ӌ&2>�;?%����BE���2��؇��XVz}��H�����G�u����0k
+JO��^�$��M{';Ӣ��gڅ���P��ƀK'��r:�iS�5ق�G0%��K���1�1��5�B��fv���9�4�O�^hŖ�b*�<�hO_/:
ƀ��n�l�w8��՟&�4�=��?��bǻ�����L��}��@�9%�;���8�����x������Wط�Y$O�t�.ޑF{���'����c�Kjȇ�V�^�իW#??Oj���|������"�j>~�
�#�����C���{�	C/i��Ҳ��Cψ$�9�S���A-�sdi�u��Nk��0��4e|�u�uxі30eQ���r� �l~�z��}~4�����m����$�]���?�\I�k�A��0O���؈u�։m��6m���ƍ��؄?<�[t�]a`�[4�?�Mm��E{{Y�f���g�욅�Yջ�g�=V�g"]�Q�� ̐�����M�M��;^�m('Ʀe�J����Ua�z���O6#q�eD�:$G̈8���"�[����Y�CKJC_h}��pt	��]dg�cߴ�Vƿ>`F_4$���?���z�gp��O��&��i�|�p����?;/�u���g%�e�bzV�tb����g�XJ�|gɎFSȦg�`\���f70���iq�,@��&���S�IE�58دE�a��<֌�\6IT��XӤ�SX����������ޡX�3�S9��N
 �����_A�?C����e�#�}�s�������p�Gf��.�7�\�(�--�G��Ν�_�{?Ο�8���+ ��!,��]�51���2��&|�}�O<ׁ{�����GH��E�xis�x���8�(Ǿ�.R[3�K��up_�|�}�������܊\�	'κ�ٍ%x��v|���xys?V-�%s�FG���^�/w#�|%>�|�F�I��-��cZj��($>G�_Uu�'�.h��7$�����$p��s�����ݷ����X�S~���!L��k
hn� !��B�bf�B֋;(j<�����?,���F�x���¶�-���!���g����o�� �*�I�&N ������NP�fFQdM N��8Rnrt��#�$E��\~X�HϜ�)XD%��UM!5=M�'Nm��b+L17���.1冉ڌD�H&&>4��0��O�#/����'�Xk�re�j�̘N�bz�"����!v+���K���	$�Vd�ؑI��Lx�o^�d�fW���+�����0\��馛p��1�I���|Vd�g��;��!i\�%6�y�尀�񤄗v��΍7��I"f��Ji����E(0z�@Ll��A��X\��[�����ƅ$e�Z��qgL{v(&��m���
}��(R�����?�9{H�NiW/e��X�U5�ɦR�Z/�T/����e-�����Y[��K����.>f���f:���_��m���6�Ⳏ��J~�} �.<�"/,*��%���ZM�PRRL�������e�,��=42�`EUe	IuD�~qx���M03Y���دd#��;���Lrv=�� B��B�2`|����E�Q�Sږ�D".���8M����������"����5�k��#����(��e����(��)�̈́�y�%�N	=66*�Ysf9��*|&���˶���ӹ���b�7��6�os�1^���sZ��5��TVZ%��1e^�����	��qcaN��PaA���b�����O����9�x".���o����M���rm�Է�M�	��ʳ;[x,ٟ�ZL��:88���yb"�i��d6-��L>��&UA��eA�S�|n�	�9��eXf-+�f�)2�8U�� ���L"��Bp7�^�u����h��=����{\��1�W�&�,�	Go0!�� //�����_  ��_�c-��-�Xm%-���'�"-���B�k�5 K
{���NҚ���Ƅ�f�q����:��(�����ܪ�yP�I�F���>��<��3�u�&'�`q<����kD�������C}b�9ydBS�M@�S����Ǭ'䗄klD�e��,�TJA/IiY�(���^���`�;g7�e���O��F>�]RZ�i�W��
�1q;|0�������p�bR�C)����{p�2r�mI���/z,�@E��M�u(X�Fu7/��ۗƾd.��"�{�~	!�3I�H�$���=��Q�l%՛�ǗOc|:����W�Ҭ|�I	:���>i��˹���P�r-L긨7�J�H����2���x�x
����'ś�8��|Ԍ��+`Ӎ���Q��b@'��z��N��cid/^F�"�G��~�9�嫐k�K�8��G�*�g���W�;�zLE����2�p}Ө��n;aCY�J��q�r�����!ݗ�VA�Ɋ��6l��;�m@'�w��,�]��a����ψ|ϝ~
��eu=��xiP��n�'(��m~Gں���S��5�}_���QW���9���~O�1�o�eĵ�>���(�9�'::���6�rك��;����X2O������Rt�=�������Y������A�EO�����5(i�!�G�͟�ĺ&�l�
i`6A�'���Q��W����b�������0����[���ϑ����c'o��u7�j�6�Ͽ��{^���7c�(���Zs�$�?�w�<����t�C$�A4�}����/���	��G�&������&��Ʉ/�����$�x6q6����n�+4)����4�:�Βc�`iL���r�֞��B�ۃ�HU�T~�%��L��Թ��(��Nc{�?a@C}%�n��m��R���Yh�$s�'�����)9���f��i3�W�^
 �o��eI�<�����6F�8�&�T�pʃ������߆������!ޗe���Jh��
�k$�q2�5���>(��;dGmm>��),z�mp�	4w���o�} E���D�4�g�p��X���h�vS��R�5E�_{_C����Kho�3�9��a�<�*�Q� �"��N�U�z΅p���}��/��7����#��;VIp9@���T)�r���W���s��.���̮%I��+\��^�"�΂Δ)�����CX�����&��I��R�T��7���0C�6�63�O�ۜ8����!�d���>���(�z��^����a
12��.��`�{�=;I��z�I]9~����BJ9��e��O"�,�z�q�W�`96E4��23��_���Q.�2yA��F�sHIe��jQ�2�r�    IEND�B`�PK   ��!Y����7  �  /   images/2b66d102-ef9e-4dde-8ee7-817842500f7b.png�XwPS��� R���PBU�!��B	M@E)R tH�J�^�JGH�.ҋ�PD�@QJ	
�}��͛�����:{�{�:���={�8c]����dddtp=��YD��
p6z�d�>��zh226�s���v�^"������dTg	�E2�3v����3 �)������7?�s��ܒ�G��/�?�مg��EAFv�o�{�/�}yU��..��=��} �����ɋ	�F��>/��-+�>�1�Z�%��|�����p%��9�#|*xPݎC��S<�'���o�9�^>�W1L�Q3����.�Q��Օ_||�*~d �֋��'uy��j.��9Z�*� �u��+�>E�� �U�L�.5!>�n���f��f�q�7Q�>��-g�_�T,�X_k����>�:�c;����F+��g?���r�q�1�����Uʰ���r�S[0'H0]l��?�הۖrm��O�������98��W�8
�}�)��;C��r��3���&��?�.���d��ƛ�d��M��X�2U:B�72���/l�b��!�#8����G��d�{��x���m������#럀�(����ū�e��}��� }�g�
�B�!��R�����R��QD��z�_/�)��1@�2���X�L�d �IQ�l���Fb� ��yg�W�o��t�Cy =�(/O2I)IGP�yYr����?"yd�{n�y�kΊI���;���!����jx{����QB�
�����8/�<$���9_�B{���H��w���;�a���S����!EK��ű���"���l�4kf�Z����Y�5h[Y���z�_Q59:�eɔ��5
�Iu��qV}��Ԕ��� ����TH��.���F���b�	�mM@&�cA��	�)�����mگ��wD��M]�_����Z�)"�P��R3���Õ�m��~�y� ���,[=lo��� ��8,�Lć5��63�*(L|�H�	�A8h-����"Ҍ*{D��e`ß�Cy ��g\.�PK���$CX���U����a0|�.Ȣo����G��EE���Ϟ1�$��|�B�ܵ[֘hkת���(k
E=��/��-,�$bb�MLc�虅�/�6R=xW��4����ZЋ'R�Uf�8n$Ⲷ���5]P�I1ِݰ�C�d��{I��M�7��B�!�P%�A�ml�A��ƀ��$�R�zi�pT$5h��h�p�V+d��<�~`pn�Ȋ����	@7=*谭��x8-	�v�'4k�߲t�]�Eo��ʍ���\~5c�U��-�Y�Ԅ ���D���҇ӌT�L�%�I<�X�(�,v����Wn��L4����P69����'8�r�rI(�d���`�G0�G�14�k�:���
��$(�;���lEo�y�B��^z. Ul����i��n?	���L�{���S�1'�:����\ϴj����^P".�� �]�@�d����|�� [l�T;���|^^�+}T�{Y=мJ��x��]V=�IS��7D������o{_le�@x�0<<�e�R
@��Ʀ��I�Z��W4'Vc{Jq�Ukg��ʀ=?%e0W�-�TT=�	�!�fy{o�-+#*�S�OH�)� k�F�,ѽ3�L}k���n���G_�,}^]�Ԉ{|������yο-*7����U�j~�afh\��^"��h�!�`؟�l��?�g�MMc�|�S���X{7�E��!�����r�~��ۜa_�}�p��&��D��%q:��~Wh���05����v�7��Qskk�
Qf㦡!�og�%�Β��V��t� ^�kp���v73�E$��F-v^�.�*r��NbX�z���>r��y�5���+�9���9�֫Ƣ�z�x��]�@��E�]���z=�N����%~�.��"h)+�ѿ���k�7�W�u�����e�⹠�1�}�?��V�v�@g�Y�a������%���כZ���a{?pt�n�3�j2\>�e(oí��8�*��e��CU�sf&�����3�R�o�^=���ǡ�^1Q:V�n�z'B]�4"Z�\5�zH\ݭ�1�q\7�2�H�}������������O������a�	k��\�1������ȷ'<��S��VئҵJ���`��lu�f���tAK�a*d�$����f����V�8�zK֓�z�V_C��kj�g�^�l�A0e7��F�e(�͝�ga�5��i��ʘWk��zT0�MH�	p�۴�f�Fƭ�EFF�W�4�z7�P2[��`st�c��:S�@C$R|z��X��#OG^%�/)�vr��i�	>�v0ʓ}��S�U�+�Nf��V?���[�M�RG�;�]��m�mG������2��;��pk-ǳM>`���`'��X��wTtB���X�g�/�+�4��Ȓҋg�c�Yh���.��7Q�0?���U�S�zw9W��C%�6�u�mƵb�0�+Y����������
H�h2����*u���Y�>(iS�(�ɷ����4B��u�Z+��0�����t)� � ]�I�	KoL
�l�y����)���L�whm��<��-��>��=z�$��"[#b'��9!��r�������OO�h��u��vuᑑ~_��i�����D�~CNS�z�흟J؍�Pfa�~�ϊ�xUk�2�K�� K�U5�B5t�F��z�ќ�l�zO���w.�{�oj��1�xlb>3��b��F�4˸�i�D���k7��UT�X6=Dv�O�Z�2��LJ�94, n��P���L �}���mu�����d�o�K ��p�s+�`�z�gup��,ڒ�J����o�)��6��u��dw6��m
�gf?���o���<M7(p,�b7�碨��_��נ��{�)�d��2y��z�ɛ�-�2�1�g�72�"�r����k/��g���hA6�.*����T��IA{�P�4|>i���7=�%^��0d����J՞+����y�:j�I�h8w�OT�n���^�^N�s|\CZ�劻�Kp�zY�3Q�):��źC݁
��ƌ 42ji�*�}S�!�"����0V-ӧ;��e���:k����U�d�w��[\ȯ��dzzz�>���e������ Ґ#	�Z��N>�����R:C������@����ki�����e���j��1�F��\���?�J�<Q{�rO�����B�1^'m�����A�d�X)9qc��ai�w�j�gN�隄�>s
�\����24������5:��(Ǌ���d-�ޓ�=���rT�,@,d��FU��E!:S~���5|c^�-;-���:���X�)�4�M���*�0J4��n��Pa��o���\��g��ե+�z�[�)�o����Aw�f�KpK3���蘏�<���Fi���O����3�ҝp����,`-V��͊�5���EQ�n���y�!Rey)�ҵ���վ��9��j��*��v���j�Ǒ�����`���=�&��h����8��-b6m<�I��nq��9��Zb��B%��[��n^��l�%�W�۶��O�����)���pa����M\̞A_ix�쑋 џ���^�!��&''g!��x���">�V/���1�__��-H>���`l�;!}0\��Ee}ˋ�n�y��:f˻�j�)��� x5�K����u�pu�F*;p����%�@p���Hj�W�Q\����W=��������X�����Uݒ���J����G��ٮ��J��� ���DB�ʾ�����4ܡ/���%$s��5�N�fj�m��$�_RYu-�*3�gdd�J��l܋�fz��ʪ[��'d�U5;��td�_��?��ų��i4���� /5~��&b�.e�"r��R�2�Ƅ�A��FE]��%2δ����7+�,)�<��N���։]�ϯ3"�u�R��y�<����h���g��A�hr�ʡ�A�W9(�&D&��7���L�Z��$Ξ�o%C)�`0Sg��L��m�g��u�`W�ISc��W�|Lc4?!�4�ֶ�R��$U-=�N����g�r]�B��pq�ʒ�32d((0��B �{�,l%N���F��s�Cw����_G��^ʰW���ǜ������tsSl��͖�ҹ�q��W_=�[�	F<���N�5�Fc#�A:�J��ҩ�%HP_O_����X�����Ș�[&����y�n�-A��C����6���w�(y����N�a[�<i6��w(��q���Ige� l�4n���I���V�Phfӎ��8�tw*)�����Mӯ]y��Ap���*���#�������4��bq���snE��u	\�V�i�/PK   ��!Yh`Pҷ!  �!  /   images/4b60cb4e-ac73-4aba-afdc-1cf5937e57a1.png�!MމPNG

   IHDR   d   o   %e�   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  !?IDATx��}	��u�WK���hF�h4Z@�b��-˖B�b�����!���'�|b�CVs�3�q�#�lr�y/��`�1D�%����/�e$�F��=�VU�������Qk�A�{��U�]]]}����:.�<��c���7��;�a,�4�֭å��>M����O�Υ��KHQ�O���3)2�d��<���*g��{��y�>��2� 1-�C,χI�!z�����P	"�?RTbA��C��Œ��_�I��T�j<��0z�J�W72� ��O�Ua=QQ4?,����,�2>m!6��+����I�Z�U�����˲�	����?H��������'��@�jڿ9>�Ĵ��ʊQ*KFS��ea,�z������S<��2@!:�
j�Ytʍ�sc�O6wT�8҈�=�����{��8��w�}�V�2b�ب�L�"룐�,T�D0sb��zz�a(��.�sF���0�O(�	����a*k�p˵;K��_�#m�p����%�>Ҍ����6l؀]�v�RK.@�	���^ȅ�{�8_g֬Y�����&�Ju,�����'�Pۉp Ο�Ce^�Ч�9O�8?����ޡ�q��Ӓ�Qۅu��8':k��D=v7kN!P�J%C�6mb�e/HL*���7sRKe3��Y'��(�?�>�����T,���� �($S��,G���0�
Ź�|O�f d	'�?�"��_Ob�V*g0�&��Ϝ�_���p���~\<a��P��J���\��s���`�ԩ�6m��p���25�J������J�ta��J2��aZi�[� �<����{��r���`���l�[6`F��d_��-i
��G��3O�dP�rr�0u�g�����#�����CKKr�V������{0g��~��={6�� 
_��לƲ�0�B�Gɘ� +c#�nҫ)�Qt
�BTL�Bl��^�}w���ߢ�M
��(����AX����F��Ə���?�#Y�h���_<����
��u�~l!NuO��-r�*ʭepp[�n��/��H$�Wǎ�թ�\�w�u�~?���Ĩs;�r|E����� ���̙x�n������R�H��5�� z��T*����X���<��f����z��o�rV�L7ӛpk`�4f2��P+�4���F�{t��%е�[���R�r�-hjj�������9��c�p�B�}��B��d2�3UU��x
�3EX���gnGyh�H�@��l�@״��9L��_5|5���~J7��`
,�m*�<F��p R���6Q�lW���?��0�e����V� �\C�]�C����e��?0Ps����lm^�#�3�A�Ȍ��c}���=�Hs����җ��G}###�����g?�Ypu��X�-���"�=p� ��������9S���g�٧$P)�l��L`%h�P��f	��T� +.ML�moJ�+���
������
v��?1o
���*�����9���>2sC��� Fq(��"��`km���N|��8�<��OÄ́	¼744�֫7�,��������/�; s��E}}}�E�)�[o�%.굉�����+pݜb�b�޴�����B�@+[Fe1_�� H�l`V �L@<L��Ҧ*�Ӡc`J`$8��a�#̚9���yG�4b�e��B?kH������5}��ս8֚ru4�|�0Ϙ1#�����+��k�axx�� a����ǜ �������wމISf ��:�rS'����]aY�c�����V~��	f�6	�������	n��l�ထ�6n����[���SP�����ί�gYqGl��aa�Pp��Z���F���}������w�^9r_���l�2����"R=x��R^^�q��Lm޼Y����_��{()�ƒ�q��(���Ri��[�Į�EЫ>*�QP�M�'�$s bf1$�\yؑa�4 �!�4;0��B������S�V}3���`��F��(���n��=�u���������ß����o|����׾�5a���M?��$/ �E�>�o/����֮�]�E�<�:��ZrH�"����K(X�M�^�Zx��"&��4� �ad\�F�������L���$`�ۄ�?���V�y(%Ka���n�s��(ߒ�?�'�o6��܇��	qW�x��c�쫈$T޷��$P ^vp4�g����R��@	V\}�S�b�*�L  iE�G�j>N/)�����61�$lP���<�ʹ�N.S�M�O��bbQd���(A�p�!��撏�
�ޗ�;|-Ä�(�������W��+�濵�[innơC��`��Q��9�-M��ٳ�[c�e`�h�Y��#���]�l�"�$����$lF\�ZV��0�I�[�,v�6�
�P�;�c:b˄����F�X��Ӡ(�������Cs���>i�l�H!
�� 1===b��;j����H&R�1%6 �(���u��SE�D�C¦��5b���������c
�i�d���d�b�1%%�c>	$��F��$��$"1�|O.P�ML�H�Ϡ��M�)V�p$��][����,�%S�� B$x%t����M��`�hE�#��φs3�x��J� �k�!��}���|Zd�x@������yhi��h[4��%�1�����,A�����gP��Pb�x���iX�������b��lSŬP<@(�o��EJD�
�D���1%��S�����gkºoi�J���p�����?+�Ԫ��do�j`2�q39o�3�n��	0"H��'0�b��
��*%�!v��43k�d����
=��!|�/k���I���)g�km���S+ېH���H�+�uSX�x=���]��~�6+>LbH��a�l�v ղ�!@�����]"[[�O�X���nJvc�!n���n�h�9�����F$�D�3o�2���5Č�t�F�]	���e�Xb�1�aa�C���5�UQ�rE��e����>E�f�T,�~m�q�昿�?�+���3�7ǦK�`�[�������D��:�W�a�>�`xDT~r������}'+2��$�͗Б�8f�Xn?Yq�{xu�d��|�no^\���rP�(0�T�kn������}<�z1m�a�
Q�#�|��TBWC����K���KM��**K���q���'y�-k�܉�o���p��ĵ�Y��"3������v�n�d�`f�0CVj��+�u��N�VةϝvS�eN'����ἀ�^t��V:�s��8\/E�z�"�u��%o�ʦ^�������N�ZD`��NW/Y������k��`�	�����B�Ǎ��D�j	92r≎+ ��d3���긏���t}F�3�J�M6]
���	��:����͹. �����q��3�����
	3�`�A���zi��Ӷ���f��n��t��k��wh��U��~��e~�Su���/�>��z��,���F�N�5ı�wlv�0m�A�T͓ܠ\c�e��X�M�e��d��U�j�Xr3R�fȶ�e	W�/�[V�j^͉ɫ5��}{9��d�SU�,�(��`G�+���Xr�{9���-���v�_���ӧA-�V�<
��U�����z�M�q�&h��K@�@\�QU�����f�.�h�꒶���Z���ŗ	
}��fd�H�-EqYb�Ĥke�b�zI *�@t�M�% �t���3E쨧��O�߸��pDTLF= 8-����Ǔ]���?�2�%�m��R٩��Ldd�b	��T �!.�&�c��R���2�"�F>q*%=� b���b_-����.��Xܜ�:zز����5�-�"���z�\١.�z����4ؙ��a��M%&� 9[ٿL	L�2����Y<u�<Ҁ��m�t��<S��qkq�� 1�WZ��zYU�\D����.D �N�oM�܍����x�E�= �C�a�j��U��r}e�Z z0d�zE0r����L�^4	�5t��N��v�39�K�+Ki[/MT�ws��N[@��"�[P�r_��$��}���i��fk)���e�V�[_�1[z�NG���%f&+�N�1RĒy���]+�֨���J0 %�d�ntLUڡ�b܅.ƃ|Н>,����O�أp�{�;����֍��hZ%��&i��+S�+-��CG�ME%�Q���ȮG
��W+ǧ�f��IT�R'��$�O��?�&Z�_�宴/J������so�@=a�"���r�-�=k&��&��*'��}-BQ�Q���Ng����������&����M�윬����E��o�q�x^�	�v뙛&f�ˎ�҉����~����f���^aw��s=�WH�0 ����'�R5���8/�e� �C�����J)�)v:;�Ap=��:˭PLGY<|@!("r�"L~*{���sv��ny*~���:fHE��t��\�Q���S�4�>�BQCp+u3���H
M�!��" �.�3/��$d�D�{Ve-��!>'ʂ7�R�""�N3F��(9:�Hl|��e�����${԰�!��NH4ݮ'Q�]uR������[r��-�)��[i �¢�����d�i��+�t13�i�]��t�1�("r1īC�)s�In�2C��T8��a��LCދ"J�p	Q w��O��MgLKw�v ��&\թw)�y�[5bOn�U(Fy ��(�4��$]m"���b�Ʌ���cTF��V6YG�]~�͸f*#����""�.9Ə���Ԡ=(˔I9�N����{C^˰���WVS����;m��G(��*�<-�(��p#�]H��kY�#(6Q��(�TQb6���D<Rw�.��I�~v�9v����kKrx�����h=d�\A�423u�"\�۬G{���fQ�Q>���~$X��I���p&P��C�g�H�F<ڮJ����)�#J�o�$���L����R�(p��r��m���z���l=�v�El�ퟏ�.���p��;G�=������&�趙�F��mU��tB|��r�����Va‡�`��<f���Y2����&�ɹ����u[�ܜq]�#�${��\4[��|�L����X�yݖX'M���V¡��Z���~����>�v�J@�R�hȜ�QN#hDx�~���S.K~�$��OF��H�{/���ȏ�!h����S��@1u�3�i�L>E�#�H�ά��WH���9Ч��~"�����T>��<�D2���S(��T4[c�b�"wRM����vtH��~%�[�D��Uo����idɒh�I�Lj��Y�ODt��6L�o��N�9��?��^"�_P�MeQ��s�a��J��-�$��&J2��j́�b
s�MXv��ZQ��8fKSya<A��{fvu}?�~��z2��"KF�*A@��"�%s���f�)�5���<�� ]���/�IC~�	8r/?p�&T����0���:݌��K�,���ò(a���-bG?��(��RAgOr��gZ_�;3��n��^��Yb��H!�����3Y�I��Єi�O���+�`w@��y�x;�c�Xa�a��x��*�����cO�
��k�+�\�����8���������I[��f�Gd�S4]҉3j�`���y�������|*v��w�m2���Q��#q��C�x�~$��^�aH�c��0��M��j�H�o����R�x#*Q	����"5���YVh ��ޖ��I5�o`d;x��p[3���&]٦K)I��WÌ� [��O�	��J���h뙆�-ܦ~l,�'�$��d-n$F�ⲥ8��4}Z�9�~Y�%#*^9N��U��H �M�^������X�-�`�ѥt|4�U���R3p(�i,,ya4K�ܤ��T�[q��[R��
�V�$��EU}v��qŶT&�=�]C5bպ|2�Dʼj���M����$����+>؇���jε�rƓ�����`�$�I��X�:3#���dO=���GN}l�>& <~��SvG�A��P�r��>U�%�+Ἣ�t�M��
��>Y���~���T6�ALۮ�e5���Φkؚ�'�k�_�<���#?�t�`T4.��Ay1�c3R��3|r)#�/$;4ME4����CCMC��8�5���-W�+)<�J/ΐ/z��L%G�[��~Bt?�d���2s���3z�0W�nf�^�gxVe~�B4���i��_���2�{
\�ȂO7��π�)��!s�l��|��\9{���\Bb��Ǔ^��$�1rL0#͊���|㇧�u`�lnb*�b�_Xi/��W? �ɟ��դ��Q0(��.��ߌ�Y��+����"�T� �G$�_�����(��?���;�8"�^YY!th@�� ���o�.���;@���w>��ddX�RN�|xb���Ce�����)}"�Z��[���&�wx8���t᾿8�^�u7�Ry^�����Ւ%K�q�F�`b���IL󋵫(ʊ�&$��S?��-z��7,�M�f�K�}�����ja�L]������y}�,��d���_��=�"�����;g�]�`^z��&M��իW�W^�q������}��u�ҋθb���81ԃ�is��.;��[3f�&ḫ��t ٿ��a�_��0T���|����GĢ`���Xw�5q�Z ,/ ���%�(⭷ފ'N��^Y�?h�����3R9�,�٤b����iW#PYw�q!�$�y^D�F<�����N^�������* ��9��}�D�y1I֙wAIg��|��Çg,L̨�z�>� �}�Ylݺ����� �������r��%A�}H-J&�B��6" ���+�2Qpɡ]0�����������$�������ʸ�������^��1W���O��{7y�Ռ�=*V�v��M|��p�u�aӦMhiiAdd/�
莖��?Q1���^w�(v�o����]�U�k@�j�����'pD�y�~.�Tt�����<Y�%��)Y  m�|>�����/�CQ�����X�{�ʕ�o�C���F��;Ώ!L��_��W3Pv|�ҥK�x�bqq^�o2*Ƕ����4DWռky:�p]-@�r"�Փ)T���[�d���ȳ��e�Ć�#�G>"*�Γ��c:����/$���6a۱e���V���P>/�̫l3�׽e0����j�cɘa/3䩧��}��'~��qH������`O!��{ёX����Q�wg�O�0f".�_"�'�B�W�fb_I%��W�z/���Y!�=��L%a�/c�`$"��\����(5}����#����q��A,�U]�s����\/+��'0:::��}c���y�Ν;��ى;�MMM�B-?�c-�;���|3�o��!���9⌋���c=g�m��<��C���'��|A
�|�39�����Sܒ���c%MzxLڗ�!X�Ӯ�L���y�'	+������m��^�X2�P�����Rb�Z�[�l)��}6)(1lmm����E�6}�t��B���3-�j=n����(1*�/Dέ+u8A!�@�<V�0/jƹp&���y.�������=���b���DL����_W�� 4u�Ykl�'08R娴 ��ɁJΡ�l�����K���~�m��~1,	���V��LG����(�9�`��1�uK���aC'��v�?��%�F��܀�X�{��W�O��8|�E�r�N�X���r��*V5�����(����2��xy�D>��+<H�?HS6@�b������F0o)��Zk��7��zWW�w���W��e�������U�V����?Et}(�3^���{�?�)�f4��Ť�h��
��O?�@� �����&F[�Dno�ɞ��QZ�`�J��)J���Əo�����RJ����.��vG�|��$�!Z��CK�)�{�^�Ϗ�	�%�?BZhT���|¡��vv h�"F�<3cjK�T_[�%+c�&tM΄�\r�!z��֭[�K)��B���5E���Du$�
<���ϕ��<)���2R�5���m��Z*���s1ip�0m�項�>zwG(�����F�wM���_�� ( ^QCyz�_�:܏�s�GI���˿s�E!/O�9�J}VGʭ�RAʦ$E�c ��2B���P�$ :)�kD8L�%��;фCgk��hau�@Xt5�H�~�}oL��5R��Q�N9D�����O�	$Y�t��	E�`��E�o��R�]�<���p�]� ^�Z�V�yoϓsb���gw��=vƫ�[@
���6�y��C��&E@ƙ�0Ǽ���b�    IEND�B`�PK   ��!Yv��� f~ /   images/4d249bba-3190-4770-b321-fb8fc027a237.pngl�	XS��=��-��P��(We�@�U���2)a�)2�\�N�'"��@9P0̓��0V� �� B � ��oZ�����<}�޳�~ǵֻω׎�Yl�z��[1��9HH�TKHl	�,�䧙�g�|�+��f�O�f�����ly:TBB�9�練�'�*�9��F8�-A t��C=�{���f��A�ۡ����辱Â����{N���N������-Ү�7�g���װ��6���������7!AAQ�}�C�����w4����K_��������R�{�����j1���}{k�<��=1�VF^x�/8o��P�p�[L,��^Fi���0UX�����W�C�ʰ�e9�N��'�"�1����J3�����B���Y���@�ڌ6Fն|/e���YMFb���7Q��yp2&�(�0�6��j����Հ���_ڟF�Ǡ�����c�t��ZD<$����}��p=�bu�l1|�m�)L�N�Z�ش=�Qm_}* �5�)�6�dK�.�
�}s[\�g���L�
Gwj��Yb�>�T�n"X����m�Er�$	F6��fw�oV�`r�������AU��b9��X��E;Y�{��x�nް�m��C�qF��p�8ƽWW��^�tO{���1����?
�1�*b�~��wң�(VN�[���i{������ ��91��\�-~�sA8�O
���R�x��BL�ġGgº���j�� <��qx�V�{沴1��tfo��qҀ�aHW��@p��H��׳����*x�
&Έ��X2����]��;_�O6���P�Z��D_;j�g�9f�몫�fQ�̩��22s��ܾ`_�?���0H;�Y�\�ЮB� W�?G<�-
�ѫ�С'�$K�<�lɠ'�����D^��@�P>�p��9۸�妡��(�n�O^hb�^�a��:�*��GA�0~���A�̨��r/����
� ��T���R�>�z�
��2��7G�jL(�PL-y���J�#ݖ0|6\�ѝɒL
��/�=����FZT�GA�`���[�8-���P����B(���0��+:���%��<XǞ��F��ʤ֜�����t+�&<у�R��(l8r�9��~�[���@r��2�4Qs[������^J�+��s�
P�L�|�H�$t����Gl�5wZ���v�]7�௠�2����'��|n��K�NcB�������œ�=�O��7x��̹v	]�+��6�ryS���i(f�=a!Yx��b�;�퀖3Qk:�����m
c��AV��/gG�,��WQ�e��^
(��WupA,��}F�o��5�()�75�t��r�U�eo<I<�s7/��a؍;:�-�J��c&��>��:� �H�ys��q�5�oO��Q�E�1�h��h��~���p���/Lg48'�����yb��J���;�70�����Є�8�)��G"w�\���*��á�|<�1��Oq���5N�7��3N�	M�	�x��wJA�I�AS�_{�ǰX�4f"&-�nӒ��Wh7q�>�\,�z?�Ҍ���:�
���M({,\���-��\���ip������R+np�4ބ��������
��(�Tj	O�D��0���.FAÖ!X| ��(|�cA/x¸�bt(7��$v�'@���d� IܑUYZ�<E�F׬|�5~_�j��l�$��p��l L2�$��M���U�#܇�Z l;O�aV�\�e�p��8v�*.�-ʜO�%�t	��bA�3M��s7A=�	*e�&*�d��c��P�s�4��w � ZJ���2p�$v��ʵ/�'��QP�N���y�r�S�$��6�(�{��)�Ѣ|�1 ��"ju�౓؆�)��q��	��!�fd<>�B,�#5{�'��}S�;��d���B�x��~*���۲4�*��%�ݟ��0puEb-�����}����,!Ḡ���3jA�X@�{��9ǰkA��_u���C���Uv������8����^b��`���Z[{{NFN�����fR��M��A"
<p��O�̬Q���@7g�C����L*/���g�Ν;o���<�x���ӧޣ������fM�7�.w��$��x�p�G���e�\i�T��=��-��L����Km��*���'��m��t��Nc-�O���0V"���&����������Wd�nl����j/�~�����Y 02�s��]*����E?�'CY:ї�)�//'�������K*舃��mɮu3팆�t9��\R1Qy�nv󐁢�*p{�>���=J:��a�o�S�ʽ(���#0.� �-�����F��赶�֯i\L��h6���Nt*�*#3��H��ȵ���>F]PLla��a���㞞}u�#M��ȸ������ᄞ�R5^���[<���ZҴ�Uߕ{wt��dge��v;��� �ȋ�/5�LO���I���ynO@{?�.�,�A~6u0G|�a��P�=q��P9h
ix�~��|/uf�Jls����p�%���XGz�ٯ�8��Og��C�ePG�*ãQ/8��z���0�C��>��7��6Ӏ�97>��&���%�j(q�A`L��<	k��L1]`�����}=�R g}yᖸ��J�=��� i�A�탢��^#{ל�-h@��)7�2�K��W�^e�K�ڔC;�@Q��	ۤ��1����+�NJ�ݎ�yL\>Azس�Z5��k��@z�H� d�,.x=���Q^iS!�F���ȕ����4Ǌ��:xB8�Y��&�&��Zԍ�۲I-)櫋�����<6��
�6�i��W܍��yF��/�N�^TF������=�i��t��|`F�$˟Z�Sf@��t�XY>	*n(lچ�Z*,��C�k`�=�E"L��{6[����S��
B[�~e�*�w���`O�6=�8t�!Sq�����^}������fO��"�I���ΈuHޟͱ�Ep�mS:�#��d�F}|h
��V��o�/�SOF����8���$>���Q���l��N��3#f)'��rCe�9�Q-��s馧`���)&ô㜾�tHE37����wS[�&*�cJm�x�MY��}�cl��7�E�����b�A"]�.��^!��f��d�d�����Qը�2nz{e���-��w�`�s$z�%���E>�qP�w��y����d����`V^�Y�D���œ����˙i����| 7�yy�"h�H0��_
���숙����r�C. X�誀3��$�6Ͼ����R�i�ho�c��m��ZsKQj��I�4T\�$Pv�ހJ�C�r�jζ%��7p�C�<���.�㥧H���f ��AT"��`~�ސ�O�,��Pw����[��6��ͣ�
��(GnW9b�����T_���}�=�������b�� ���ct��2jؒ�����U�cDW�pC����$���c�A�[���ױh7���ⁿ���|k��4�&܄�@y�,��s�*w~�_(+�X�1x��$	~��=�u��aXL���F��;��j��&�I;�oj��ωf�D����\�3U#h��S�s7ܗ?���Eb���(5DaIf;��}opn<D~����D��F�`���s��s.�*M�ܺ�BG_�
aۺBx*nP��ǰ�4kv!z��u@,�(k� 9�/���)�#_�..m����2;w�;�L�uT�?�VL%�<O� �jv�"�J���r�kS��-��X,��a��s��%���s�Gnl�f�]�,�K	R���#� Y��bV#8������ќM�"�L�C)�YX��c��lT[�/(~0�L-�4�96�VP��-Ud�7Rf�9d`��߽@	��+z�_?:�;Mq�� f5DO��$�=b�v��ſ�P��KVA7F�����~��T���2N��~�0PE�F�O�췢6L����<�nw�Vr�S�&W�ϑ���^Pa�Ą�sR�������jf���j�<�p��(�'�4�Q��zZ�c�̿X��F��7[q�U�~@t����w����$r���=�S�=`�. �2���i;W�7N�wD]q�����Tz0
����O�0S6U�KQ��j�KjQ �LP�17�|p#��L�ɏ�@=�����?Pѹ^�� ��b�޻/8�0<uS:E�;Nw%�.�u ��椝�w��3���MI�X��h�L��t�)���i1s]m����F �C��oq�F�9�qh}J&�s`�-P�N��Yw��'��YOM��y�/F��� ?n�KŨ��=[����*-�?M3�+^Jb��$�i�����M��u;��~xJ�`'�o����������a�3���2��R?���������#6'1�"<|�:�%F�`���	�h	Z;VmxC���#rbR��O���4O�3@́֜f)�?O�vm%��Ew�#�����ϑlQ��9�J�&^n�_~����G��$�%���R�N=����H�6.M�Vt�������|������}�#�4%������XC���@���P�뢒�AMӏ�2��<݋sv�⡬�:�f���%߬�� ��*��b�r�N8���7/{��I�8W��r"�3�xܱ���ίw.wH�|��G�m:f�LH1���F�.��]�3�0:�!>ÏZ�ʽ��J*�~8�=�ο�rB�G�}�1��%��uci�v$z���|���ypq$q-t��V�O�րB�v�9���Y�:��>�VyJ�W173[�ĆG�g��YԺ��S�a�
=f�ik�M^��'�\f,�ԟd�Z��	5=ͱ/I���b��8�|:�.(���(��v�E����\��XҶ��ҝA���Q�d�j�D�:2�x�Ǉ/�ƻ���e@�L\�t'�=R��eN?��LX��͉l_f��_��]+δ\��W�Ye�Y�C�-(,4��7-�2u��5Fż��}�%w	e~���# Nt��6.�������NS��wM��:4=K�z�2C�5�Q�_�4��>hl��\\�M� |�2�����U���㙺 	��3�qC����j+Wz��W��F�B�@k�qCC��|��?zX��y�_<l��8X+X���u;���!	��|/�~�ƶmۈ��[C�����)[�ϊ�z���̹��8���KՊ�@5��Q[^8
�\baVH���XQ�a`X��PE�����t��ZrD߇W7̣�ˁ����&2� ��������sZ��.���v����TaHQӈ���,��$�J �zМ�P �ߢ�[�}o�io߾dh������y�����ϰk����N=��a�29J���*�ts l8�(���q����!0;��E�ʁ�ؙʡ����	�I����b���â�~���/E����ViY~
ls��r+�q�ن��  AT��u�"g{m�&�L�?C���H�{��6���j��:���FtB�ٙ��D�|#�fw )�Qmz��8��afp�0&�Gʫ�h�	��ʋ��)�JY��Ճ�΋����[���k���i�����֤�*Fk@�gmA��{0?
�z�� y���K׈���0Ú��68�v���61�C�c~��c*�'�n��y�FK�ݼu+�2��e(��u��3F�nTcO{(P�{��G7gh_��Ϟ�p�O�8z�Dό�	홹]�q��b+#�aڻ�(���k�_
���R*��.���G��~�〴�(��܈����^G(S�n��M%�젩i��˗/��}O���-t_�vm�SO1�>3�عx�"�?�o�4t���u�D�Ak9�KpT46���,�UY��[dj�����kY�mО���TS:s� �Z?9��oP�1r�5���;�ewLw	<l�� ��6�(�x��L�����$aإp�So^N��5Pw��7�Q�������:bL?���D���vgݻw�����o������)� �5#�/�F��|,͍��2
�~�c��d�;�/�w��0E>'Y*͡�i�d��? �k�N�
'���+dj�9�ɽ§��w��a:�@X�j�+U׵��z�
Lz|Y�B^�'4l�eS��M9�l @�@��וz���^l����>�Q��o��B�`w�b���b��2�[2zf���^�L&�\�{����[��d�����aܳ��/��>���쵈�5�S���d_�:�鄧��;:Db�^K���])C� �~_;\���k~
��X��BOZ)���ĜB�6��whWMۖs73�|�Z[�^ ��lfH�L���;��H���tJ�gV~��dV<���~��0�%>�WL���kV��FIw���FO�+�\4��M�{gMF#��cfӑ�S�2���7�^ݺ�@�����"2�Q�'��ǆ[q~�}Ip.�'!��\�<�n
�W(9]1n����&�z#��PB��y_� w����Y�^\S{��}��B��u���=	�̜�{e�cP?��z�k]��B��g3���2�5I��L�\�w
��I�m��|b�Se�Sm�~���O.lB&4ۼ3�sW��B)؂~y}�^�S&�b�΂�RW�;��|�ra]��i��r�k@�OQ`���"�;�I��&�4H���ʔ�_?�]{�L�1gϞ=S��i�����5�)�E��c&��dcgɵư���84J��N���f���Z�+A!��n�|˼#��n��O�<��}TS���YY1�g�.�V� 1� ���N}��D��5J:8�;� F�b,�-**JW}�N�OjQ�]�p#���x3���j$�A�ry��L�������ٗ%�- �f����F�c?+���M���n��:�U�L�	�B,��fJ	Uڌ\/	2����u��bX<�^<��8$�I�:��n�n<n��%֏C�:a��	�O}��%��G.{4zrL����C(��>_x�+��\�%��I���;n|�{\���~v '�Pz��{��޺�۸؊3=����8w�.'XrQ��p&<Յ%W�o/�c<G̢�_5ǂG���+�yV<��C'��[�f��{������h����*U���o�F��`���ͼ򷙼D,V�ň��d9���^�B
͝ȼ&�_�w��	�\/�F,�	�g-�0��}�di #��>�WRW�3��irdw�H��#+�H��/��N܀��R ��b��(�VG�V	I�y�z�{l��K�G�5d�ʟ�_�3��Y����Co�c�zz��o��Qڈ1$x��u#�C�>����t�4�5_�������526!�=HƯY@k�6����';��)�b�,L�il�VwZE��[O�3��g�7v=}�tkϧI
�<n����~G���΀/@[���d��1�ӈ�|�.S�9bs�`qp��O��Z?H��\/���I+ŀ��>��FI�3� ���`���1ڒ�z���`�.ؠR�UC�й��.�+�@�'����	�>��.v#ԸSV�<�q� ���S����uz��X�{��v]O��f�Z���=����%���*��Щ������������e���}��X�O���f \��+U�:WNw�������в��v7�im1��r�CAq���d�ۘ<ώ<{2Ԩ!�w�ͅe��f��ؤ��/�d�K,y��9u�=��hl��G�t�W��|��fϝ��`�k�`�0��A�l=�+v�}�6����'�JmJ��+U��I�q5	r��E΋�z4�*\[w�'}'��m�o��U;.���:i��$����{��'��w@%��q�{1�s�oL,�Q��s~#�s=�� ����}et�Z�Zw��J�?eKa�2���pGlC�}!Y��$��t!�G���a	�))�������\��~~S�7SRxv��wPj��]�V�{/��`�-�o]����H䅶�]	���DZ�f�;E�h�����:>�&����8: �I�c�%��0��0:%C�7��c��Ka�Z�0qY�/y�8b5Q���j~��Z�h'��!7�%��M,�2�簈��������S�]�ČRC"�6NHt�:�Gzr��y���rA���
�C�A�ȈD���,4u�����e��w[�Cw�م	,��}�b�����`rr2S:�����@�;Wp��#r�l��O3Ж�cF��ݔ�x �����֔V�0/cv
뉬[�=K�ӟ��rҨ)�nXM1]kt�燌Mٱ�P|/������j8p��&茺�D�w���6�(�4�9 �f�#�k5��.
���^����j͈8�f�����B��K�̓�=�v�\z�R+���I���v�7��a��-$�^S�b�*}����>�&�E׳2��%�62ed3�0�i�51��i�Ob]�c}?�<���䥘�>���}f�	�}^n�B�n��o@'H��Dq.�������`x^T��@�?���yϦ�E�vj��q/�܋W��Bb=� ��FǞ;�r/��gg
�'��.~I����k?P��LdVN�eB��`��6�R���K�mb�f.	�h_p<ΜȌ�I�p�eJbZ��$���Pkf�0P�K�"�l��n>xY����^��Vi��l���6.f|��Uf�]遗���n����/��͋���0���r���Ϋ�1,�d��{�5�����+��[H�����		)'��/��a����r+C����ġv�"�������}�0���-�)�lKfhU�� ���r�j����	�]�W#!CD��a��ń�l��D*�J�=T������=&P������U��ow��H!�)O��Q�Xm���|o��� $VQ��ޠ��b�Z����/:u�C�!���[�4��^��	��:�mE���7�H=��/���E}3�J.3���;�Y"�^�R(��7����zP����j9G�&'�r�
.5�~��
�������{ٲ1�L'��[ųQ�V0��a�(�0썝�F�ڇ8pT=�/zC�"7�N[���Q��755]���
��{�]�F�ͻbK��۱�0�
���NK%�����IO}mo$��.���R�k���|��LO�����5l�0Z*
����wPN���%n�����g�=e�tP�;�οv��mz�j>�a��bx���W��®�@h��o�&�۱k��SX0��b0Ă�L������������e�5>�7m���d�ơ���>�34Z�Ʉ�r�fҿ��f!&|�Գ�~NNNW �N���0r���<l_����'���b���!Z"�����b#@l6C�OF\�*	�#�c��P���٣��p��K�M�a����]���]�1&6�X��)�-�v�X�6��r��g�]���Q�|:v�>c�'�}5���(w[��-CB�@"�̖[� J��D��j�%�6�kn���a<�/v~�r�ޚ����U8ه� 2I�.Ҿ}�����m �9�b�D<�:/k��/�EwL�!P�|+���A�sJ`)�� �te��);t�frՔ{���xjZ���shttt8�r��xr�v\g����<^�ܰAv�> ��n���7� ��o
��H��mL�ڶ��N�30�����aml�3���u�]��(H���&ƀfkx#���.�Ef����i �Bw�@�?R& �;6�V�<�����%x�����<�M�L���1��w��;�JXn�uA���g���K��Oa;�,��~%��#V͆k	�h��}�\�c:�j`XgJ��D��_�tu����%ڋ+2��ȉ���*�Z@>��Ø��2�h-���1�g 5��_'�jFt����̣	j�<�w�չ��T[�_>����:`��w�~�u����@⯵�;B���FW�8dn����1U���R�/��En���
m*�w]�r���հOnq���?r
����x]���Sߝ���yݬ�nS}j�r\�J�͙��;�C�Y��e$��!��8�$O yݼ	L�F�;����x�ꗒ��z���~��*������+7{x��s�0�?�+���b�<ɭ���2�=T`�F���C?YB��5�¡=�V���Z3���E��׈���&��҇]�j��z���0��R�
YulX�J��!0�H�z��i�O�g������{*m�ּ�M@˟���bʟ|�W�cV`.V|1gOݒ�%�(����3�B�7�U$�C��w����5�Pi�u��
��B;�5i����M�L]ҙ���������������u�@�s���ߤ�@1f�y�����5~�:�'}�탕��F2�KS2?5�$�oO����9C1e���̎�L�����f���O�;��g>3��jD���*:$HQ�yp�;	�IK���5VJ� ��{[��r��_P��d�͘�:���'��d___�4����19(�C�Ńhʩ	�^P1�>/��P���;$y?����1��yq=QԊ�[��=;�lb]��������N��%(��LA�E��Q�J�c�}�i�\+�3��Ä�z��
G�����au�O͒Rl��q[x9�6u��ӽܡ2�Y��]��OR��-]B�5�\��X��7jrU�8<2�hz�BGqv�+Є�{�k�z�\�2��5�ĲC��Y�:g3Me��v��2�,���Ĺ����Kw����H�var�x�!_�7־�Q;^ߏ�-z=�k�L���D�**U�����VZe��<z}d���xzK������cv���MgY���d���\�J�}|N�����~��}w�cφB0co1�	�Y����2cv�Y���K�M��tp������j���I*�n�!!!�D��kmGH�%<�E5�f*���m@���:l��zs{�y����K��0�ѷ	Ԃ�('�'|�+)<����g��Oz��5��e�j嵅�k�2U��� �_Ǳ*v
����^#f��H����hN��PC�#ƍȤ�X���@��vIp�$��u��ܧy]9		�"s�ZO,&7�RM&B��<w�OM�e�L���m��-C��4,��1��&\�k��]7$�g|T5~y���N�n�8妀�����Ж8��o~�dovv�­��㴋�K;p4���n[^F��%�:�=��H���yM�8����YZ�ڊ�˗�߲P���yyO*+%��)�Js�%��]��6_o�|����MOn��L�����t�ȁ�EQ�x��{�c���E'��'IJ����-�ٍc���5T!�=I�:�5��}�"E�밼�����~���u'�I���C8Qjvy%'�M�5�}%��|�z(�?ȫ1��p�mb��$�}D�$o���]�����Ę�q,�m*�Fŉ
���cIj9��s�j��Ir*��֛$�b���0!O�Q���G"Ӄk�6�4���<Q:�3�$`&;�I�4��7�ԥ<��#������)@��?yr;QZ^�oT�1���T�CY	9�,�"4q���Q�ר��SQ��??���*'�p��;�	b���SQ�}
�V���{�n����Z�[@�^���֋�,*:��=���/\��.�f=IM�J��{�>sÆ�qP��E^�J�[8���#���O#������D�Yq�p��~��q�6I8���ar!�SǪ�'qo�x�l&a��0d�xJ]��cy�jl,9�HA⺈dyW��r�ti`R�h7����������wČi�e�t�f�&�t@ZN��k�4�Xہ�1�H݁���X.�\u�RÚ��]�ݛ�bs�&��ƀ}�*��͏)QIޫ���i�Y
��O����V����@�&�A��9���4�c]d	߈M�$8���fh´D�-�5n��hK"�d0����>\O��m��Xl툺,�2]I�/�7���IB�%B=�z �$�p��0R�NI�+Կ��bh�i�ǇIR�h	���Ƚ�L5�ɫ"��Z��|^kf(�l���	������8��.ryq�/2��?���p�&�w�9� �R��`����.��*{��Y5�/XM�_��C�*��$����$�覠���  x���#f?YiI�Tkex��;�,�b����zJ�)�>�M��I�=�^c�C�hb#�ʂm"-1"k���G��ʊȫ��q��'~u.����ƍ7����]A�զ !$>�J�l����0�t��O�����~���Y��r�@>���Rjm����G�~mmm]-	o1l��E���."W���8c�MC�p�ed�w�o&6i�$O���o8<�m�!V�m��w���Ν��/$�?	NB�Zci�.ߣ�Y�r��J)QH�8Uň�#�A�5��|�z( %=�����r��N\mxKU,�y�=���v8I���V��R�'Rq�x��|�؈kp���4N׎�m��}#"�S%%<0���߲��Q������8��\!����h�V��m�6�#ݦI!~WK�WD���Mݴ��*��ȳHOs�$ʛ�3(���d�K�?L���Y����H؏�d%kV���>Í��>���|��7�I�B��űv���B6~��|[��q`&�*��6ܼu���\�	�9���<K)!�=�gy�v�&{�3g~D�撤t�q�7 ��G���~�&��NR� �%��.�b�A�&��ִ�m��`���C�Y&��:Aʈh���n{3`a fՖ���4rn����'&�>�i�"dnǥ:�;��v�Kޝ�'O>1P������{i�S����d��[�閍9���������̝�+T_Ϩ(װ�&*=-��=4"�!�T�2�:�T��$�aN�����٢G`#����<$��L�.��G�lB��-�]�T���*	��[;��!��W
��2:�pO��HC��!��p|�K�7NVEJi�����u�W��B?��FZ�D��L/���Px&D"Eo)vq3j@,7RU&�>�ΫKsa�yi��m���2?�a�Y�۞n�/�ޡ���f�ǩS�΄=w''']�^�;h!)��h�MF���_<~xc�u��ŻFQ�?~�tɑ�4�\Z�s�j8�.i��(�]��b�j1��*�Ӗ�-�b˦�>˛�Ns(�$��˽;�?C�5�R����Pd�(�겟�͗?�������o�$Y3׍���~g""=S�*�y@]z�c���Iv'X�onnn�Zk����dz��545�%$~��h��!�t��w&�<��u�Z�C����r�����]i��8��� �|���U���O�v,	)ֵ�]Mv����W�\A����ݮ��<�U5 �!�N�c�Iᶢ2��'��	�c�y,��wi��oh�N��#H��Y�� ��V�oDF����V���Z�y�Yic�����V9��D�ѣ��
v?���;�x}^���J>��6�|	���QU"���Y��?ۡ�Q��S���\���G�m? s*=��d)�;�w"��ݢ�Dcp�Ν�tL�3����T���#v����D�0���0o�-� G�����'~�V���x�('2[�qFF��pcC8p<+YW�e�];�|z�����b�赞�

��؁99&؄�܀���/���bAK̐5���[5��e2H�R�Ϟ�)44t�ə�>��k�= kk-ށ@�aR�e�h;v��g۪�o>|�P+�;X!����	�u-H�濔L+�*QhN}� �OL�c���X�ہ�T��{'�!��
Ę�a�0�#.��sU��:����2D"q2�.#+������*]�o��/B+#�dx<��g��OU��xO=�YN͌�E����	��

A���5�F��S�Q��������,*�����ۀD�>G��L�Sw�J?'yL��|\\\ijH,�A�&���"�~���v=�
��X^��b���O�\2���*��@���8JLL9#?J-ph��՘y	m���[մ�ZS��e����L YH|��cPx�!;Ā5��`̈́����>Fm~���\F��G7�� .j� ֓S��$!��� �����}��6�_5�EOe�`�pV��,�ʖ���i֘ �i�JI�9::�/*���֭���6�DG���w�h�� g�u�	Y��x���Ԑ�B~b�XzN|ej�Jr��{[GL��cW؋$5��cv�i��zN(LnI�sL��@��hP� d�WC�|���@�)��PU�[tOxS��,//�h��օ[�� 㝀,�_�u���.�c^�^π���J, �\�����+=}}��PUU7@����{�V�W�
��lSz��|�x��U7H��Ջ#����tedd�#h��(���Pl(���b ������R.�Ҩ �gQ:J@~�
�q���5+��R�zzּ��`T�?��Qw6�(�?=Kw�LN�`@�(۫I����Y�D�l�����BUj�/B@b#����u��s���UTz�.���S���T��>��}ܭ�����R�n`���Χ;�{�]|_J��8P��NV��������s�� ?��th7[�֜}��*P��?S����'�o�����ۋ����Q̪%�Z�J���d��'���0��֣��¨�{�|�pVN��= 3���p%p�,��?�G�c��~���y����������{  ��������Hi����b��X�@E�p�r�wՁ4O����������A����>y�ys|ǡ�WQX����� �Z�bd JK��B����kV��o�w�n�\���u-{��˸k%Ф::bڲ����_=G�����B3w_��+@�;#nݺ�`������y~��[���C�r�a��$�`���~mo5����C�� rZoo�9K����c��z�:r?77�Nk,�6X������W�Ԕ��G����$om��+A��y	�q�8�E ��a[.c��}�!�>H����D0�u��볏�vQ�0��ͯ���h�g�B�Ɠ�0�����v� ��SK�L�Y�G#�w���#diJ_��2��� P�`=V���Z7��E�oL�*!5A�s��X�/\k�G,i�K�R������	D�i4��Pz^eô,UI�U����@(E��a��)�[)���O� a�`-�B�>�-�T�B~R4��"y9	�f�)���i�	�O-9��W_9A��k-MM��8�Є���%�P�2 �ҽ�u�z��o3��VA9��1U [O]��f��E��ٛ�@��F4G;� U�yz����DϐG=�p��s�As�u�Z��*y@�21q�4�,���~>[:,A�jڥ����7/Zo�읉�73c�����k����E {r�$�h�VCړ��I�U�V�vj�kf`U�F�	�x��ъT�c�lA�1�n�3�o߾�I\Ɲ|?	`rz�8绮X�,��h"V�Ov�Ծ�-� �a���e�agg��Pe�֫t���u��9?�$���}�NG���Y@7
8��~��d���u=O�w������Oh��)v��I�?@�;W={13VG/q�*E����W('M>ɡ=@������g���u�"��;�5ѝ=P�����70f�����Ѫ���)�j�Wfǭ��/��I��-j-2Lu�L0��]�* ���	ľ�Ӄ�݀%ש�m�%(hh�*+��H7��k�ĭ�1�4/[V�!纈 ���6vv���X�?�a�Q��n�$�l@�t�իW)�5�;���n�-�!cO�� ����%	M�NB��z��m)��R��C�.���!��D��{)A�g£J� k?�������])�)���Ǖl�g��
���ů�aD�
2U��i���6�b��߮��҈�H�]�R��8Vڡ̬,���.0���7T�t���N҉��Df�H�����r����B�'�����';>������ۈ���xfcqq4�I���,P陃Ue�P`��%�cJP۵�%!R�O�4��H��ȀsF�t�Ò$k����K��~?��\�w���\%;:�C��}����2T�3��*v񈼭h9?�v8�k���sp}���~�uua;6zz�$h����M�%�{$N�DO��R�Lq��Z�v���i6S?B�lY{~��ǜ�ˏ]�x���WS��!�?��c ���G�0�1G�S_���p]�)�8V��O@�lml�� �\/�u(�~۰��o���
M���͸�Z���ΚY��YY
�������7ե����}����?���g�����|�F~*Oc�Z￀�.�,P�����EYr)VB��moVI;fm4�j��g���@��q����s_��'�˷�⦥�.0+.Z��}q ���F�(��2m�S�	���̈\ǃ���2��P�4/�;J]��A�#N5��fv��yg��?�Y+�(5��v�o>���@��m��x��-,�R�'�������{�� �DjZ۹ҫ-Ye2�dߏ�gdK����="d�x��I�u�,϶@����߲f9�_�ˡݽR��e��T��Kx"`��T��g>]����{�A�O�UkhxO�g�KOj��[f*&4M���4����NX!�QPX�<��PL)5�S�OjJ�y ��HNIq�f�#�EE� ����J�����6��r��y�왯o	U6�V�4,�z/�t@O!�P�0�PP�� ��=��F50�,�ݨm�\�%����B�	jCnQ��S;7nQ�>���|��������Pf�o����I�]��ѕi�(z��'f��i|���	�A�w�Ø��&����%b��^ ���j�ZBh��!��,��

@υ#��-�E��^�(�(CrRg��"�&�A�~���Ю���O�g�qu��m
 1l�E#o~D#)�Z&�{?�h��af�� c���r\�"� �7IVA�$+-�Ut �xy�^G���C�`�o�k���eW"�1?uP����w�T����ű�� ����|�f���*CD��]�a�/7��;�h��T@]*�;o|�o��s������#������k(}dI��`��052���c�%F�I(�ۓ�Q�k�$`�ÿdkV�6��m&$~�*dl�+wD�W�+�k�4U�������/. l><}�7�����Dy�#������)�й~��\�vє���"��h���pav���"�� ��k��^G @�`���~([3�<6����9�뮃��S9����Y��O�7B��t1U��N@��5�k�B�<(�`'  ���X�W'�]m=*��R�^�X)�f��5"��  �4��G1��ф���z��oP4��QZ��By'�Ҭr�l50�X�׀Ð����ue=q�"c�Ƃ����/�o���-WT����Iȟ?UiD�j�9�2�
J�r�@���4��������"��P�'ĮO���~��a��Q�
�1!����0���zP8h��(�a~�ڠ���=��D�O���\m���h+��.$��|��b�.v���В�SG6q���D��+��j�Y�����G���e� J�n�?�̆k^�z��)�j"�	�{�\��#U�5vQ��K�_ׯ��)��0O�Mg�Me�0�`�)7��d��{n�D�3�'aK@o�q�=*���̊Љ�0�b�!0��vG���w8D�����k�������&�^c�o:G����ˣy�90��Y���x�-�����	��=���̭��2�Z���*��[�5�/A�T�_o�=����^ ���O�G�W<sZ��o$����ǯ5U3!k�_4[��:9�(>�?ȍ攫^
��O����p�F ���fh�+��������W���^����k~��Ly$�n�\s` �@�=0��s��,�GGyG�)��mC�* �V�"�qB�Z��m���w��a1q0A�:�˨�uؖ��3�4 �/hU������ �r����8-��l�J!22^�4(Y�d+�M�^�SVHB�5*+��{UV��[F�����_�����r]]�㹟�����>���s�l⋞;\c,�ӛ}d���9��B�г�+f˃�r$�X���lV�~�����Q?YQ,�cҰ;ТQ*���R�Bv��/�yyy�'Q��0�m��O��.� �ߠ�j[�����~����1��T�*B�ё���Rav+	27���O���0�z�Y5S�}�1�L;^�3ˆ�)�B� w;���QU\�[Ā�\7��_��2����ō�T�O%� ��#��o3��ބ��ɾ���_� ��y�8�����a����DTV$E�Ë������О�I���nc������9]���F��%���9y����&��f�+�av{��������c̫�vW��t	9�E��'�~<�u�vt��x�<0D�����?�N���9�Q{)^�~��P|S���]>`$�I�ɹ�B��VQo���	���{1�/�k��3:::�/���}�����I l����j^-��`�4128�˟���`�k���@��bڹt]�O�����ׯ_�S�V5���	�CCC�	u;4QUIde��������d���zy
���p8�d�Y8El��
t��leuu3�}	���&obb"%%U\T$6]|�/**j��ډ2J����]W���~�)m�{K����p�J���Vښ��W�J�2w5���Z��Bwإ.Mܖ�i��O
��������VW�l���v�I�17][�n@F�2++��H<���N~d�]��K���c�q&>������:�iu����}��FI���eJ(��&U�k	wn�dV���x�1��n�U9%��T���c�(p/%Gd�(���	;�����wmy��e�L탛�h5��Tt^�re�⩍Ӗ7Y-��˖�l:�^���jְ�`ee%��2	�U]�y"��5{��u��J��ˑ�\���
循�*�P@J�ǥJ$b7!�?���?u>N���2<���L��sG�:�`ĺ�����E����p��)t�,e�X�H�2Z�R�T��|Te��TG����ġ��n���O��4�@a��C��P�Q�!��3�C1m�JDSS�H��*a�FZЫ��g�K�[s��4�F�RŴ勺��7�z���/�G��kH222z�4������kLyQ��(]�گ?-��KY��(���yTq���P��4o}���
�W���KPWv{�wKB9��3<�֩��|W
!q������@��}SS��
���!�f���69g�w�MHꡃ�����-,D������>ׄj6�����.�rN�y�Ǥm�>�:αa���go:a^T��A2����}�D�c
�q�����1q����C��)�Й��r%w�x�>��&�
� ykuyzE7m�@��=T��@�op����Ẩ��������9Q�}q
����l8g�t��o��$��l�����Ə�\3�&r'���ofȝ[Ӂ����𗖕���g%��,�ro�����T����'��JK�tʶ��b/�TPP`������P�p�x��d��hB��V��-;�*��uĸ���F>[�ƍ�s��z����J�?���r��>f�������7�A�nB��]����3P�������m~�
�K�ӗެ��`g�����oE�-�]���>o�\�7@Q���޹��41z���YT�Pq[|�+���w�Q˳1=Q����D���X����J\JN���W�ޮ|��,gD�?��(�ɲ��Nc�zո*dqn��X�N�h����ڧ!�Q��w����CօG??=@��S��%��>���-C�%Y��9Q�+|}L�Vm�x�8&��(la��D���q>�}��5��FȖ	��GM��}%�5����b���;����i=@��M\��Tmc#��t��ř4�^^����"U� pa���k{컬fq�&Ϋ�+=��8RL7+,�IF�{466R10�LLL4�%��(�L~���rW�4��0�+�nß��c�]��g�
��sW;,B��E�iM�}�:M��
h��}0����^�:��Ǐ�UVS{θ�T��)��w�������?J]��̉����e�D���l��ᆠ����iJJ�m�~��b�U͔��x��տ �N1^
�̲���`y�*ȡ*<���I�pZ؈���r/�����j;8���mA�ϕ���o����*���A�-�����qw��(Agno���x��VE���O����(��R1�u�gƣ���!�F�X�t���V� "�g*8ʼi�vNL'v� 5V˱����x��x7hG�x������@�eϠϹjjo_�/v���|�tj�:�����C�E1�`�^���(\7�}BJ�p�XS�������������o�/��0�2���������s555|���&f��V6pbҘ�w�v� ��@�vo	������?{�l+����E����ܐ;�'E0�y�/���{��#C�����7x�;���+�
(�H(�lg�%Х�S��u2
�d�����a�1.L)�w��j�%�U��M+q맷���WVVD�#�ܻ��|8(����A� ��N/���+R ��w�ې�n�&^��ݦϛoa~a���Ԇґtt�=<<�&&P�|����[ $ 2�^V��Q�at>�Q��N<H,�G��sssrr����/�;{�w��|��5vwo8O�h"���gA��~ӈ��^@e�`Q �/S/��UN�s��%�39 �nBn��J���;��:��)���3ww3C����8�9T͸��K��M�:�Z�ߚ��`t�]i�Hd`F-��]�cQWW7]k������x�J�����&Hy\$�=C�4����@��;T���ۑm�\P��`�kbW���7�7�4�x�.2��"	ג�=���S�����H鞞�����n��L��5�U`�a���d��m�S��o3�5��S��-#?�~�
�500��� (;�D�UM�/utv��O�� �FA��s뼽�t�ҡ�C�ng`` �Ծv�����M����Ɔ/���$)���O��]��k��nr��3��Ҋ��֒�Q��bW�p��5Y�^Y$��T�p�
y�n���;w�ܷ� �%�e��xҞl���:���E2F�w��qt����{�yB+	�ʊw[��/�?��,�0f�|E�3%�#� P�gϞ����E��1�3���|�ŉ�աx5������@�>���Z�#����u���wܤp�*ou"7�{�M��4���M�AJ��������Oʄ�л��#$��\y
-�z�����������W���վ����	��,���_
��I��ʁۥB���셬�^R��ɐ������Qo��8���1�nX�؍щ��͛�?�K�����:��W�Ǆ���nN����b6y%�5889����[�w�Đ�>zmbd4^}��Y
T�/_8ED� (N�%$$�#=}�4�r4pt,�ﴶ$�I29��n3�V%a[�E\��&���V��>Q�X�ӽ��`ue4a�;T�g���C� �_`�`�(j�Ns�Z��v$��&rbk���ٌ����' ,,-K��"'M�~+����{'����jd��ݏj�Y6�?�l���[��x"oh-���Aac��I  3��[0���C(�}�����|轠�`�S�Ay����2e�<~�]��{��FGW�RV!'�A�����!;�=�%�jW:k��8\ы�Y�񣚔@�@t�c���+�"�&b#�v9��pjh��f�o��^�w�$��������|cWX�5�Hl��9.�&���v����E�8߬+W���e��D�B�t�����!��3����}�gΏ�#��O�s��j$ߖ��o�D�-�\�	���ZX_OJM=|���w<Ӹ���o�=((�7XK��0��Jo��@�U8��P�;�#��ZD�u\�?��>�{l��Ī*^��6hN,���GM�+immMX�����7H(�HK�O������2������ �c/o����v{��������.M�Ak��5�xM����,���[�i��ɫ�iQhPVn�E�$Pr�M]�(p��p\�h��QPQ�L�6�iRS{��T�+))�a���8Y$�k,�\�ZK�g������;�*�Ht�qT��W7G���U�G��0�3E��^+P�����ؽ.d�YYT���(��w�MQ�F���*���������{���A9G�jNh(����zH���q��@�'�$�6�+��/v�" P�Zѕ��
�}�ɯ��<4�}����*��E�,ⴚv@�JJ� 
G��T�B���'�AA}3���G�s�E?i�uˊ,?pX��E:]�t8_t
�n�3�*��@Џ�͋&)l�V(���
12�"{�H]8��)�76�J��"!l��U4Bw8�y�t�#;�|PfGZ��-�z���E��"�DD6b(����A�8&�re4nn�)cV�@�Iw��H\L�pL���*�qd	H$��sS��6>�d�e"�	�)�e���!���P����8�@��
ٽh��~���P����%I����*��RQ�����E��Ӽ�Ꮤ&O���J�� �!:�Ō�t���%%�A0���l�G����ܔ��`�#,�et[����Kɓ��D������n��I$" Q��Ĩ蚛s;M{i��Y(�76��҂�C;�nP���Z��J9[�g�ys��$�&x�ʑ��E�C��gݗ�A=Z���7�)��co����8���84}���aI[�,��/�W-<V��^��n�y�51��΢���qT�/*�q�p�>e��ԕi�)4]|��&�^d}��b'V�f�-_VVW�PNM�fCk����n�)))�E�>����{���D��<y>�{J�o��8L��������Z�a��d������Y��#�[a�{�w�WƖ��^�D=��dٽ���g�pa}cjj�_]}�&֘746��Lc7N�sv����$����5�܅���W[O��R�T�KS?�+���&;on�;,=�^Yi�U��o��		��/��-�.W$�IQi��*�Rhu,U=J~�:�q�[CY�*]BSSs�c����ӭsK.�����V���7@�A=��rC2�"�C�j�А.�����c���Uv���*�!]�Ųq�iѫke�?A��[&����������θ�*�)��E�$����@���*�����Բ�΀c��u��$�i�D�Бz�jΊof���C�8��ބ&ˤ�x�Y�gXXX� �A2_���`��`�k�~����겎5dP�ۺX����w� w �Q}z3͕�&��z��2(\ˁ����o�$A�K8;;��a���N>�Q<?ڌ�F�ҿ81! `i�7���q#`+o�����.���'�Ք|�Z/ҸT���z˨H�_TTT �_�:YȈ� Y�񶎎�qqqw55}��;��:<�?��F��xd��c���a�N�-���5:hk3���}��sQkmm��\D�{�=�Up6�[������Q*0O��Yr-���KI �����g.����|�!�vzF::̀��p����Dc`�&7��z�L��@~�ZKq�� �������Z&� ������o@�K%��zO��v�D5v�(����g����ϓ��"�jI&V�k>XEM��>
��ؘ!T3-���B����o���`A��=D~-� ٙ`� ��s�� ����^�`QI���h៬�A�B2@\z}q#���At�8'��v[��I���w��J�f��,Lv3:::��0v6���x������E���6���$b��(р��ST�̈́�I����;�P]966Vܙk����P�.B+�u�Q�y�)�\���ML116.���s�x�8��6K��l%__%_�s��,iDԷ3)YY�H9w��]_?�Yo���W�Lj���)4�Q��%hC3��6.�H��b�� �M=�� �z�9As��+�m��jl��@nף�H���r38��6w,��G+��>��&5$��t���=n�_:Θ	P��F��>
�x�΋?��4解�a�"��螁ktt�[�:��X7T[>􂔨��v�JH�e�{�ZP2��V��*C�c��i�хJf�E8 J�M&����ʥ�/�} Pk�����ZZZ'��V�Gwm.h��%ݔ�i��@����P�������u��Q(�4o�#���Crj�?�4!����R�[����N�"�� �v�B�Eڊ�L��l�9(��Pȣ���\\����&0h<,!�r�l
�MT��8�7���ɀ��ז��W�ve\`W��4�{z}�z///�)��Ɖ!��h�A�"�9�epx�/�`�ʊ��Qa=@՟��}�~[�\�E�� !턷�W]N�`"tyk\h
ncf٘u��2����ũCp2��`�C$c�R�jp��8�%:��t��o	�a�]#�����.��������h���{hӾ�����xS10TU�?�Zp��Y�c��Y�r�X(f�[oq&(����x/AL+q���}��࡙��J��?,���M� LH	`r"	
R�č��5vo�v�ҙ34��08E������i�pь��_4.y���W�����1E>�*�Ϗ��OG0UVU�zqPm=MĶ����:	#4]__�мB.ٗ�l����0RH�Dq}kK� �! ��e�Ƽ-�����7tn2Q㍨�H�t!+��S(�FH��K�� a�U˷ۡ��{�dS�������a�� �����C�K({|ᆝZ�Я�$�ddd$�Ő���@�+q24>0�����|Ң�vU�����1-e*�F�{���A���&��B�8C�{Od��y�6�A�$k�ՕN� �w�����<6qS�=;�5�p�����������#�T
�ךlik�w�������#��d3���e������0b̾��@ƠG	=t�٧O���ǥq�S�	������� ��*��:r�9��kME�<8�
��	 p'(�!(nh�gv8u��~����V^��&B��^�s�NG��~�kJB���]�r����G��i�j&��;���w����L�����_r�(䏉���j�!�P텄j�¸qqK�O��6��g�F=��������넥]A0�`4��]:�t�x��IgǺA���z�����o�{�#�/pp�!$F��Y:%���V��dcamSu�� � Ը3��C"N3ҥ�����J�7G_A��U,�W�p�Ҁ�� h�t�G��j�M 2(!4V�{�=U�z%8Eꌻ����6�
k*�i���̸��ͣH�C�HZ�&g��K_b���l�TUU5]]'<����ߗg�
�����g�3e��=|SX�t.o:��32(�f��nQ=7T����		%��f�E�6���iP�}NK��yP�W���3�m��r�"h(���Ω�O������?A�CT�,?1\7@�q�	c1(W0x���cʢ���b���áw� "��٥Y��\��V�C(m� ����\�=zb��q��Q�/��ǃ�Dϳ���r�|qC�A��<�5�,�	x����?~t�E~l�GJ{�1���2��lmQ�r{��q�K
f&���@#֓];�最R<]Ũ2�oCn`H��yl�N<���E>V�V���ٞi#C�u�z��j/abbf�=Q-�0������lcG���6P0T����l]II�Ɔ��iW�	?����c��W�[A�11
:��=h~A@ݗഠ���]�yn���_���6����'̡b"x72�G8I�y��iq48]�����4:z�o���;�Z::�v��/,�]:��T�����ι��a���&m�3���J����9��.Bq�t@���|e�W�J���}"��<#>!6�;�AGb�1 *�ˑPgF��@y�:xSD�
��-yQ��`8��/#��h��lg�/o�Q`K��"�r����֮.(R�x:1�Ah 9Z���q>Q�B�m��> ]q��t�v<�������t���ߒ��M?Y����� V�����Bd�\Aq�GNJZ:�
q�!e�	Cؗ� �)(���^dm��z�s9}�yb�|��볝�vTN�w8�|�����'�R��d?�v��yL��(;�h0������
�1�r;Q�VG��V5���e�����`�F�2@6�����#uޔ��#P�28l �L&�\�v�]6GX7���:+?	�9�!>��I������QU`u�Hcvv6��{���Qȃ�Wv�3U�;��%���颭%������+�����UWG��	�6�o�����)�d/Zлv�?C�=��;bw����������X?uxS���+�|�SC�"�R��^\II	hN���{@�Q|a�؅A�I�����j�F������L=�S����}���L���1)���jW�.O�Hc|rZ�+lTz���ϲ�s���L)��V��b��:�m���2[dX=�%?�I�M���^j(�����kK7�5�9����][�1�G@��M�j��I���d�����.���Z�ۂ��:�U�:+++���$+�����7��B�=D��� j��\_T��qW�c��V��O����p��`1�b �a�I��^0�=��ȢP��[Ղ�&L�I0�5%^ǵ��7�~��%�!1An3R���`��vA	h'4�@�L��A�|PSOrC8�^��h��07���iu��`�`ܑ�LxAgҗѷ��J�`���ҁ��oϚe��"��E��%Z<z;�Su��<�0߷����9
&�m�=�S{Uh04(xW{W�-�k�U���v�CGS���E��~zn=˰w� Q�w}*��Q�������
��eTO"](X��@�`N���?��bN؞Y<��.3���٢w~t�q��7]����)�Y�h��l8_t�A��N�?[L����ڂɦ����K\�a �-���g�@�CR�[/|�1TC�3��bAae����ˊP;::�y �T��,�qu�&Y/���n�uyC�7V'c ���-^X ���ń�`�f��`3���3S�E$�X��j�c�z����e�j�۷"�T)�i���L�aN+�H���$���E��z�4�ʦ��9����mF���G��`!S�f�����Q܎��_���=di�}V"�P|��B����o1���	����`9W>�ss��1�]J
�c��dBL��x�O���t~���Ѝ�3���c�8lQ1cj~�Qzd$nL/�$DBJ����'�@oQgΞ@z����:�&��_hh[@$:�s#�v��?��/���n�-҄a���E�(y`�kQ��L\`T���6�/�:R�ܘr�����F�8n�QH�'bޭwn�A�6���7�����	��y����)�蛚r>��!<Su��uZ��@����B�JCK��ލ�����)���1aD���7�`��"�G f����Y�}�̊i��VV����`?�8^q�hw4 �Gc��}bh+=�����Ӿg��7�@9ޖ���-,("�8��-��
*?7����`s��MF��Aa�u�bkӑ�8�r3�Ss��(~ m{{A@�ʔ0�+�FX��sp��J�s]����q[b6���*�p
ӣ�%oB�N�#�>e�u�����Mq
1hԱH����3vqG�������j>���~GE֦�4���+'�	SfNNzr;������B��ނUP�����
�|!	� %������c�� Z�P�����C+Js�����"���-��in�'�m ��뾈�^�i,�7�&�B�6�މ�|��b����n�l7$f�O�	L�
4lpp0A�����^�8��	y���G�4�LD�3�)��Dm�#������C£84)ݍO�:�����_�gKF�Vzy���Z�ݽ2L���Dg�ـ$$�����S�����L9@}^,�>�}D�A
� {#��P��ܝe�%���z�IP�;%�uza.I#����,FA����[��$koF���1�K5(
4%'�����(�֢pp?�.i�o|�V$�UE�	HjR�_�p2��r`���]@�-�346��)�wuuE���䡥������XѴ_�5�ݼ~G�9x��|�|Ԓ�N��%s��|A(B��ZQP�&�]�+*
p��x��H�x�E#a ��(񥗠�A��̘A�.� ����h_ƴ=�SOwC���#Z�0��B�!��V�-��ZC"*��^�03`^x���޻��{_�sy��sg��6���PЮ�**��=F�����<$1�@x����&g�R�����D��A�:땶�w�G��X���p�&�̰�8R^3҈3�AAڶ���&=��������Tl�md ��9��NdOLL�n��7�Uc/Csä?]�x�B�-�\2?�G/ds�r���Ɣ����]��&$�/ɛ赌���������j�?4�>c�!�R
 ���b����:��ZrӁ��-�~J���U`ܝx�Yh���=_�T&�]�mA�>������$ㄟ*�UȰ���dn�"��Lp@��i��--KC�7o�D/>�&�������;�������S��cbb�^�����(��			K=O�E8�ߞ�V�*#����;�V^��GS:�K�-��-YU�]���]7�N��|{}���QVzU�#�~8~��D�2f���#�q���<Ӯ�/:���VKb�]�wN��J#O^��9�R��(u�)���8�f�j���d��1k�������&IO\��+HxC1X���|�lZ^�×U� O����YJ�V��~%!f����!s����u�?>nxv9R�wJ��<5$4�a�B�HFr�q"�㈗_��'͹�����<�#,l�ů_F��󧂌���J�_^�����mV�^�����)l7��Y��	�:%����2��#��;�Q,-��AC}}�9E���R���s�D���(:�����F����������. �X�y;;�.��E�(��� &�����9����� 8E���0+����[�>���hh4��}Tk���C�!,��9sm���T&1���<��I�}����+`��>'\�!���9���w�X��X$�e�������2oE0 &��e+(;���8G�=��P�F�al�ii�
���Y�ZM˙�9��Q�G�����Ճ�SZ?�C����w+++���#|]YYId����Pv>��R:��\"�� cmGG���̔��_500�Vp!nnn�� ����o�d6�p���b@�<���>��k-	b'"���*Vy�s����&�r�h���ݻZ��-�RS͕�냥ġ�E��K���e=-�$<����J:ndd}��r.!_\�ܐ�f$<��(uV[����<�r���b����~N�mX�	�?������/±��ۥ�����t�w�@U� V>�~R{���{��ͳy��0�R�`Y�7����[>��Z�E����r��
'�ko����,������Þ�4�,**��"L���3_��냙�<�4f��`�e萷8:�þ|�^�L{���p���p{�T�պf?�����c0��g�.������f�ıCE�o�n���T���fA�<�^��$K,�'���|^[�3�� j�`�[gfR��
D�WF����w��
���=�,y�����]���(aSuk��A�0����B��������8���5��H�����}2��q�Q�⁁���X(�R�F3�����H��066V`�J�ipSc�>�H�mu,B�������l�Ν;<�����onEɃ��x����ZJ��T����zz�.(f�j�-_e|���(�$o��ڍ(?Q�jik���K۪[I�����h&$�����`b�0��>�ty�|g��٥���7��N�WC�A���::�~85�iMi1�)�3=���X��r��X�����Ăg�I�=�{�;V<��c"���xx��3Z���Y��\�P}##�}�ϒ�k�8���LcŬPeUKh%Ði{[ٜM���X�n�3G`Q
�����_�lJ'Q�����|��.W����Y��b\F���b,��=eF&&�S��7i����V|,GXQ<�g���jJ'��gS���/�cYH���l��'���se8��
�	M��Lz"�;t*͆h�1M,.�rHH�~l'���{�?��!���ĳdگ�����x���KJ����#ƬY;f9B�4�/�7�hVh�"��?6�R���5�[���v�r�dJPv��]-��{����n�Y���Fo�f�O��E�[����
��χv�L��Q��v���6�y�7�j�R�9gBt���H����y�`��U�Mglk�>��턺Ї�7�� n]r>_��rHܢ�����j�E�;�}p��풀@\U�L���c�(7��;q��-3RlON"t�+�(2Kz+(3��sT?�߳9�B�q?��ˋ8W��i���tK❺�f�S6G��o�'�&Jy|����~RZ��1oIW��t\�}��ʧ���$�^���,$<[�l��*I(���+�1q��GM� �1�������
�Xa��={��+> @��̛��֋�x��xE�������QKX�f�5����8"3]9�)�7�5|�'���K�^����w�ry�����27�K�=ε�Z�h,3�z�K��#��ŧ�Y.5EMA�Cu�v��b�0�ЍL�ɯ]*�r#B�DU���$4��4v�x��rE]HO���Y��Ve��U˝����T�Occ�������P����d�Q�q�A�h醸Q�gƆ���#����2`-�B�����uu/�sV�a\�+�z^=%����~�\PŌ��n��%��O�J(3!������M�~`���m0���*-}v�ϝ�l�q<#�w~nn���xbe�p�imq�O��I3aAA�fK�������QQ%͗232(���C�1�HK{��ff����R��Y!�+�UB�B� �Z:b�j������}}}�P�f1�~3i@����y[;_&%-M�������sO����{���n#���
<?�A�C���&Y��h�14�F��$c�,~~���g�d�x�ӉB���^�G��ѽ���<�~�E'?�dd<����_�6�w�����3B�wI1</��-�o�$}����'�aY�����a� ��.�3"�j������!!\"�V�-3+r����dv� d�N����E:�cUmKƅ h\j����)]���А��DOu���XM>2M{�\qqq)�s���?_#gR0Q-�me�t�y>~������%�j�Qo���7�5M���O��0d��� �ߖW{-��Op�N�0��HMMͱWic?�I7��Lח}�ʘ�(wn,���7l'�	}!Ng:�q5-9�� +o��e��_~����~��Pu}[[��I3�y�t�X�(� ��|E+��e#��-H��2�q��!!3a:��`_�J������ᣚ�������ZFj211Es˝;
E�wY��ExJHT�R�Z�H|�Qgć$]=��k����3t��O��J�s/CU�c�>|+[����d�b���0R))o����y]���̓` 𡤤��I~�y�{QЛ=�b<��l7�`�끽�j��8�sxCo���;���W�����*��c?�0|?lÚ��-�ܪ�lho��;� Kl�c6��V��o��_�43��:��
���ǧ�'��K��	���{/ji��T���MN�n�z\}О�A����v���%z���=���1�%?ٝl$.����%�-�$%�ؒ�\Z�tc��=�ٌWIJK+^ĺ<�iɰ������^ ����=)�C��SU��!�#�~' "�Bt�14wt�U�=��{��=܊����E��b,_mQz���x[=�,*���'�5��5�헬S��gz�k��\��Z�O�o*��L����(�1>Cup�	�Z��su�2��*jj�Y�.��l���c^?��~�.VGS���I�s��]S:$D���1�P��{��q��o�C��c9�E�"TTU�u����$j� Ny��O�R*���c���bUkfr2���LHUQ���Y�-������X�� �ђ�6�h�,ls[9�X
uuu���.�v5]Y-p[�<ǋ#Ɛ����PQV�[��a��ߗ��i��6WW:p� !�&p��򰔙J�D��7�A`s�92�XA���ܯ� Ì�bqw��>����FNN>Z�:��s-�eb�y���WC�z�y�n&�
!ޖ��2��G|�5��F���R�&� ۗ�B��AvQ�6�h5�<z�訷8�a�A��1av���v����(��N���u��0�[�W�[��:��G\������=T��X����3g`b/@w BS�a	�G�={�bgɑ���N\�^4����qk��F9j�2vG��lI/�:�ى���3� Rd��樨�7�;�����-����n �PU����Y�9��D�7�
S���g?��1��wR�  ���|�I�,��]?G�'�{̾�O�����W�%*���s�/~�˦w�м�̃3��Z��kM��~|$l0�k�n͐����	���j�1�.]�,3S	�`=::����Kz;6!A:|��y.�ı��+�a62k��H�],&-�+�����D�6���q���>����w|��ʲM��SO��W%4f;��S&$�d�L8�����d}�`|�yv~�n��E�z���5�|+^ �g}6�:�G�
���=�sUG�4�V����qT�dFr��y`� �qxlZ��y\��RA��u�1S�6G�Ջr�����i�ή�WՂ��9��'��7_L�B֗\	����m\��􌌐�i�仯*�02*�����#W'59
�R Rï��%�pB�/��Ƹ}�0s�on�6\5�>d&R!F&��Hl�]�/鞃Zos�x�u!ܸ�o�?��x�Z��̥���ӳ�C�p�L��m�5�+�SDY�F�%�V�nt�^\�&�7��*�S����It�� ��3l����0�7�yp0u�ǏPF+�uD�R�S���6�ӻ��_�g9�](E"�� N���K�(�QW����J���<oE������
Ik���CGSf
V����P�ƶ���w������q�y�����*~���J��kkyH���\�f�f�<X���p2|ߵr�V��×��4t|����6@O��B.�`�=�'�؆A#��BTM�	vԱ�{h�|�^t���Y!#C�!@HPٷ؛���>��>���Y�Uy`ֶ����R�p�\8W �dӊ�/.�}O����1�w��u��A��ǽ(�Ӻ�~ԡLZ���`w�~�|�7�G�$P��pݙ.\��v�Ú���� z�6@���?;��-��(�� ��*?���Y��l�8]p[H���P^^~�مG�� R�����'����Qt:==J���@�wɨ�؊��賎?hʁ�>�wH��7��ihQ��`��U b���7N��I.��
�
��x���z1����1冚BIӱ�b�L9>>Pﶬ�/		IC}�;�Z�C.��]P;���'�[|����?�Pt���6w�^h�7Y��4��J��@aP?iE�42���f������94�����"C$s̫����5�P�=��õ�T^e�c�6�s�IBd���:멃H�(��ݶ��\m�#,Ec[��f��|;">�f��haUO��<e:ؤ�A��n�٭��D�����jV��<ƹ�p~Tj�oI>���d#�xЇA[`/T� �vTS ͜>\=un��=�{e�L��n�}�ؿ��fd,�?���^�% �t���t����R��>�@��Zu��a�=�>�||��~�~ݹ%�Q=�������kk �ޞq����G��\� ]4Jq���>~�f� m����1�e>q���4.���$�%A�/;���-�(9�+Y"�F���Wv��ǿ����T��T�v���'��!��Q����ʨ=��EU��a:��aYg�)l�� |A��~�晓�c��SUEE*��P�hn�#%m�_��+�H�`"��ӬPĽjW�)��݃q����iA�x�%JF�g�
?16.�z�
�W*��_`AD�97�f�fte�5��nq+��4��>��{־8Ϊ�cs��;x� �(a�*+��LC�����(��L�Mx(CCG�05�Ǯkl�w�p^+s�� b��ydhbb �|iee%j798D4u���<N�\���ڔ�Z�^N	g	"y��2��V�$�8:2���/G�;\?�r������䍐���J]�\��JKPDS�=H���ttb�����+����A���H��V�RQ��V��32x�ϷD)��i�X\��������	���t��:���q����4�,33�7#9��F�j��>B�e�g�&��[lj�3?77��xϾ�扣,�_��4X���

D�+4�j�IH�h�#Ӳk�;Ah�!���e}PD4��
'�����y�"�GD$��K�^�bOG��J�����%���9p|�8Ey�4|]�j�c����b���[3,��K���z�������ߔ��M�{�����3����~�)��gc��隙��C��n����-� ;��:�;_��t�{�'���X����Yɶ��|�Mgg�ys�8EH=kh%N&��>��]��Z�$OG��ȧo߾��6-p�)����哖�� F����~Ձ���F��x����,������}u�6����ҫL�r���@`��0񸆍���K@�����v�2�r
`��ǈKHX�-���uu!������Y��<�@Nb���I�.y�ß4���1I��¡q8�ؔ���@ZP#f�t��d�ț����T*F�W��~ffƈ�ɪ�����R��"�'��E�I0KKY�C`�94��3�OA#
�ң
<T_z����F󬭭G���FFF�4������ai�gb] [?����ly���8���|���D��b�n����\�ڐ,�a�����{6��WU�&>F6�QlƧ�A��Z�S����J�rq�IF`i��h���������}�ͩ �vA��A3 h419`YX���Ң�x�%i�ezJ�Y{ُ�Gv��u�u��q���4�}�MMM��u״C?}'jp�E���68m�LzON�OH���F VUU���N����r�΅WO�d\h����$.���\12<&�L2�|�x��9�ү��ik�
iȻ�R��������~��O�������8��k���ݸ:l�fAf�V��@w<M#�ZF���$$ܰ���MM�Zu��6F��Wd�Ӓ�z��LmN�������l�hs�Y�ǫ�LO����ұ����]��c�+W��ɷ��%�=����E�:,�,V���?1��n�UoH���y�з8����O�������R0k%!!qe�����A�ḻl`@���
b$rҡ�IG��bvu\TT��~�/uuu����ڻ'��h0!�~��aJ/`r�Xz?u�fJi��F�it�̇���`��z��z�����z���Y+�q'�f����$]@�(J��V����@{�������S��[}Ǵ�֦˲9M�ą������h���M�:##C��Q�8D�g�v!c4�b��(��S��������'�Y�W�G�L4kj:禧�)s���p�l?��gI�'c /����Bh��lR�D�� >���*jjBI}>�Ze��,r�[3@f��A^�L	����]hf.q�{����걖#�6L6��LY}�|�PW��.rB�k�-	r�\Xe�~�嘀S�)�0E� k����-ӳ�����1ܸ��22ζg���t0���"V�㰇����'O� �&�Wy���nl8�L�>=p���ňµ�BE4� ~�H�ݭ������Ϛ�v&��m��}���N� �AE����3�>}cy��.��W n���r�/G�p��s������i�N���7^o��E0Q��M--w��+��$��}U1��Ū<�姃��7(�(nj�W�����h_���-	�~�*��lh��,����� Ɂh\��x���3QM�CKg@�31.��lL�v��Ӥk��NG�>1&%����>_i(�R0��D����c�l��E�S�%me&�㝌�{Xb��u
� '���ƙ/�7iL,�&�ھ���˅�m�s��M�)���9Ki�ugc�˛��I��v���O�#<����MXA�B���8�c`v��Z�2Ѓ�͏������ݛ�ݩ��Ȟښ��q�r��呋���]	_���X��?�/k���)3��(��:������K��(�W�]޴Z�=�š����/*��%~���4:ON�}5�:G��{�W=x��-��t���Js��R1E�bb�kIN��Ϊ��p��{��R��+���xn����t7+��)��:�9B��C�iA�ZN��Iթ��̙��#C�R�y�������ЩE`�ȍ�±�b���u��/|��e���o�W�Z�C)�;X0�J_�  5�� �Y`�~�3$4Tz������h��&K �x�of�UV�L;s�% 5r]�}hd��B=�]�n�"b��ě����^�2{\>XO�/�p�/?������U����m���LV�] MEG�7XfZ]$\i{h�'|~qq1��V�H\2k:;��*�R�E*��C����ݬ�L����$	�x���_I��$VT����Sʠ.�}��E׾�6�����=ˤ�b�D�`�=�5|/�+���1�L�I�[y��/��~��(9qqq�>��aVIN����q��gϞͭn��t-�8/9~��)�[X�_{?�;)��`�A���­@&R��7G���]D~�P1��d��c���j��xᝐ�d*4�3DQ�FCJ�y�H�Y�n��K���hB�'�Y�iB��V��Y�J��.=��ο�:�9���^��Z�Y���=��ֳ�=��{�+�ӢEV����v���5h�::o";���^->&�d N���(���i`9L��?$"�W1�궏a����e�p�2����cv���N�����A�d����eG sl۶m<�yB�m$%�RF�1~~���N��iݘ��^�N���6�6�����Qm�~� 3"U+KK}��Cɜ^�|�wl�2-���
��n�_sm5�+R}~?ȭ]a;M���խjo���fXW��D[A!�� L^����✚o��C��1�Twg�h)��F���x�cn�ea3��V�ͫ�@�VS�=W�1[�6�(%Zn"V_V/�K�򼛛>T�ϕO��+v��!������י�������Q]�n�|�6H�Fz������|R2�x���2�v�{&����ì��/[��˫ԥ�ye�W�F����Tl����/_�/fa9�A��ݗu��X�=���@�� /�`|L䤕+Vt�F�}�m2[t����П�����!Oӷ�^��T��[�04���-U d'�t��C]�Yx���tR��f�J�)YPc5��@rr �̲]k��������R�ng��{�3г���H���]g%+���S�{�u�j���˭k��]]���
�9h���Z��~�E����P��~����$~���w^$RW[��������Bo�Ϗ��Mǖ�^2[��D�����?��u(�ſ��233���}��-fƓg��O�ך��>�����k�j�|�{��}zTz� �s5�U��?,����W��N���ލo���{{V-	R�q,Z1��P�DD1��B�T�#��܍Lc��:���+<�r~Oˏ������'O8�
p�y�n�֛fK����Ր>ׂ饾}T~�< h�@���C�� }3O�)z&�q��А���t�2H��7c�x���~��x%~�b����YR2��G�o՗I�F�˺�B��S^��`W��y��y���䏐�t�SP55�L�v�.�1~�-2 ����5�e9�YR��J�*�|G��l�6�Ns@MX����Ǫ�Ĭ�J����t������t�LR}�uѳ[�����,���l�	��@1ǽ����J�>FEw%V>���GZz:��C�E��8 ~�-�4褗����ֶR�_��nT��h���UE w���]��C?�!v>�n�d�C�k����z��s[��1Qo�<�5��_�	(*.����1V�t���k��FD�����O%j�/�@�K4f|||T
A���6��/�Q�XQud�\������
���n����@��-�IH$�%8�!*�9�uq�?A�u��	4��ޅ�S�$C�.�_YI]��g��gQ�@�r��
�PV��{M5�Q0�1��!I7�NI�RɃ�6�<�x��Zvvv�/���}�C�����QTTԣӑ������^/�7V���T��*J�ض�O|f#b�Zy�X���Ǡ��l�-�uu�ϕ� U��1����lr|�%ϽG��*9�����p/��}x�T�����>���Xy�&�h���l]Pv�\��#/^SZ�@Y�~�+d���t��0ק�Ŭ�[�8B��f͚5�����1�9�w~������Į��a`�i�*�3>%*3��~��Ԃ��4��*�"�MM�C��#TK�S�k�轭n�����\��U��J�.�jP,�����h�։V�ǿW�k����sr������f�̋-^[�>8%���f���D�V���!��_�O+**Z�b1����>�Q��_����g���v�C�~CƊN�_!Xn�����Y��uTħ�R��6�{��,�11뇃< Ӈ�QBq�q�{������X�<=#A��錭��!��#6�t����]>Y�4���W8Q�^	Y�E7���}���h��4L�P5�O�$�Ƞ:�9G��h唋�%nnn0�D"q�3�a��q�l��~�ePYW�L�ʚZ��ѥ?'��Ǎ�	(��z�<���q��b��:!��W���s�b��~�&7-��OnߌMi,פ����p��aze�U�.��¡L�	M#��F����c\��3��4X̽�Ƶ�.����V��K_��ж��w��&��{Oʏ�ܸq�WH�`ҟBϏ��|�����/���R�Fs�)�����r�	k��N�x�.�ĖKL "�F..��6q:,��z8��v:�Q��j$u��W^VG���t�D�}}^���܉k "��j7�?���ac�n~kz$�Y a\��Ũ�N��M8���%}�"�<�Sh��{�)m=@�κ��)��ҥ�k<�C�^�*fG���jV�����-�9@�E����Hス���ǏAm����Pz���Jn���#A�۸iSJ��j�i�Mר�h�d��|���e333Ә)����l�t1wN�w"�a�b~�g�t��|����ml,���~�4�KxB�m�-�ߵ��$~���c?��������=��|T����J���b�}�>�C�9� YR�k�*H��
���g'#����աq�.$���W�x,�VRR2�i���]5���u�t"�ENm�V��4�����g��p�Ѧ�"���8�)Z�B��ӛ�>��?�.��f��:���:�O���)�Sh/���=�����|����1�
�A(Gs�����zgQ���^ul�,9�n�~�0�������B��Ç����l���4����*n1{��C w���g�
÷��]�v�*���*�~|�

"�km�N�u��=Ŝ��,t$*�������,s��kEa	��O�v�:+�$m��o�}���ѱ�{����;��]�Gw<W���C��mrIގ66��Y��=i��:�H0�P<:s��`��dS&��N��ڨ�?1q���;��4�B=[���˗c�8�0I�"���nڅdY��q����Έ'O6@�������]vko�e�R@�I���*(�7�Q\^o}&���.�����H�S�5��Y(�])�}5L�iP���]��#;�w�ccբ7�~�Dgg��M�D_�h����RHTsg@�|Z�WE	 �!�"P"��\�vM0*H����6�F�_�<�o$���E�P�qM,���
*��+����&)�+�W�Y��U�F.�l��P|���T�[�FG�!oٰ���*���XdMŁce�WXL�
��``FT�f����Z�%��X\Q�_�8�Y@�Dhҿ�;i�5�	����Í�w��RE}�$K�0���Ϸ��ٛ�::��>�YI%B|�=��ܶ��0��&�7S�C��Ϫ��D~Z��8�,~�,����ɡ��R�hNʽ�:Ff�s
E#1)��]NZ�fJ���f0-������Z�xr�ӧ
L^�C��qt\�s.$w���� s����,�p�m�{g>Pu��صV��eܒ����4%�q<�t���^��EU�gve�������l��-����q�YN||�5#��O�[[/�5��
����m�\3n��_Մ:
27�|�����H�6.V� ���Q��e��F�u���0`�6&����಍1I������j$R�=nq���nxt��Kv*�kjjR/t�6bvoF/}��B�x9""���/j���|���R�:@G|L�]T���V 4X���<�t��#E�OZ��}� [__��[�wS 1������Ȏ
H8�3�65���:uwPYt�����t�BtC��kb��3{$���b��W�f�s\�,���&'#�M?����h=��[r_gō��2=lܾ����ﴒΓyw�.7��x߳zs����<��O����ٹ��'�f���_k�2�z�ȓ���q_>�:}�כKm��ٍ�ο/�l+5K��� &M�A/�v�e��Z�}�B�!�~o��5�ͬ�=;���E�t	ޮ��6T�O6Bexb��8���WUt�W]�b�ϟ?��탿C3�&�!.�{r/�K7H�H6̻g�H��XTL��\�0�1�hYhX�lt՝���b0/��ab����mTӼNO$�6��;�o<lڴI�wɛ���֢>?��R�&�������g�����5݃#���~ű�zw��*憫Q�<�����U  ���M����7�GR��7䲠��5��+ ٸ���o�+V���%C~<���DhI۸b�`��4��ArG,���f?����e��A'.�uX�;�=S=�������~d�P81��60 �$��<^�a5W�<V�5wV�%���g�n����b�Թ�"��^���G%�:��vH�A��W�o�� �.4���͛��Մ"��+۶�7�jI�����s�>� ���녚�����$W�U0=��F������{��N7\�1KEo����Rv0�� 0�\��Ӫ*M%�Ƣ\Qā��y�~��'�7����B,����v.Xk����j���F+�$��4y���BM��C������hD}oT����Xxcd؜2������孅�����������d��u�'�0������w�SbEm6�#5Q�r��g$�\�$ �_��X(27��'�Ӷ�l��1)f�ak"�{� �[9Ւ(0	��&��-4���M�����8��$\�i!/�9��:8:��? -zخ����yy�����������{5�_�*Iz�4<5ԭi'�fҤ�zC� ̈́B� �s5�e��C�o�C&����?�oMp�/J��-�2�Yfә��y���u+�����ՎX4�E���k����u����q5�AېQ�ɬ���<��e�MB�x��5ˍ�L����QuJ+�����%�o�OV�r7�n�4_@hX{"+;��g.^^���{�J�宵����6��U�����o�h�;�p�%i�� |`��r���Lw�<!.Vko�ת|�l��7%���N\\�4S2����@ݠ�X�|��6 �<f�k��3�%=%l�NzOH�e̴���HMZ�M�7�d���o�k�:�y�ff��=�e[��M�M:%iL���'m����$3C!��j���ߔ�G��4/����LP*&��#[�L[�|�� �u�U�;��{	B�0U?�iQ!��o�%�v�!�I#���C��=��O1������z999d ��V#�:�>I4�s^�о#a��Gž�<�Q�jo�#�B�D���ߎC\�m�x-tE�����"�����F��l��5ݑa��9�sG�V!e���헃�
[!����'HȅN���H����&���ڮ�v���P��TI=W��ۜ����$0���2���O��O��	���Aw��Z��m��Wq��s�F����*�!
���OW)	9gut�NR)�N4�ƊŞ�DpHXX�]��B��,�Ѵ��g̢�R'�$z�]d�z��qZ7��ll��1�������6��_� �p;v������t�fټf���>� I�9� ��Zvc��NـK��m�cŤ���=B�V,��-�'����߿���F߿Q��p3z�����|�351�hDI���ېEYXXl�]�J>�
>H௩L޽Y,e�����o�����ϛ�jo� �>�^��F�m���ݖ���h1X�䇢��4���2.��yr�ѴHک�|!�V�K�EFFV��<�tjj����WΏ��UyB�m�v//��h�������{'�"?��^�fS&靘��h�u���8�X�����ޓ����P��b�E�	;�~��� ����t��
to}	B���ӏW������_e>��G���A|m?�;��al�R��OK^��#1�~A��e����4_�$�='AX`�K3�$x�b�\��#q��3��=t ��
�������$�
�&ל��;t6�x��$t�%��ˣ{�Sp�h���>���% �?(s-�ԽbJ�L��q6\
�[/���*���H���*�hs<w�T�2�ߦ���e�"�����h�֢
��Z߹������/�t#;�˙��9��!���4�c=���if��}���c=}}E!�Z� ZH��mn��!Q��[��OQU�3w>$.���2s��XrTV� ���zo$��p%Y w�@��� �:�����f��=1118�g���i�/�il�T����D�n-m �>�N9��X�B2��ja[��"L�����%�J���O��\�����D䱁'`��Ā���/�{�b��v(?A�N#=:��h�ק-����қ���~��A���r�g��2%o��ܹ}e���tw	@��$H��s):���X��N��HKKS�Xв"�Z���*��I΁YP){����c7�y�c��D�����pby�ZrM!��=��� ߈Y���+�����F��Yc������2����@��������6/^���[����0�����9]\\^ggo�k�4�	&PUU��B��\7>���H�e�O!?<`�z��P��@h8=�.�lQ_�eCI:   �>��3�?p�^��v���雒r�7�O����`}���#@��\~~�S;#��橲���=(�!��8��
�%�w���{���S���$�w���;��;� @��O �u���ޮ��E���%� ������w]�zn���$'��#�h�]�Ҕڜ~�w�~�.@R<9���#P�Ԡj 4�yidd�U����Ք��j`��>A��[��AF�#j�!��C8L���*p%栍�a����w]�	� $F7�E����<�����Z(�`�U�fA��I�cp	���g;`�ɗ9r�|D�_/]�͜���H��RQGJDM:p/7�E�L���ӎ�v���Q�Ǖ(#��_�^F��|4V���C��y~�GHL���������;��]�=:���� �ֲ`�J�t�و�q��iH�M͏0f��"�7��E@�i�����aB(ף[��F�ggg�NIiSw�H~D�@��#w���'~3KE�p���X��#*@TK!%�5���!�T^F_f@��@&������,�ѯś�?�#D
�Ի
�84n6�#�IW���yHYzTy�+��
�Κ 2ˀg�JJ����D��u���@���r��\cJ��=߅�|SLR6�K�::���k�M�2�3��m��Ex��,u>H��@����@ ����T+��E�(f��t�������@�0׀oxX]�[-�V}���
K�6 ��+Qso�����E�Y���������fS�����U
i D�p��I~l.P�>�:V��\����t�[G�#��lZ�.̈́8�>����F�H7�8�$%M� ^������q�v�q��֓t�*I��*�<#@֐������n�K���Hˍ^�O�k ��W�R�fl�X&:��'������ad�]Uѯ32��_P�L6�ŷ�VVň����V�֜P,�eKǥQ��P�
ڛ��kH�sD I)\ʗ�L� ���n���S��߹[��n ��y|p22Ǘ�ߺit�u�7%K&:��\E�[vVn��R� ^ �|��ƿ���C��==�WzE�W!넄�>��1�V:���p��U:e
��O�i$ҿ���Ħ�êw��}�l-T���1�5f�K
�N1��zR�u��$==-]��d@=2�XI�!<<�f�./C��!���q�\�&�i�l6�������5��7�t��������_U�������\� $�E�<�]���"�<������t�廬d!�B��Uϡ��=(_Ƀ��^�'B�)��ucTkƯ�zݿ�.Giv0�Y	�--��`��F<�u`@Ŏ��p�F��^��BAY/L�y5J�|��-�x@���۵(�itH�c��Y+DPd�`F��Q�����q$�ҽ�%�c�h�&77���l$�)3�@��<���mX�=�	��sXpɐ�(��q�&����ۣbmpl��Dt�LdY�4Ru������:��)H���B���$���S 3��_(��Ӄ@/���$�ƅ�}�������MdQ2uuu�zrss��W>UA��V��'��s��ZL��_�ta�#�𽍖"����� ӏ���;{���Т_Z�z����L�i��������z�p�D{�ʻ�A��*Fx�/i[:i@��PՋX@�ԺLaj�f�A���ڌM��5� y����kz��~1vv�҈�f�R9����Li���+}j{�zbں5d�U��U~� P*d��VB���<$S��sj�|���r?@3���^����Ѹ��*:�����oL�h4��Ż�v����s\[O�U�"�u/��mP����/?�[(�$Z�����mT}�&�`%�T��e%��k0��Ç/XX����./�<$��$�M�':�P�zMl.m�M�F�В]˦PP*�
!�|/6cK����9Y��Z���'�6�'
�H�Kx6�~�ƿ>B5V�
�,�S��N\��zz��b��S�NA��������m��R,dK��h݉�D����3�\'�*�̱�q�y�[�Ys1�Q�A�(��8�C�jM۶��`oOK�t�re���c�]=��/�ӈ��6����c���9[jB����������Q��Zooo��,� ���'���(�Y�N�\1�Q�>�}�a�aE����C�Pa`1����X�r@5����Pg����m�C�9|Q4
���NCCw��!p��O�|뺶��MuU����V��]s�E�B�օPf�����WiƝ*�p�9�P�c����Pۻw/���Θ�������:G'*�iR��' �_�H ��L=�y��ә~
���z�ȏG�c�˰���2Ʉ�X�����󮀇 Ę��y��5��=$$� �����d-5QT�t;d���64����/��W@EĬ�e�M�6�'��9D�� �4Z�ԛ>�Ґ��ⶒW� �9��}����T@O�}R�����҅[����PG�S�w5��:��
��@��yANW�(��sp2����_��Z�	���4��
Ҏ�԰���;��37o��տ|�r�$��iG�n>0�}/@��$q�3	����Y�b~��Ŵ@��.���s���(��z��2��(��םṞ즡O�t/;�z���ʌ��}��95ONN����%�g�i��xH���$��t�4�����F_w����+��ď�y���OG&u����{�v��#[lA�`��QH�NÝ*��a�vV%Kq�Y��i�S��Y0�����pat *�rDq�66*l!�?�so�
�E&*x��;��èbho33=�?M��VA��ϠSȼy�" N��::��$5�Ԏ�L��hAC!aax��������
-�))�z��������VQ' 2���3�)�.���n��}Tcע/�@U���)��"�>h��0��w�m��l��}l��'�X��U����DQ@׀�燺��~f�� ͷA|E��u^�Իz�\�A9�@{ie!���^�9g!�F��-���N��V���m�����Pe�/נ?�EݧŪ $�
�h��o��Ѧ	�}[[�6-GA1e�Ж�7`����%�y�oDA4�J�܏J~��֡r�w��`�eAw�n�U��c�aO7��<H3Rh+
���$:�y�R? &HۈŹ�[���%��o��������C��h�җ��1��#	&z��h=L$-=�D���h&���Uu���9�!��բ
| |BϢ����������	�DM$C��qdn �3�M������+ShfP9i(J�l)������:����V�� ����𑲵��E2��xI���"�%�=��=��
��h��F��NII� ?��R~d�ٷ��[�r�Κ-��o[A���wݻ6l|���F�'1 �C5Z�S�6���NJ(Ix���px��+�6 %��_�~@�D��\"*���p�P�#�DA�~��̙3q����� �$�����Bݺ��V���`K ��� v� 7!�@?��}��IE���9#}�w��&d��Dx���@�/�w�}Z}�s�4l��!g�d���
=�C����γ�o�:m=�w>��}���`] \Q�z�"�� �@��
)�x�PA��-.ix�[�e�7�vȂ��s�� �����f���W���D����^DU[2-Oח��P�N�u���ٰ53�Dr���9h��6�_oq�ҽ
�/��;��Яs!G0x���iՒ�o������8��Z`��|XG`�[��+���Y�*v�*Fw�
,���m+����vvB����y�o~��l���$Rds!���
zO[-��W���&%GC" �!W���0Lu�F@��UY@��G��s����RT݃� �A� `A+ kNHN����`5��C`F[:���蘪	���`zE}�2y�������ޤ�K��������ab�A�Z�]ꍾ:ea��;-+k�4
|�m]�ȥ/R\�jq�2d����U�o�
�,T�� �DD�w��Ǡ0)�l�i�s��R	aL��i �/GNf��Y���hi���M~ŕ�U]�#��s�=����^[����P})PG|||���е�%���4A���谿���A/L��ҧ{n��� [��V���V2�oiu`c�@�[�%L�DFtA��\ 3h��H����}�>���~������6�mk�~�<�=�P��}���y���>�6���V�E��[�[9^ۥ|�l��X�~��haa!:������`���v5�b���`�ԃ� �4_-4�2���YX��W�Ջ����b@�M��!��T0`h*�c����㗟�[O��� ��7\���y;1O���X��TU}CCïz��e7?"ɒ�6(	`A��]�/}�xA���p����t5�p�r�>{l2�EŅ���̒t��/��M�h5��m���[����
w��/<��%,��7ȩ��&���=�F�y��������!ˬ½rBd_؇{Va�u܅&�5���fw��3kW"+�|L�:Eu$�Θ�>�3?�Q�Og))Qѱ�~��������͔���O�d����*������M{W�reZX �Μ�9τ����#�y3��M�,�#ˬɜlҦա%����S�h5,�:K���%�����深s�2�3|�h�V����c�(X}����%[Q zG4|M:sz(�;#7���A�8�h�8�]��K���,)�%CP;�1_��F\�8�^�uN�i`U�����!�Jg�:�Ƒ,C$��c$��^Dr5F�
H�. �Ia ��Eǥu0L\g�5��L��%xg���Z�L�4\����wFNM7�z6����K �
��;ܕ w
8��Owb�]
������0�>l���3�[��F���̓r=p�r��I�Ϛe��^��;�L���⦻���`��܋{R=	5p�r?� �I`�6��|�@=xX�ql�z�l��5�����Hr�Sn��-f��'�?�`�Ӡ�r�jue��?���A�Mw����,YƦ������VC�m0�P��П��p���:xă��<�'��I-�V�E��`����$�Q5B̳��k�����5)\P@�z�Y(���@�M'(�{�a̐��&�P#;��@O5��5�.V�F��Ƚ;-Y2��!l�<o�� ���&``���P��}Lj�,6�G7��;��)�}����ܛ�]?�3� ~�0�S��A��NO2�f� ^�d	�Q��1��la܂��:5�Ђ�p�B�Q����Hg;X�#(�I�,�U^"�ryբE_ާ�~yY~������	a�ˍ�'D��ě���n�7���^��bG�����%�7�~1�f�}�x����{��4/�bhc�'�lw�x�����<6݉��>�0�U��Ln#�}м [�aඃ�+>b�k6�d�~�m��}��,X����]�E���Q�o�Q���|�:v�(�K=�gZS��x��Jg.���0�\.���a��;��<Rs�9�`s�	�+�0F�B�� ږ>��C�%����дݡ����]�G��ׁ���8���@��9�3q���v)�tȶ���������J		=0OP�X+ a��9}�h����A�L��=A���ى�<�Q챫e�d�Ŏ8�_Q�I�Q.VL���jN_�7�=��+0�1�1��0#r �y`%6;s���6�[���+�n(ja%�b���0� ��-Xo?PhK��3��XC��8���P."�c*��jw �|�qr0=g��<��D���9Z^�q�8�1�uI�  ɂ� M{� .��b\�(�ԖJl6���<L{=�E�� �3B̯8����A[ڠ���V�A�F�Pg���A�0�!Ѝ��y��`�o�F����EY@:�X<�A*���C��zй�GN�1ȡ��=��������64��M�]n�`����uє7�O���d0�1x<z�P�I!xyV��z��<+-���j��G���!~@n+�ۍ�J��7���6z� <&�=�=���[�<�#��t.m*hT\[�=�6Nw���2kAL(�H�2��[��f�"��K�{Xg��,��)�A+`�3�rK.�� 3L���<��1���$�G�5�&*����a�%
3ʑ0иBἇ�\�t�� ���'���=��@�w�F1�-��߽��y9D���}�fl�ϐ���V��F&�̂�l�R.�}������Л#O�4�ڽ��]柈��-ւ��h�y��	���롣7p��!x,�ėNK;���z���Ή�)����߀��7���o����d�|��,������o�����?Tyß�m�$��q�M7�����W�v�(���(��%�mp���Zv%����.����)��<����1�R�25.����w���x�,�[������w$�R��@X%�����~�O^��v�����*���_ծ�1���#��9���F���,�o��l,Y�x���nof�Ϳ��:���������՛y����d!p�la��"�LK�:�I��v�\SS3���o:{��#:�rqq�`�s��U��\����w�ȴ�`k��+&ѻd��;��`N���І���C��&�ᶌE�mĕ�\W^�m̑'z�Z,�;z����&����f�u�3�8^��4�V�naU7����Q�*e@�1�
/PAGq)�-�w;,Y΁D�p��Jg�]���HB�}��gqcK�NgN��2|;<��eǵi��8g���4���ma�mÿ�o����2$.'����G�a
�Іی?z�ؠ���NÌq��|u��_7 ����m�9���^���#�����q���pM�ΞH����t��vVc�@�hÝ"��m��w:��NK�Nk����V#MK�[�vǷ�:��9������fh�yP~��ݲ�8ۑ%|]�Sja�q��Ƴ������#}a�7�3��mE�V�ZZ$U⒣��n罠��Pb���P �X/���FÃ!G�}�AA�����xP�]�{0�A��G�8	�S�Ծݚ%w< ����H<��=��u�ʊ����ߒ%ȟ�ݲ7�r9��P9T��n��Oa�5�!�ȴ�
.��~\Hp+L�6�nq�G��6�U�� �5@�G#XA&��0"����x���&���cp,���~���ha��Ex� �p���J�����v`j>�
��aj��=(^D�8FG5A��q<m7�m� ���Q$��ë��r���fl�0ƅ ����	�@n�	�����6�{���XW��~8�͒e	Lc�6�9���K���/��w��1�P"���k`���Jc�KnN��cx:� � ��Q__o����]ϴ`��v���?Y�$���q`�3fc-���i`w <�a
{ (�<�Jm���A��_ ,���n�%�e�EϘ��Ā�� �g츶�І�ۂk�!.߇��6D����6"zH�*�6D�w��:=����:��6f�m��D�������w������^_?�Ӕ��ǂ�ҟ0+7箯��y��E��������(�F�1�^� 2; 2��d���5�hǨ��D,�n��q�ȭ���]n����[,YZ$G4a�J"��Vk�� 1�� (�bFM�F�:�?`Ѓ��..lv���`dn�Hel����Գs0�	J=y�/=��a=n�`(�l#N���"�K�vূ�ԭ��у�@����"賥����v=�6(�C����{9@�W��a<A�@�ژ>3�e��(k�G��|sB�������2�B��`S� (9C1�W��NDp5Fp��>�wb���gG]]]C`>�!�%���b�3�][oς�bzр��J�`��w�L����T�
q��U^�D���Qah+��]�U��GU��]L2@O���6;�:���M~�; ��,Y�f����<"��Wɵ�}455���ߴn�q�EG��)�X6fa������bbډ(?��e��چ��xR���� z)y�$P`���*������	j�A��Sy9 ��0����R�|����� �P����c��)*6"h`��I��bn5����*�
� #ڸŚ�q��gv���-���P�ȳX�j|�k[�� s=;���$�`y&�z:,f+���0��5g��C뮑n�����c����%����|J��Rn�W��S�qmm�Xk]��̞fB�ۉ�����؟����F���c8}���|�Q��׌'�e�u���E�r���i�K<�$�Ý"�l���g:��%䌗|��Sd���c���D7C"����_$t�2��z�J�?}dE>�������Є�O2�����2���_���+�ꔈu���?+<
V���4�㿎��u��(ϑ�2��&�F��n5ޚ(�}}�ʢ��ݷ���V���\�S�^�����	��U]e՛(&f�O�}~v�Nv�Ԕ�?v�:^`m��v;d�jSM��#K���G'&���KM�.}�Y�<6�wf=�;@��j3o��?�N2��W�B��蠣�YV����c���7�A������p72�ѡΧU�5P5�ᨤ�&Y�ώ�d�mQg'5��Cՠ�i$��rO��믧����u�	h�E�'��1t�4�fK�R�k�{�>��A{���n�߄PR��$���I�T�W_=/�g�q`�{w�E>�LmB�"Rܙ�?��dN��q�ĭ#S[&������yǑ���\{��ә�C1��_�Y��/̮��aN=���d���=,&�!�a��"$�
�VX�ߜ"ߟҠ�����0q��lE�������h���T
��B�"�������B��_83h�DPVN�?�<�I�[��ş���*9C��Tiq�*T�|�����R�
U�lg`x�ƈX���t�r����x���wP�T�7v��A�aC�c#"����j�_�:TX&��hμs�g�Sf��w@�X#Z�/��ԟ��Z�P�i�y*E�"��k���4L5B���Kz�%�uӷw�7��v�t�,s9��WLE�7)ͺyvq����J�.?=���oi�xs���_?prk��k|��G}��a�
/+�C�ŚV��IDC��wޢk�2��ag�{��?Q1ȑ�����ԩ���mV�Hځ����>:S���'JL���3p�}P�O�?��zvh��l��=��V�Q-([G�a�\�^-ꬦ���u\i�@���-q*�z�2�T�Z����n@S�M�ۂg3��-)uFa�I؍Q��#���@3�pJ՞ZjW�����d�ԭ,���(��4�"�.�(ƻG�Ѷ%��c���,�!�!�9u&k�d�S�'�*�2�R��s/���zn"����Zo�|�d�5;4f���"���db�fMigف��$ܧ���k�f��>�x�?-)����I�y)b�N^���ՠb�㿨��ء��rxF��}*P\�雓�*�^v
��k9CU�.ػ�.�k���1pC�\x��v�eӡ�R��88#$)G(,q�Z$�����z�V�7L(��.���6���&n4�n]3���'�숓9�5rr�oRs(v������X��@���8ůT�%��o&>�S�0��R;�z�!�1�t���ܤ�
U\�a�m'��IԎ8Ǘ�����bQ��L&:��L�RT��_��F^�"n��ݺ��{a����xn�Ȝ�_���V%�N���U(�Dq�հJ������B�k��$��fe$��3x�����cмǌD��m4��Rg��UrS洄s��W�x���]V�$�H��տ�,Խ��&;�j�L¤���J������I�(���g�m�#F�|*�)�)��"��t���T��x�֦u�J�12��<�A�]��<�ϣ`�ie�'��W!�Lt~X���r���[TZ�ckB�ǉ��q�8#��Ó��s��?Qct䘼���JgS4F�8��w��eD��ΉC?�[iB�[tU�M�&>��^�넦Nn�w�7ڀ�o.�k��{{L��I���Pqd*ى�E�HjV��	�7����K,���E�k	�yo�L�mr/�-���Z_�jo�1Ev4�}�3fI���o����s�د��l�zpb7HW��E���eP�+r��z�)Vገ,�/6W�-)�������ɚ��Yo�?��4����(d@o��|�J@,{uo�h)�9�2@Q����ws�M�L�f�(�i3Pg�ӵ?ko��8�5bQȋ���Ϧҕ�Yv�r��HRS���ki�(���g�a  }��Ώ'Y�ޟ�|�ڞ?Ш{��M��X�$����K�����JN,O0P�yK<fok���lG�w���IW7��LH2[�Br�>���0Է?���SY�9�Q�r�VO�,����Z����씬����Ĕ���觢��r�r<�<.>:��T?��\Ú��H�g��2�zL\�yp}_1s�����Dt�K��3 	!5Z<��x���ZO���&��;���ニ:�}+u����1�T�<���/)+f�!"ݯrЎ�>�^��!2+͓�w&N:~DQ��T��)C��k��ҝr��UU�	��`B�wF�C�7yh�H�;�F�+�)�(�q�u�^�Xj��=�휾�L�0�����=����j���I>�xd4�,�)�lL|1����e�^��ߓ(u�����t��?��o�u���4��` ��3�&��b':x���'n
)^J쬾�('+#�]#�iYߦ�\��2:�� B�iTc���Zs��
/E���lg10��})u�a`D�Z�L!�E�J�O�� ���P����J��r�0���%ny�a8]�r���������0L�.+}\��?�c`�a%f��C�F.u�^� G����1Rg��r0v5ҍ	8�D|J��.�� �e`@:S��O�_�`@���������J�q��h�d�.�t�F߁=��=#:���Ga�?Ƶ�s���e��M�bYL����0!�<�R����d ��5�����\�\]�0��)�i��:ԟ�V�Iz���x�*��j���l��	�b`#=:V����g=��j�b��Q���<�~|��{��7�mUթv~ף�2�Ա�r������dz����NM�d@u�����b�Pg���ݓ\nka̾R8ձ(C��<���{��fٷK��� %����bf����K]�t�����qR�S�t2�g ��n�?��w�T�&yA��'m���F�~.��?�Ni�I���K��u�{oˀ��5iyq3:S?fy*f Q�3��U�u��������P�;��ș��Q�nC�72�zs������ݮ�e7��? ��>`W�-i\��:����6���!�7�m�����M��%���5�����c���Z�z��Aׯ��0&W��{���mP�7��]Kŗ�r2 ��rq�q���ͺn6O�̿i���#���l"#�?�g]x�e?���j!���z�VMjV���}#ī�|�^���K*��dEi���_�>8��4��:��`|w���	�K;V怳����(�W1��Qj���´��L�x���G��1"U�7��:�WԽ���ok��NPn&Z&5k4�;&��F�,܆����ɖ�3����rnvS5"Z�A�{�S^�m8�"Gef���.֐NsW2�f���?O\��;�_�`����
��4���F�)�,j�T��ԯ�}�3��a���Ru]���:N}�,�J�0\R�O��8w����1VZZZ.lN5gS��9���Z�=5<�;����;�đ�߇����E����Fø�/������d������s�����[�7���
�%zm��9�F�nJJ���I��T�ʹ�H��{`v��ѽ�\�NB�%�)�rr>2\}(�ִj�&��r5z�յ*��n��E`�O�Z��5N����@���~��ި���D)�)��oY7�j��rF������]��l�xy~�&Y�u�۝�3[�.A�ya��z��B����;[��X5�,�LS5����%5v�j�j�7�[�S�Sv�~ qb���늶�0�=������-w?�}N�p�	��M���2#�w�{��Ӝ݇�� �vt��Q��u��6jd���.��5i��R�6=�
���WIA��K9�YVBd�[�G)�#�(�{9W�UdI��fxh����'�U@b'C(u�R�r��S��,»7x��ʐ'~9:�fg��;����y$����:�oW(�(���yv9���Җ�Gmn/����6jZfZ�����	`�^r�F���̰#�U��v>v����L��Tg��a�MJ��+����I�f!⪄������i�I��bW�7k�c`I�E�C+�<�8�N���c�0^�p$��Ҭ:Ĭa:K��+�O�*3��u�Tza�d�3���)���AS�ī���?�t;Įo��e ;����k���mrl7����AkS���9�_��=71�$�Zu��ඳxBgH�a�)�u��R5�v���U=��[�f�FzY�s39��D|�:�\������X�º�:����q3J��x
�c0WY[{{Zyf���@�.^�¾Q/�O~�JcnW�Y��V�}O火K-�g)���,פ|Y�m�h�s�.�I?��Ԟa����"�2���s��F��w/.)�I��[��C�����B����Yi�m�@0W4�جW�A&�jC���Z�4�v��Û�1�<�D�ב_܆�Lx��*���5q���q���W#8���>_��ܾ�f,�]��G�c<Xte�i���:���5��%o2�X3�%��i*N\�-�%	Qk��;��z%o⽞ +QwD��OΏ'���#��Cuݜ�,�ň��*�JM��iۤ2;nQ��ab'�����x��db��#�������0/I�y��j�X%��q ��˰����K=8����`ͱ�׶�Ę��O����)��P��R��{�N�4�� ۵�ô���i��
�FŞ���"+�<��ˠ�o�o�T;s�N��63L�����J�먓����������"ý ��#o��j2���|L�C��`oo_�' zb�|·���
eѠ(f��n*ԡL�g��e�~2�U|b粰ӗ�9�2���/۫���8'yʱ1��\�꥕��v-ɻC���3_�EY)f�e����=����=����/h���+�Z��b��V�S7���K�gE@�!�"R@A�a	�X�֕Z[AP�%3!��HXԊ�7������|g��=��˽7s��O:j@!WN ��rDb�c�����Ȧ�0G��FI�ٮ��뮁\XBWxu.�L��,ۄm�߅�X�y3��W����_i�׻��ٸ��Y��v+�i;k��gd$O}T%�Ti;�7���]0Wft�O��w�J�5�����ѿUv���S&�nI"ҽӼx;�\����?ȱ�5k�d���C69��cUz���)l��&�f˜���ܥ^غ�*�N[����F�3��v�O�a�V9n�y��y����)����'�ކ�o���](C���m��{Yk{�禗w=ݕ8��n.����-{y����լ�Q��Ӕ����9G�\ࡴR)��G:�t|����e�&D�|�ѝ�;�Q�����.��
�5�YmVP��#�aa��d�֩Y��OSo�5d;�;V)5�cteI�n%���K���낌��C6��{AD;��$#c�_�ƒ~54��m��D���F��Z{��`�*��ȥjiGlXM�*�U����b{�"��	��fs��%������������k�g�+f���K���/���^�j�ϩE����K��s!>�/�/�j݉���k��8^��z�,���]WIxs�:B�q���dt�ő��Oޥ����'�����uȚ7��"��7|�KA�B2Ȗ78Gܲq{�$1C�Į~��8���v�B�u$=�I�<Ų�Q�w�,���gB�6��d�w#��_���re��<H����Ir(Rv+�Nw]}�x
9K�8�N��kJ��e�X}�F�r���*��D�֥x�؇Dڞ*A��s[[��9b�ӹax�б]�B�6-�ZR(3�a%��Ʃ���*{���j���6<��sE�A#���Un7_�k�6�U،����M��y?���|7�WP/�%��j��YD�9�=e�*�ڛ��;�mT�R��&y��F!��\���=O�(��>��q� G1A����Lk�������ӻ�kB���GtVd�_ݖj�B<��IcӇ�<yED�|º���TU���: {0�+�Я*OJ=x�DS��q����,x�m1:���K�<��@�3�x��6m�
9�.M�:7%y��[��-|�z��F���wW�e���%��C�k�ۻ�a���Gy��5�?8�hp)�3W��	��˜�k$��y{�|l9?��=�5�E�!��-ݎ��̎j}��@?���6ͪ]�����y�b2��!x��+/�$E�O�2�z2|Gz���r����{`���<��_1z�nq�/�ڎ�zU��}��������$[�/���������ks��Y�l���L������Ym���ԛĎ��o/�\hd�in��l9������G!b�#����&oN+(�إ#� ���\G���S������)���&�X��6S�LO!�X]�\I�����Ǥ�fo����eP���Й׏��рt>K����r6��t�ذYr?v���NӘ�@�<!�
5�'��+���p�N��^/��C���䌽<��R4� ���/ׁ��Q_�fɪ;y�分V��'�0,�����cǸi�Z�e�q�R]-2m�:�V �7O^ƍ�������<�\��=�K'��6[�_����������L�`t����f0�C��R�j�d��&E��c�o�D./��"=�hl�J��}U��(}��q�X8�xOc���!ٞ�>!M�J�h�N�(0G(�,$�񡬐�J�Z׍C�z|�Lѓ1�� �AY(�I�H�u�,q֥���B�X���m�bR/6�a��hm�k?��C��k�e��������^�7<t[?��uHorU��G�2�(s3D �3�rnpb�q:8ٖ��~wl}����5�c�
�����@�"KQ��P%�/O~��$Q/�w��<�y��tvǂ�=P�1��7Rk����z��Ɍ�"���C�ߙ����c�L5����=��O�*��̸oxH)/�
E���q��<�;���A^wQ^V0g��R&��@s(:{20G�xj��o�����=��yn��"��jO�a-X}12Y��L�K�����	1���c�j0#<Ʀ�LD�Į&�_*Ě;�zll������=%��iMf�a����w�s�6q�.�\��ԟ'���efG�H_�H�㖢x;�ĵlJ����J녲QG���i�4o�y���5Vg���O!_�Q�3V��T{fx� ?�ß���5�P��o�E��U)����-w W1��J�ŲQs˗9�uTU&u��<�(��z�`���7l��O���d��Z�xb*۴�{�{�)\��)�'[;���:�aB�Ui>�t��;�m��T�Ho�@g����)��$�x��ґ�e�u�=�&�����s�';r��y�AD'`�<d���EJB�;f=�H(��b�����K�$�"��D����vN/��XY����׋��8��C�f�˽%�#'�5lҨ'�m<���l�o2.�`e)SX/��R|͏���x�;�"Tẋ���0�N���֭���:��zFq ��]G���������w�Z�Ok|��W���an71������o�{Ug��
�}9"���!%��c��y��MᎵ���}�<�̍��(�sk�/�iAyv�Z�u��G*I�d�	��r�8W�.Pg�6`s�'�����:E�k�-"�r�[ ���s�����X9�S�����8�=��@:]�'�ZI(.�Pj����~����GDѮ��䑢A�h��4������z���F_�~��g�dsE�0G0x^�s)\�4����E��ѝ�����Uy�<Kv���y�D̋x;�!7[�^P�#���	k�4�d}��[݋�0�W޴��v��l}�\y�!�zA��x2�6��ƺ��%v�Q:[�=~� ���j�����T��y��5��~S�X�#t�����Vm�����K�&����������j7hp�+n��g�<�@�&���C�o	"�a���9Q�*�&+��,��8)��~`_k_m�Ȱ�΢�S��+�J���3� 2��J�m���h�}K�b]�Se`#�����Y˵��[�y�����?I
�`x�d��SQ3N�F�A��|S����ى����m�Zz�'<���BT��9ۿ�kc��;�*K�F�H,6!���/���9("��21������
o��E�~�f[1i�En�����aCD�!A��B�P�(�QTooRD��lT�^�}�
�|y{t�)�^E��8ޗ�f�#3LsĎD�Q�ݎl=u�1�l�ma��0MvY�$2�h]�O��a���Ǻ;�W�#��/�P�%{�����f��D�o��t_ $E�ě��"�$�o�W����Z#wҬ� i[ɞ�[�C�F�bu!C�/� "/FV_�)���P�9���y�l#�6�B��]g�p)����C�Z�\I[*�Eb=��}�6G��D�#ߚe���w5>��"2]��;��8��n$mɍ�ȩ]��Y���`���Yj�k� �ʔ�m�-E��Z�E0�ғ"�=[�?t��NA������a��U鈺�l�t_��k%�X@4A������Q �B����y�֓�Eg�U��go�e�}��-�����`��t��(s6ID�PF�ې�<�E�Q% %oDJ�C�_��j��Wp_��@��4y!�I<�/�<�k�-8�ҟH�m��Qfs�^�lYD��7L��@��]���rY%p����M$���1�m�P���T�^FX/�2�E��K�*ԗ����G|��v���Ԋu΢6�R��D��v(���G��R��FR0�9�%f]��5�.���靹���e��C���O��
z�㤠l�x��Z�Q�Ke�AE
W᎑��+.#-r}�Ґs�{n��g�~��ђ���%㇯����ﹿ�\}h�w"�J��Պw�SG��������Ӹv/��j�<\��k�!1�='t�����2ǻx�<<���?��p�O�E���t�(��M��?�&��Y�MG��&ǎڎ�!&	������G��È�-+-�o��.�o��ָ�YYI�]�Y7R��MN�:�_�1�tD���I��<��l���7��z�U���r�i�#j�l�buQ��*a� lo�5r�iQ���:�`��*��2�ʾ{�f�_�M	�݉}�LZ9-�m_���F��W����#��r��~{�N?�5�>8H7�7W}N�u�ٲ����N��ŁX�j��E�����+���c�:���� ��w����<_X%�����/��X�������= �v����z�,�� ���-��EB�����b;�D<R�Q"����]���x�҆�MT8&dT����&w���J�����D� �pn����%
��1@GR޼\����hG.���V`o�8n7� 
��7@NK&�ũ�3C�;����A�]��\ތ��k#�6��p�C��)=�)���
;ĳ��@�b�b�J��]��x��w�t��O�#�b���h�*܃��0�a��M9���,��?���Oq��zѦh��zn6،W��G�D;u�'�X�v���唂zD>��?!��m<��ؾ�m�~�Gj�[��W�R_�<���$b��s �NdJm�s�����e�"�ђ�D�U����[�Y� 6d+��a?� 
9O)=���&�U˚�lݎ�uHhd�?���"��Ȓ��9~*�=�8�͑�&�����H	�ž�B�V�]��S���s�Q�[����2^�٣]�k�19}r�����:r(e�^�W3@��Yӌ�L��Gz���T7P���5x���[,�`U%��*�As�u.[�v�z�˗-��:�Z}*�$cq�i��o{����SK���T}�I�ۦ��C�T޸1�� D�l�U���n��*&�������S�ۢ*����7������h��W�����)���HJ��i�5
}pT-���e3ƶ��I6���kp��
�[���؍���JuTY�O���	�[�>^�n�@sZ�����?O9�$�]/cZ;b�<]h�l��!d4@��{�����2~چy��8�����nha��YI_�c���Rh)�|r��ܐ����#���R���$�G���`W�v�y��eH,��ڲe�u遃H���6�'�0���5�J��!�8C�.��
��lC�9�0�	�}-��d#�Eٚ
:�x��(�~���S�ҌH�^q��Ą���p��c�����@��*֢�_GM�6���K���W"M�B	_I�İ��
u����*4��
v���PPXg�H�L�j/#g�s�Z���wD��|}1�AK,F+�#�JjĢq�m��
�������m�OG �\��,��RЃ^
NƟfD�Wz��^x�z!�U��;���r~�=����t�qҎ\�������U���+m��v)RZ��f��@��_��L�.�[G�aǅ��8�E��xV�"�V��U�$�"ϼv���p��!�_�q��x'#��E����\f'�_y�Opp�v!Z�GF����\T��[��v��O�v,�M]��zq��7��]�S���x�o2��i5���~�]�v�,�q��=�\@���x��<_���N�A�����R����p߶Szj��U��]�\ND߻�O��˟�W$45�.\��]���~�Tg��$6��,'�G�I�r��L�c�ωA�9�:G�C� ���3M,�0ݩ5H�ޤ��U�w��uE��|��vz��P�<�o�c���Tl)�Q~�l���ކ{�K�P�A������̃G�v��U���Ux�i#�el�Y��RQ$�%n��x�3�<����Uu�Y���+\\��R�/�Q���@�K�{��zZA�o�ޮ��f��2 7�`T��U��0\;��
-$���TH���]0���4#��B���?� &Ըq��]Y� b�Ĉ=X@����{�
3�u��4<�5�d���U5��`O�F�,<,�kTCS2*�Yf��b{0&��M�^'��.�@dg�WŽ����I��u��3V���۪j���N%F6���iʟW&Y��#��ۛ���ɼ�G�%�$Fv/@��lG"����K�#�B�ݗX��&�n�\DT���|�^(���yQ�3��V3���PQu!x�?���f3�A�z�w�&Uڒf�aѣ�.�V����ƕ��r�{I�qj,��~(B���0�Ryܦ4!Ʃy=G"YUH�[uƉAo���*ũ�I<�T�_�rـ�[���]=�V��V�����#�Wo���ǽz,�+=y�]uI���4Y��ǹ��o�'�-�kqA�$S�s�u7���D��O�X�c�B���ϭs�ղ)M��~���QBl�OꟌE�fC���,�VzcF�^� T"��v 9G]�6�}@�gVD5��U�.�9}Ű�F�
Ծh.�;��r���u�8m(����z��Ge�|���\d�D��r�	gۣ6��Q�b���H�����"+k~_"�l��Ȗ�әTH�(�c]�������0���[�g�x`�k��)8\5��C�t��*����ߍZ���\T�N�#L��I�o"w 5��>�D��|mr�K�S�������-h"���(�>�i>�d1�!���]6r�+�
���c��l�J���t�B���OX%�!$k��s�?���=]v^��a�ݔ36���.tw� �DH�Q ��U����C uM1x&��
r�M�\K�yj��u�N�ٺ�*�HU�L����r�8Q���\���b�3�?�v]���2�^���Ħ֮�ф���I����ee��벳K�dP��B/�!?]��&o򅎒i1��!�":��-QfH�b�֘Dċ5��f�����ش���^�����k�"��3��T�d�����~��(�Niag��� ��V6F쪮<
o��ȡyaO��XD؀?�FfDv��SB}��nL��#���D�q>����Bn�l5e�¡�D�c�҈�0�Er� %�������+}���fL�[*ۦ�};�:1�EB{�#j�&��ʑv�w���g���x�׋rĭ6��]� ��uNG.Æ*}7A�����s��}�LX���$�£ŋ���}B+y�.-d��T~��F��:�e`;�mV-�a©�F�J$�[����uK����m'D�ݧ{�a̭ƥQ՛s�N;B�3��j����2>���1 �Ͻtq�|�X|w�㟛�xr�TY�������|%��P lC��.3)$����^��Nb~�<�=*id�i�nd��UeKx>ԹI�t�"ד�rh���M�Z�]U�����U0�p�/[U�a��~�*S�G��.A��.���K$�X�|gD����k�R�)�&O[|q�w�kb1�in�r<L&���8E��G4�VkJ�&�^c�����m#�2M�Ew
C�*��+ݕ\����D��]K榋$^-5M�1�=��#���a1Dҍo^�cX�-�Co�!j�s���规��Gx���lI����)k/S��� W��{�E�*��h��~Dlo:��(�"M��h�������
m�`�I��RE�b�UuP�o����0�i(6��#'��5d�I݀�s?��W{U� ,�VU�|@�*����+�]����S�,����r��\ :GŐ�x\�^C�$c��j����W*�6i4\��{�����|M~v�*�G6"�K��cYˤ�ċI~��k���rrE��)��i��|�ZB֘:#�"�H�zMӐd�=7]`�P��K���D3��SV���7�&��S6s�Z�KG��h+���|�w�����f)_�s������I�����&����<2����׺z����؁H�qC80;����rF��L(�݌�6��r�e��^�z>���w�J��9���
:��p���dFBt,d�1��1#��,��i�g��md=��n�.G�7�{*��_~n��ly��c�A�&��z�/z�q�ŉ���9C#��g8\�5m?^�Iq0JC:P�@�mg=�Ƞz�Y/�3(C���A���+S"Y(�%d,XT� ��@���m���@y�E�F@iTz-f��`P�l*�r,( ]`=���
f���[Y���_�px���۾��Ȗ���t�	�Y7�%p���_t|>ޡ�!q@b[ k6�E�i��}��X@�5yhdBgȊ��:�tt�����]��`lN���/�
$�@M��d���=���KGZ�[�tX*���~�ʑ2S멜��O"bA?1F��N0H�������L(�H`�,�L'�Y>�H�r��:z)��� ��9R�eS �2Ћ�P�N`�^�7�Z �Ӟ�`��Џ28��~�o����xM IsA�
���z@e�ס�^�@���FA�^���6J��X�!%���]����r[��7�!!$ƜaL6~n����4۱4�����.�jP�{u�w+L\���E�Xyy��Ɵ���WCUg�{%��Zx-�J+��ZBs�O8��.�i�����?�eLǧ%'�^��bT���1�y��mF�4���]pu���FX,�~d`[X��`�F�f�ʂ1�,�Øq��.�>�X�V�_�Lj��}irh��!��>9Q�S{D��1=&%)�,S:5�q�ʑ�	{�>��n�6 �,f�- +e�΂l��lBg���j�ME��/�ě� �8���H�T ��R0#)���p�Mt�Ft�7��m�IFtp�2�����8�-�����T|A��4ͽg|�e�:�B-�4����t<0��H��?���':V|kdv�?���J�t�q��`7c�:;듟���� �ۓF�s��a�ǣ�FR)���-�n��h22�ĸ��P�s�m;M������ �m|�E0'_u���;��\T<Lw�������`�DEL(��f^�c\m���+� ��Oǀ�Mz�Vu,C@�;O�p��M ���`r���
~+�$�-��Z:�Rn�k0��3:eB8P8w�NS�gƅs�н���J�]�LHt4I6.���ӝ�|���h(:��h-��e�J�ke�o�ŧ+��
ş��`�Q�vC��@rAрQ��5 ���v��g2�0�p�s�av*H���OK-���`�!��Kx�w_�孍��k8��-�5h�`�c����44�g$������-&3
�f ��e�{���k�����i3_f��з"�C�|8�����į4`+A��v,�8��3�b�q ��'�0Gf���eƁ�ǟ6�x�8��	ֶ`��_��-��>n_7j3t$ �m5F���r.���΂?~�5�j��O�r��q�QT�����Qmw��	& ����/��5�3!���#��	G�m��杦�F�ݗ@z��{��Go�K�L�H��K���ß�- I�	R�$cC^V�$Y���?rC������޽�d޸����po��?2�[����r����PK   ��!Y8�Z��(  �(  /   images/52e5cf08-beef-4b5f-967f-8676d3f3880a.png�(׉PNG

   IHDR   d   K   �"�   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  (�IDATx��}|�W�����WW�˒eɶ,�H���8�'N!$�&$������̓�f���ҲH�Tl���*ǖ���e��ۭo��|��˲�ya�?��~�|�93�93Gֻ>��p��Xa������^#�����X��[��ðd�z4�����Â���N�X�l�&;�Q�\ ����ڥ[pM���o-������`�{��y'Q"K3�X���V�#���+;��B���`�1C�ަo�� {��	.���E�c����D�e��v:S�6�Ug�Sð���8ÝnZOm1,�g&�%�u��{f]����ˋ��D8�+�6V  `f���<�ݎ��^����
���׆�G�QܾР��ߠ�琽�l�ȗ���^z��N STy���3c��l�Ə~�$�jԡ�~�^D�F�|�����<.�S�NYՀ�eW-�����/5lM��-]:��J4K1���u�9^Ùα*��e�ؽ�F��V�8J�3D2Rf���!	ܱ�W�ƊW���|�R�N�Q3�+��z/~�r��Q��N�@�ܗ�a�F?(�0�f�1��m}u�w�x�/pE���gՃp�v`�4g��.yn�\c��s��2�N}o�M_�7^�˵��_Ɗ�;�1��xeM*�������n�1�	�gMEm�����k2�ԗ+����X��-��̉ r�;� ����8�d�����2˝2�kR��Nk��"���0d�ZMeo�Z�ni��x<��hQp!���0�p�-�*�ܹ��#<P���Y���O�;$�1 ��ig�ak� �rm� /�˒{��Lf(}6�c��4���Z)�S�u�̈�I��k�g�O��av���O#4ԉo�&�f��#�Av1�h��j��@ԘM�j�H-�.� ���ү�hu�S_3y�ˤ���"�D��E%"{�&����l�G^�I�?Cg�����O����c}t:�ڇe�w��WpM:�_��G~W���j�/��;M'34y��,��5b���2kp16Y��F�\	���&g��1yyJ5F ny�-(�>*~�sSF�,�;�/����QX���%��s�F`T3�x3.��Kl����b�������QBΖ��v|�L�0���[n�	M-�ݍ�Y�8�W1��<x����=y�$kE�!�W�Nc4�E��s6�ܟCr�	t;"P?V{���F��ș���Ȥ�1	�ĸ�M�n��j��,�^��Pė���	�Y����k�`����Ϫ�G�ǉ3�UB_��)����gb6���-_��[��:˫l����3�]�� ��+��u�n��+��j�a��a�D�{�#֡��A1+$8�W��뇞���?IIID��49gQ����$�U� {rO��K�C��h}`*�����I�rZg�8Q���F��m�����<b�_D\�,�/l{I���ŷ�8&��l6���u��uXԛK��������s��~����1�9����k'��K���P�����0��.���8�'���v����.���v�f*��ϸ}�":��Ł�^)�C����!���<���xE���4�
�H�",P���j���X�ue",Q#3f�����*��F�YZ}ubf\� 6�_'O$��˱8�j4�֌��:�=����)���X&Y����k Q��;l�j��a���%��5-e%�*�WX�fpJR2��ٌ�Ɗ��&
���Ʋ�E�0W=��������ncs�Q�Y���!�_������"�����y^�jC$E��!���T]�9e���"�]�m��j�.]{E�N�۴���<U(�#�աT\PPz�:Ǣ,Έήf̝���B�eGB��_�����������S�����*�5��p�[������]�rQ"����ЯdB]�j8w谸�}B�>%!K��r�0k{o�#>�A�h��#xu���PQb�Z�k
���� �v���$��o��C��b�a�K��5���F���1�?_��y��P�������̨��W��~���JE{D'5��c���]���V,]�	9�/�Y.P�KrM���\���0贡�1�S{���(c��0��T�gH��)���4g'h����rx4Έ����n�j1�{Ĺ����n����X�x�2�^��w}�$.��Q^�QԪQݢX�:7�א{?�P�W<�8�zF�	��txƅ�!.��/��h����]�b��ȯ����n,xz̍솨���?뒅�=�!�B�$��ځ�H`��+�A@R����_��jn�D�[T/�\-��J�*��"���th��c߼��Z�1�[�M�����!v����}�{FMA[_4y�ީ� �D��144K�U$�Oj��rNn��m�@ThBD��ފ_4����wv,-O��E��4�j�$Gi�e��W��Ռ�D̕�%m��D!���ͬ���,/o��6JB�D�ho�O�(�ׄf_���?���g��,A��v.��T�Ѝo?}^���wbCV҄��x������*�A�"�^;d��Ć�y&k"nټ�ߍ���?�G=[����c�Q��nT՞C悥B�A�B��k},��{C�H0T��ҧC$R�0��_Gi�I�UҪU�L
�뵍j�+S�P�Hx�8�u:�v�GYޮ%�Dh���L`���dP�(��	S�g��a�����γ�{¬$l��.u�Ÿ�#����,s�ۆ�*��5`˦�bi�Cj2�I��U:l4��<����T�B�7�!�pW�C�5�!��`�I+�m������^�ώZ1�L�����.�&�Șv!~����s4Ѣ��I�ZJ։�� �;,��|���B���d��0�����+:�9���.���ߩ%�a�8�?J��{�C@hp�Jp���B�t
���4VS?��0�N ���GԽ>���3Y�	C'���cg&ʲڂ�6���	����$,@}C��yX��-"u�z!nC�����zv�.��!�~qc�&�E�B�ϥػ�����+�{�d��S�)4K���&�'�x~��k��+��,ܛ��,.d�Iܞ�6|�s�}����A!(o80aMdҤѽt�F�O.ਓ>��@ecs�H�l�<uC ��?�c�7z���!¢�fB�`�o��>^�up���}-�f�{�YM"��Tm�����,�7����}�|�|fJ�fd>�mSc������c(?BI�g�E��"���/м��N���_�Na�qq̈́���D��,�1U�oe��]�������
1�/�$F��'�V����V��B�x�f$�_ۀ^w�.�\{ϒ~^8���c 3j|_'W��#��H��B0G�L������G�x��4&_�Ͱ	a�����RT�����f2��Հ���~�X�t����9##D��
!�����&������)� �?9&����V���DEl���~���g��Z� ��)1���c�����N����g����]hҦ,��=������W��Tz�k����%�jV�Fc~��W�+_���*t�$�Ю�������1���y��iՏ"�=���߁/���m��V��s��>�R���i��کF���!�O������+5j";*}֪̍i���y�oO��|~�R�긞�6QM�Ѻ��3��ňN������엹:S�R�o����D��PQU�_D�h״�lܴ���C�s�9>����ziy%v�y��9ۼho�ǲ��8��o�%\�Ӣy,���z
�s��ݲH���4% �k)�M��;�7u�0��lM8z�ץjo�x�\���؆��!L``*�G�C��ft��m	��,���ic���cߘ���^����1"�߰p�A�#x*���@��t�͜'�$/h�\����v�՜M�:�o���jhh�o�ڦ$�g�@oo��cƨ�1*�%U�K,c�D��=�!�Q�WW�f"��-�>��+�9�h�Ck���:�x�^7y�R3�Е�b����N��
���rP����k�<�L(0k�Ȱ���|�����aD�:��M����x�%�=j�:�+�<W_4.,jz���#���ȢSV	�Fg�(z����R���	+�*�[���h8�,������%UB�9���֒������W��U��:��N��E:BƐIn�~šjM؝�ZJ���'3kX3�F�(T����=��D���(��Z�ѠӖ-_�ł�t��}���Bj���8<p���|r���wx� %���1�=���`ߋ���^,JOS��i@sSR��gę��6ek3�Ȉ/�V����żC����r�'�8|_��'r��MUC�E�����[DM�J���!ƶ�N(M�}�F0E��b~~L�5J�U)�9d��x�l"�����ۓ�Y�#,L{���љ�*�~n���^�2��"��ȯ8�fqz�3ͷv4�x��hlӋ\*jQsKX0/��bb�O����� &,��
.�"��(�]7W�+(���״[!^l�S���Xq@�O��ý�Z��<�=3Q�I�q���o��mu�7�7}^K�W7jw�Q?"3��S�]���s���z��q@�\� B��͚��EI���u���q�����z�%?�1Ô:�qq��*.*k���F�1�����ȍ4��
���y&�{���Ι]��/4e��"���u�+�����u�Eͩ'�gj��0�LL�ݫ��={����ŋ������2�?�!�@>{�1�)Ծ��菞��6�ϥ�"�����/U�y���ʑ�1a���a?�&Q<����fg�$�M�Z0�(c�k�D0�!3I7�.*�	vT ��y%9�4�����85�a��j_����w�w�b�Ix߽>&��5�j�tܭ��{ɏ��!y`K�P���+RB1��a��v���!}Ba!�b&ĪA��^=U�� F#��]�2�\|���}���j&M�S�=C-��4U�3u���Ѝ.w�z�K]���!�d�p��/k��h��y:�˕A:��ѫE'�i��0f��	z['ǋ���4�⼓L�;1'�H�°*�FTˀv�V���0y��b]}MҖd���I|��KbʤQ�0�^wD��{��Q#�kDl
�:I�����R��Rj(��r�2-^;�<g�M�	ĸ���:İ�z�q.� �_�� ��i��H����`�Ο��x���0�1e����nv"��݁��Dsw����^�fhgOl3�_�6�(Q��'����?�
J���\������_@OkД��#͂��3x�ZT7���:�=1щ~i�����Ѥ��$,9���0Q�.76۶avl8z{�ʱ����h>��[�p�������lc�=������7,8�VόjG���m��5��0�JQyIaס��Yi�R�G�H�3*���@y����b��Q`A6�\�a�6��$�QZ"b؃c�.]�ԌwWS�zT"���PTZ�7w��݁%i���?�����N踕!3�?�+������W��U7#��(�g^����ூ�/ᆆD��;/���4�i� ����P+�	�,
�~��wq��L��ߗ�����%�>�5�cXZyO�x-�*�6�O`�Xu����݊��oBqy��f�=B���xE��>��j��2B�Hٌ���&��Ivb�����*���f�^�r�d�q\�c㆕�����QVH� N�M|�������5�'��.*׭��g]C���N}M{8����ޤ:�I�q:�K&0d���j�Z�+oz�X�й:�D׫��Z��:	���Z��ܼ	Ͽ�t�P ���"v����~��œ�typX�y3�@9P6��yM�'{&�{�m6��:/��@�o�<���R�f�=0 U����~���@"3)�v�*�!X�O�vYx3��	���
^�Dq��y088�Ҳju��t�L�A��aJeY�RY�$f�x�u��fC�6(!\�`�|�Ik�R;B������Yw�>׳��FE�	��}٘�f��'"��O�����"��Њ�~]�;e�H/��t;�'�@�U?�|2�ʥړ�ę���F�%1v>��S1N�=-�f "ãq����{�l�q;X��G���/�x�6��<���z�)�Q�r9����:Q��EGļ�#R+qa�/cȞל���f�Y��gB��xf�>��^��>��k���\c���1����:_���j�=48\t��	1����bTbW�C0���'�}����V1�X���6��ڿ=SGg�bJ���J~����:���q��	�$}p�b�$lBgƖ�btV�Yztr�BprnA�^�r��Am"f�<.f��>�@�m4���B~rݞ3��gD8!\��3e�u�n�;-L����z��K�CBL~��>t����~��̸ ,2"�}�O�!J}��Gڼ��154W(G�fq�F���!��֛���mȬy��QJի�����ehܷ�na��HmG��w��Z"g�(Ӈ��@&���>�[�a&K�q�/W��u[��3���E&�j����,�c���t�~�i`at��=�VC2�[FKӀ�����As_.�+�A���U�:��]F��ybBJ)z`�I�<�2�?�)�WH+{�F�N�!S�[������X��QT*8܆��a�3�(%�Z���7�!A��4 f2h�5w� #���?6��Bf5Vu�F��r˥�V����ͬ�:;�×�`���*��b��n{t�aEZ��P:�f��H�ۃ��8�o~['9d,\�O|v�bV|L
���A�=�W�O}��j�q�V�a��kBٙR�]�U][�%31ٚ�q��ho-��
�[���#hw'�$�N��G�2�5gl���s�����X�Tܪg1�m)\|��bN��bJ��=f�:��Ix�#C_��ҏ�zb�=���D;�k��0G�>�O_���l�OK��c_������3�0��n�U�f�ݽ��O1T�!Ǡ�fH�<�{j_ŗ����,
�1��B`�u�k{=��������p�"���᝕
�y��d4�O�*�f8�`d��\q0#�E��zڊ�&�;Ž�|��0��W��C_��U3�yY\��-0<s�쯰�1#S]d^��[�S~�?�^�T�$�eI�M��sʪNa���uRǐ[��j4�V�o ��暻џ�;����i�YC��E�y�L�t������b���:�Sy�@������;��AT���z�m  `����6�jcdnH�SlN�����X4�{�1���_�v�3n,]��LGz� ^a���`�U�#��8�/t�Ԯ���N��9�J�
KK`��}v�Љ�d
cWDBL%qO֙ZJ�[)*�Q���q6�UܾD���k1�g=z����mn��E�C�Qۡ�����m�}Z�����;3���t-���w��(XPG�Ck��q�Xv}J@AnA�7D�h����v~̵~�n�����r�ۤr��hD�u!D=$��bU;�F����C�&��� �>q^���]fM �K�i�8ۙdǢ_��-5�i��O�0N�ɩ<���M[��3j���_�_��`;J뺐�~���=]�^�Uf����ݓ���ˏ#y��1W��������g>�����|��i��YN#M5E��@�x%Q�xG� ��j_%��U�n�-z,:*�6��k��{���И娶����P��U�=x`�i�=8(�nZ���lO�<�}䗕(?�y��?}7���ba�*�����_BF�#��z�j܆<tT֟�aZTyث��,���CVou�c�'�0?�[�u��3���_n2�i�TҲe�Dm0j���XF�ݩ��F`��p���O���6���A���J}Z.S,��������o��R��AN�(߇�E��7a�
Ћ���9���A�;��3�y��
��np�V�	��5��{+�l�֮Tg�=�!-	ĴP� ��|{�NR���������E�xփ���[�i[����6���~��̺E�2>�3��k���ߝ�x����)�8��M:ld�����X�3�J����9��P̜��Mhj��"��!Dl���q��\?�J˟�+T�N8c����	C��l�Boը���������W��^:��4O�-�|n� �P�k�Ƅ���:��Ħmb1Oe�.%S��K���}M&�u���gr������9����1�/�e��� �)��������)�İcb9Bo_;�SW*ߗ�9�!��!Nq�Ox�!K��kXQ^�X�N�a�&K��x�Pg�c�FD�� ����,(�Aǐ�T5q:|B�M�4��)��1'���PF$f���[�A%dI��� V���=ϞČ�}�x��Dh?�$���׾���Y�	p���Iz�~��X��5��D��L4��M3K�׬��%X��Z�}x�_��!��^��=�S�#';�)sN��ز�,�D�Ij���y��:��I"�|"+�t	a�{��П`�>1�?�|i���oL�e��?QyW�V�*&dѪ�q3�ۯ��'Mח0��,L���&S}e$i�}!�Kf$Ħ`n�b��[�U�R�T�3�?~������Z����g��F�bV^��r'�.}U��=�̆e�3㤤"w�9��ފ��
nѡ�7�X��3a豧�oލ����Db3��*�.�Җ<%��_6j�R��r]��U��1"2J�DO\Y����=q�7h�v�\Jg��^�R��Ct�;���a�FX,"��@��J�����X��v���S����Է�*[���}]���/T�����ůE��cn�u�V�֜Ņ�=|�e��������{�â��[U)@��U���+A�Q���/#���Ȟ�V�����Zq�sf�s�T���j!Ɖ&m�N��t�e����xM����8���ɭ��p����p�U��x���٢�2��'N�:��v��Twp-_��h:~y3�Q�%	�ڳK�l=�ްTU:�nߺ˸���e�O��9Ah���e�4�J^�����ɍ��y��gy�)��Dt�I�C�B���;��?�O�7�F5���w��c�b����+�"oYC1<܋����m1�^��N��ş+,�"[tSkN?mV��wU����$ﰊ9�P5�m�#L�Xt�8&PlN�ط�0����D�zվ�%��"Fbe܉�z�5��*��|7ӠEg����jtd�;.&���)��ܢ�����V�lR\*nY�)u������~�*�f�NHSu�O��M���εrl���:���a�㈊��lQh�w�;~���U^+k����Q��"����D��+��$���c�cغqn��~|�gU^,70n��V�'}�"|��Ư����z�z��~��1�3$8�]=S����	�CK*?���H��Yiظ�C�6m]u�l(��ի ���f�RrO��d#M ��-�w�%��M��ܗ��`16o�G8��|BJ�jdgnF��7���n�GO�Y='����K_X���nxހ0�IY%Nf R�E���hi��M[�����K`4�^�1��.�O��s{1�bѢ�(m�bb��7PTvr�-çj2x떭��;�9��p�n����ӯ���R�h���P�xu|���J�[����^P��K�_�uӇ�:7K��q�A��@G�HG-�ˎ"5%K�������/��)/�P�S��ՄsE�Z��/���������m���Ƶ���[{��yYJ2"��p��P�߭�3*2A$�Om�7?eBB"�At�sl��c��PP�#ؾ�'7��	y�yHΰ#���58�~�V�X�x���T��w��>���
o�������V�<���ܡ��,#��0�v2o'N�ۥ��p �n��ٮ�PO_7
Ks/.G�$�ϼ�Mu�N��)H$9a��xi�c�2o_���3t	����ǟ��ړ�������g���"2"^]38ԋs����dz^�>Ũ����Y��0�Ezٴ��m5��j���
2�7F��s�Oi�[V؏�f��+��O�����!NZ� �v
i��HW����4�x���������knR�;���Dea�!O�c�|�Uklr�Ш��|�z���g+]��u-�:�����c=���Wl�ʢ�����C-�����J��_6��<E�1    IEND�B`�PK   ��!Y����+  J  /   images/5644ca41-1cf6-484a-bb07-c2f9a6f5b19b.png�WW0 �]-�+D��DM6DKV�Ѣ����Al"�Z���$z����:��V!z�������g�=3w���=�:Z*T��  ����[��E6ٝ�L]�{K@OUco ��� �����|�`>z>k/{ ����x�Z{�xx9��J=  @Sj�r�o3v́�I�L��S�g@`
�\���EG�T<e!�����DʲϘ��|���E-	:3עt�&^7Cx�-��
H%TH��!�U����������C��ח��(���~�|����>��`����e�~�L����E`"#�n�����bng��0�d�w��f��u���R?	X_�B����������`؂v�r��I���ӑ1��ԙ��*3~��_��:a���skZ8��[;��"���� ���p�HZ�������1�d���g/ǚxx���L�	K��%y&�Zt�Q�� PKI�!����O�Z��k�>)�|yX@8ҳ�́ߖ�N��+a�i��?���m�ޢ�[e�O�M�����"si�n�4{f�g��!l�4eqz� 4W �J��(����3=�ͤ�;[AI=�� �Z�G�'�Ci�55���T�eqo�Z�K��T���/���m�p��&�5��(��sց�ѽ��;�:���v��F3��� 氉2��G�;H��1��"�{I6WY�#�JJJZZo����gKJ]����p�Y�*�`��&���i��&�k}pp���F�oʡ�t ���>�x���n�3c�ºk�����Vq�[˛���ai�ɢ�L�7~@�ĩb5�W����`S�O�=�\"�����j��oq[��Z�ޛ��~z�G��/��G��)����Ci�h�k����i{(z��_�zģҕSD�i�����SO���"҉5\�^QY�u��6W-"RoMaJ�`:��󸼝�@�&�GH(��3wkװH<2�wgv�9���>�M(�Ѱܢ�k	u��WKJN>��`�i�꒬����Bfxn'�R��c`P1o�9��T��E̵��h�ޑ�OZO��F~��nL,"�h��UO�����`�}�p�P$v�"%Ʈ�Y7;�>��B��Q�2��'�З��>Q���ߨ�|��>SU &N	�}�C��<&�uDi�ƴ'�5_��i��H��dƱ\�7�[�i�^�6WŊ6G�M*U����o�c|��3��g��4jf4�퀋�Da���B�h�bs�H��Lu���_b}���p��9�ib�h�Hm���I���� ��w~�:�Ǚ��(�Z���iaa��-%�X�0n���4�S�P+ҙ=ߊ����D��BmvI�Mm>���}K��A�U���q���LyKHk&��MjB��}���A�f�)���D}�ü����{����h���xܞJ�tW�&P=�a�kw�m_,#����rׇ�߶<J��V�vg���^���ҵO4 ����l�IGB��L��PS��ڽ�����	�;m�y�}a�.��%\o�jͧ�g�# lF�<���s\RCj�ch.�5O</[ߖR�̔��{o�Zwu��H�UV�E���_�#>��N����1�+��Ġ�E٫�ͺ���vub��Vt���9c�M�j]�򏻏aj�(p$v&�99�r�ئ(��J��Y&躙l��u-�1�}x9��x�=Y��絗�<D���T͢Mxf6���Ȉo�����{�W�������fF��Oʁ�����w�7���C�f�<�{a��ḡ|̴n����*��V̶Q�$��e���YWc8���dO΍��$V� =�z�z��!�Nj��8�H|������~@�����;/4��ʽ}�Btnb��D��WsV�_዁�tPY"ۃ�t�����P��~/�9žcT��bQ�F���n�}kM�F=��(&�����<�{�W���i�1Ӣ3F\QJ�"�i3���%��1�ixjF��aƓ��r�*:H�s�Q�"�@�g�����������$-x��d�۴�D,hO$LDRS{�T����ib�7�G6CK/X���7�ɣ� �)��֚��tWDE��+�9��R�dV\�Ѽ����E���X�;+�[���P�a�Ze�J-s3�~v#sA�;~�sDh	.l�//��ܦ�:�S���Ż��|������ᬹ��FO�����h1 W�f�V��e%����\+C�p��T�8�wʄ1���l�5k�a6�|z��j��������2�zX��:�ϳ9	���P�������@�UlA��0Ԥ����\[j�4�r4�j:UOz����'y)c5�����;�u.S�����t�i��p�*y�0ؾT;bg2015A?�Wj�l��ۢ�$1ye��K�����E�^-����T0���8��� ��p��a
�`h*�Nj`���S�^N���dB�@#�*N�CK����9���R���૕V��v@cy�;�K��z/:�,Xi6S|��궣���M��v]�� &)��\�4���9h����_T����,��u��=�n2�O�R$گ�[?&̽�W���'����>�޸��R��q�ݐsW�t�)���9RqP�`��]�
� }5
B����g	k��g��wf�Hf�1bt��}����8��c�N,���.��)��֩LS ���5���梓EjP�r
|-�������q����F�(���5,�y@� g���Z WMP�;�,8#�]$.%'g�^��!��.�x-z�\��������NQ�{�zAz���Qr�����-wT�1�,T��r��5:}�R��`Ha�ځ_��K��������`��s7}��3���ڑ_�129kzV�0��� ;�#+w7�p�i���L������ xT{�^W(qm���_N@xGY׿�<�F�^�FNz079[WE�D����i5��n����a�Į<�={�ܕ���V�i���ܬ�K��$�GȰ��ץ8IU5�D:9��W�Ռ�,!���%l{)�8Do�P�H�~5(�\@��S�mmu�e�m�ڥs��>+��ڃ	:=s�Cl���Q�X�f	Ǒ�V��a�<Z�5#u&r8▴ ���c����~��?�j����Q�EB���C��C:��h��a��L�І������l�z,.���'1yiV���F?��K��.ϱ����"�lC�&A�{>�v݂���`Ԏ��:���<��Pj(_�q�e�E}��*Sy�ţ��)�E��k�����N>�a��Ȼ�U�Mċys|���_�֕�d�.#pѫ��4d1�&@�h�[�Q�����仚b.��W����M��R�k9�FY=�t�fn<O%����\j�l���t�r+�����Ñ��T�(E�@D�����3jbT��hy��b��A�`j	�\)�v0�	Ăl�r]�_��_�%K��*����d�PS���ſɅ�.��{ӕ�#�X���b�\6��K�g��,id�dQ7�o�|#�p���JN��w��
F�$L���2-x�s��`�
�,"#���ށ��1'Э��x>���
#����-�|a�M��^Zօ�Q����q��>��Ւ����v�Ur ,��[���t���(dN��z*�Vvq��}zR���j�fC�;<he>��4�d�R��f�Jso���|���_����|	.���۷�R1?����#�<=���	�of�d���{�-����k}2`Q�5�����/���q���w���t�B��a�˳� N��%y�{�es!}̰B�crY�	5C���ņ-5+z �!�K��U��9i��hE��������$M:a��Y�UmW���JU������R���)�\�Z�~[O��-#���b���T��\p�������O���h�_�fR��L�����WNs��B����z���{Xc"]���oMe�X-��sī�M�`��E������[���Y�T��0�:������ϟ?�=�
^p�>f��ݚ�4v1>�^���f��"ȴ0��^�f���J�j�M�ZŐS_B�M�/�������c;��[�sCT��#�܆���b���?PK   ��!Y}�� � /   images/5874d651-dcf0-4a98-b8b4-9fcbfdf83d7f.png��uTT��=�t7� !�ҍ" "�4JwwR�"�-R"��� ���!!�\����~�y�ǵX,f�9�v|�{�c���L424��TNFA��@��P�Wx\+�/DG��j(���Q0��NN��l��������I�d5�TmM�\��!�����6����v�����"d5䩌��[�n��N�kҭ��8&	?�w�����xXh�j�y�{����B3J;���Њ�4-� ;I���TJ+S�|�9���S��������P�L��2��>S_�D�Ǌ���>��l��ڟ���ڸ�*�������tq1dOɑ�Å�_�@��/�� �(��H�ER8v�):������W����W ��D���ӧ"�����E�"Dl;H0\�~����`�(��S���ʜ��*	gy����<�J�9�ڍDf
9::jqlhدv8o�}?ޡx.��r8��4�>�7�ӧ����ĺ���%�!�#�p�_F�O��?הa�e��p5�\N����o*˵�ru�av
�܊<~�$Ѧ��!���>ʈ5't";���Vd��+e�U�̛��[o�z��-~����,ٰ�ή�ᱱ��EO���<���II��ZcY���cn��t"")[�$��B��Jů��He�HeF��7
K�Zs������4����W������a���A�j�$���[�9v�����:�ܽ��)w��]+C+/�9�9���_vv8�z�����#"�N����&[�$$(>>>���0tsK��H|���� 9����v�Ņ �e�;�";
���2V�7u�����X����Û��t�{���#�ө�����~������9��U~2t�S��qer�&��m�͎���\Q$�i؜���GV�1��a�747���)�,���>Ө9y�K�a����x{��5�H�W<� �}��U��C���f�|����H�K���j4t�2zT�Q�� �ř�([���Z�d~[��xH�	����#>�94�#�ݏ�#��E`�t}�_(��[���AXVV�4D`0��X�*`hhx�w�{G4Gӛ:�W�{{"W��E����(�Fx�񀄖�B����F���2�H1'Vb*Eے�������n���_Qg�%��������������7"aSu
�6FhW��������'�Q�i��RjF��t�մ8(PUÎ�Xp]h_
�M����Ѽ{h5��0!���(�|�QØh{���̇=9Cp�Џ�U�:�8լX�"�Dǋ�/���V"�a�Ѻ�p4:�\��\������=*[&�R``�;���ڻۓ��ۃƾׯ&d"�k����\�L�[Z��+�lܲPsK�#
�B!�б���/��
ܳpѡ��g����O�9��,�ϟhy�YDT^l�&��v�1�3KJH@����=b�!�x�W��ގ8�Vv�22��ʦ�ϙ������w7������� ��}�T%����^iH��dL�p��w:	���-�0�C|�׷�=��rxt�Rо��#$,�h�2X�v�iM���8����{P˛��>��|l�`�S���۾���?~� �GY]�	V�m��� ��{�[�i��Ԑ�^E`z�FF[.��DHe;:����p|����-���'ևn"`+1w(�����|jvU��zFu�p���f�M���3�LW{���Ɓ>��HD���@b����.d�X�xv̬0p:�ap���K+9Qs�I1<�e�bw9jW�{��	7�������l�@	�"���x��MJ�Ch�b�[����alw������̒C�\c̉����ꗱ�^�A����A��1�R��3�}j..\p�23ǘ�X�}qlme$�}YC}����YF).|uqA�������f'a,��zjc���(�wO��h�k�fH���sj�Ȯ�0���]+�;`ە���#2%��\���|�\vgQ_�~{[__?J>w���~����B���v��B�M.~���G�����c���P�;ع3�F�lmm}..���2���\:��̅vLWZ�rƑ�6�XQ�͊��;^N��͙��x�60�&	r�=||��������?m9k�ˈ��n�d��dVW��z��
_	,��2��îT���&V>sb'��U�cAA�S#���%
TZ��2#�����Đk?/�_e�r�~:%���+-'����LN�y��ׇ^`^ Z�А.1���!CM;	�{׋��׷[����d �M�9�`r"w�'���tF�X���$F���8V��2����q$be��ȱ(o:8���0D���10��J��Ky�6 _]On߷� �
�����ʏG��F����	�F��
J>�i}3�YQ�Ъ�93s�4����R���Q�Z���$��0ځ��vH�'\�cx�f���ke-)�Ar�.S,�Xy'��Vw�<A�m�%��7�+�D�$�/��>��o��ڙ9GD����c����uq��� �H�>��ͮm��!8?����7ܕ�N�~��,*5��@ "�������1ۢ]x�}zH���ST%J^t��:>b�`��h�=��{চ	�磌qs[�=�6�)��F�ρ�����l�58�S�u\�T"Vo�r�D�V��a�g�S�뛛��^����rG99��^g�*+RpDࣴ�mow��g\w���֡���iiz)��S�R�8ʪ��F�`�5:::8��mq�/e��jNK��	ؤJ��r$kʆ�����x�����<�,��Ё��B�#��F�\��~����{qq�����B�lm������������f	&������> M�/3��ǮV�I��͉�� �\�1w��Gd�%D� "GD�+����.i�n/����ĸ���'v����FL�pl��\��b�2���%������9@q#{�9�F��- ��������)���K��x�Wg�_��xG��C���"������R���qG�k�X��jݖ{W;#V� �V"��466�9�����J�iۣ2uݭ�1D:]�xo�Z0M�..R�X�V���a�
ҝ��B�DI���UTZڇVZ����A'vI����#�YҀ�V�7�u_�x�����+C��~�u����ˇ0isR�E�����v��7��Wk+F.i��h����aD��%�FO˓�F�Mu�S��;�����P�2z@��� $,��i�v��D����ʅH��������5Z���g���q���܌�OJ�0_ƅ�V��qC*W%���+���ґ� D[�'Z�˽���q�{x�><�����@x_b��w�6 ((��Q*sH.��#��ox�"����k\�
	}."��ow�+퇺���++k����۳��^j/��-����M� �T�̵̿Ŧ�.�6��H$���Q@�yη,�G���d��l�2#ԽQQQ&6����w��X����^2]Cw���������zz�_���aW�T|�_�����
�n���Aa��^R��%u��rE���o�>����)�$�`,�rG����������n(�]s�v�D��ڱ�ӖKLl��28[�	U�~�LӲ��eq(
�΀X���E�Ivv���A���1=�� U��F�9*Z�n���/K��tϕ:�����5���qS Ѕ}�L#��LVA�H���z�N���Gm_�
ت?DF�,
#�_��~��(_��t������,����7-�sҘR�QF̑v�P_W����̵?�N�*���Gô�����V��s
h��\��*Qhӹ���l9�B���E��FL �#{;���`$�XegE��'�A����j5�*cq�L���iK_L�^p��J�efF���@u܀�smb�P����R����T�j��s�� �(�Q%�`�,l�o�p��(Z���G#��ko$���5���O�S/,y�����V��G�j� ������,�˗�].dc��HlqEmǓ�g��E��S��k��Z2W v{+�tj�:�'�����;���;����K�3�y�J�����s5�}��v�'e6�S��S�=��(�4�B¯�]3�g3�_H��+)����JQS	/H�=e�qt�''5����k�}�������4��"fd8s���'��i����_1����|�Nz`��I���(���r�R̋y�;�%�'O��4�uR�Cl��po�����F��v�$�I'��P��^+~i�<GO��L	��(n�J���"I�� q�w�@b�!w��қ�Q�O���ȯ�'溷]]]G�;���įj�]����c��0����F�l�-!�R���)��Y��;�sy9���c��7³l��߮c�V�8t�b7J����b�<����шCu{�������Ro������b��R�	�\޼��sR2kܳJ/�n��g�����iu�8���dvּ6�,�A�Ϫ�Z�FFFovά]:���A^Xy4(�g9��iɟ�9����͕p�I1�z7c�٘���ō��g@j���N�6��.����A�!>��X�m��P�P�p���C�ί���
ö��^��C{HjY�+�G/�)` p�(9�
>�<~3��ccF�NJz}��B�Rf��J���K��x6b n=�>����Q_��뵉R7�ت�7�nQ�Q��*��w*�@�;��J2dI�n����	����l���"��itX>� |)�Yn��}2[~xvVuU7f��sw9xy~�V�@��j� h��?	{�+)�3O.��+|x��>腖��dAp��@��_^b�=[� 6��>���v����A�	������;l�cU�g�E��/��vU\}س�<e��GqC�7�,�X���c��s&��'���K~���H��!·�=S����D!��caHC��ΐRQ=y��P�(��q�'O�Dh���v�՛]$_���{�/UE�G^p�*F�(��n�waMp���08���T�>Y��/:�FjYR�����%���z�������|�7��,+{Tǿ..$rU���pR)��Hb?��g-�����"������r���tEJ�Qg��*�G�pnb�қ�8W<S����G��	��|����.�Y?����kϑ��7����H]��.++�r�	�Q��&`ߑDi�W�a i,� hcE�T��k}�G��ܾ+�H}5��h�I�|�g�����"�G]}�����\=�g�Pxti)�<��ok}�E��ֲ�zM3�ń��b	c��ƈ��05u�U^�O̮��s�ԃ��������.$��|��b��-<櫨�����Ф\[�a��RN���P(8M �#yE�vK��c6>��(�)6�"pYr��0��m�U��tP�^;=u2㴝o`�ľ�Ùw�q�n�r�Q�����v��)M�h	�xi[�7��L7�g�	l�L>J��6$��IF�N�,س�ۿr��^�C.�W�8�I�_���q�r�T����2Y#���!#�:'7?��
�El�p��vu�E�.V*Z�v&JW�D=EvQ2Ġ��Ų��P^ϱ��ѱ��5V�:3\�5!!�tsA�k/�5����'���1d:���r6Wz��/��~�4���m�s�'ܺBBBC��Y`:'�������$Y��2&�sm`�@F;��\�����#��@�9���'�� Ƙ���د �~�s���ӕ�/7~lg~��q%�yt{�=Jb��<o�J�,-�����6�(QQ	����q��_?w�&���Gy𸙒��8EDVW���cХ��J������7�\����Qn��� ؉C�X�T/��4�J���ۭ������O�=$
+���Nq��ơ��tu��!U؜c�����g��=/ZtĲ�+;W���*i�CB���A���圼#^H�H����Q�c���J��[or���ML ˆ����*�ZIڔn�`��lfB�f�|��� ����m���B}��~�ÀAK���""�af�q��Q��[�&����mS�`́Noϡ�N��Z0&0�=�a|��`V� "l�I��6��bx�k�����R����ޤ`�f�'nל���le_���  ���n���uTjjD�>�����(V���):)���Q���^�k��@'���r`�'c"8~�� ������7�?w&H���C""_v�FE1[~�����r�^xddvݗ�}��/DÕO��U�Jq����/�u�H�����Ag��&'���h��x����f�uc�,��uYq?¼�ȶw^D��<'*MJ"��S�+'/���9""�摰��H�f���y)�����|�ڱ�;�@�e�Fޅ88���~	ǘ�P��=Ïq�;8�m�H���T�r���4JP�^f/������nb7�wi%�&"��ӑP���~��222sd���qh�33s�z���^hV1))�o^Nf��nx���iFf�C ��؂�3EE�,�,�����6\4\p��*��\�q��yl�
1qThdR{Q��,��P�y0]�K.�)"ei���'So���ϟ�lY���P?�K��-�+�k�a�k�L�eՄ׭��B�ٶ�Q�v���d����^**��������$	�&zF4��%��R��/��ڲ2.r�=����n����#U���Xl44���l�%���8�N��/&'�L-�&7�7������*���#ɐn=--2��ǝ��eo1�����dޡ���%�IP�h�;Q�ö7���)9(�>��0RԐ�w���R�ꋟ�^A�G�KӲ"Us����R�ۯj��������e�1H�'���V�u})�d����g���lhHW|�F��}	؎�t) ЍS�����rOl��]F�.����Rhb�ع�M�z������O4k��_L���1u�u-F��/�p��I�!'��>==}.��]2�&VC�F�)�mV�E��Ѽ��{��`�����h�j��
�r��)�|b�WV3G{�m���ρ�i����d@9��|�R��J�\�z�~��/�s��4h+�a�ʠ�m���9�3GU�{�Ȍ���%��HR�d�w�7ㅈ-'JR����� ]^��-�x
��L렗�[��v�*|�~�'���Y�q�|ͩ�ݩr3[� ڵ+?���$Κ�#[[[+���� ?�r!�VǑ"� �,h��� ���Zeァ���rG��.Da�M�	��. �ֵ��6�j��T
<���T�O����VVV�V~N���&
'��g�<����U�;4E��	�>.���9Pıi?�l�����L�$�"���������0'���A�b�(�`���~@dd���S<^�O�*o�pg�M�fX��t���$��h�BA��c'�Ta~��h�2]C_�ݣU-�Q5��n �'��9�}��6Y}�2�G)�����L�G����
Q4��8��'^����١P�Ĉ}P�iş�SӞ=R�k�˙\��6Ei�Œ�Z��3���Q�A��z^�зN��ݬ����:p�̲�%miT���k`�vu����'����z7���bC�x9%���F�
���>�S�*�4]�s�'b@\�L,�]����^��Dǥ��2,�t��:��u�wrq��P�#��(���@EE�Y�!&fVy�3U�A��خW��U��<�q^e(:�ي ^�2��ޓ�;?:¿����?FZhn��#��Q�O�v�J���^�i	Uv��������2��mJ&6�Zݎ-�|�޾o������𾤅�[Q�N۫X�����>�D�r?9.bj�jM�#k%��5�a�]T��ߨ�F5��[_T���*"�@�_@ ��r�j�]��&��5��]��������yd�?� wd�`(T <����Pl
�~���E�ݎ�x���J���F���J j�����_����U�=�X�� ((8���6Ez�t}R��*��5� �'�%Q��r����61���e� �G%=����yp�I(2Gs�w�B6��sm7e�^����o�,��x��_�z�C�k��j�/�;B�*��$%%��?y��ؗvw���r�.ǒ/2eFqY[K�
c�d����h@Ӽ����`�Z{z7韮R�;<H�c�P>Yv�4ޙI���r������459+���z(�����	/��}�M���^[W����kI��1=�I��L�W�h�� `e�|�����+�Ս��wU5�'YX ��\�AS���c�DEZ�/v��"7���5��7��ֺ�J�T��`�F��P��ڷ?e&��*��n�y�㘀k\?���Za$��^��������z�]#���47��	��xEu5��ԍo��<�������8C��iE�Y���F����ZYm3�K��.rs����W�$���j�DO���v�@$*3���L\�#�-��~��4G�"��wdإ������2� 33���X�ssv�Ł5�����=�ͱٻ�����E)�̓E�i�%C��}M>iP�c_7�ӠB�ש�A��+��wP�f�%RQ�682���e��n��j�jl__�0us�� wxPm��!���&�ӽ�An������;NO+� J�zN[����w���D�vq�v�������ވ����r��3%�����t���i����y#I�/�q�������ʝ�	S�	�|hh��N�h��Ѳ,y��ɣ��pӯ$&M-*5܂VjD?P	�����J�/�K����������$pt����1_�e�N�;���sWS�k�5�R���!���
�og 
�w(v����x/1���{����3Qqsۏ�A��2�߶�GI�osK�'��
L��
��R�����%"<ܧ��Ъ���M%@�5�*���k%�ۺ����ommIJ�E `F
I���GX�O�4���<x	]�	�ry��b�fI=_��!�nC@I	��[��mԬ����R�"f��L��j����]O��?`�����3bO�N�Jx��l�8��&<�r�i�#p����0R�;��A5"@�K17�����]�P*'���H;��G� .��A��A��)�_S}ǣ'W!NB��)sK22��R(����@k���4�i��֙�В룟?eK��lJ2�(;d�PA��bѮ�[�#��V���9��)����5�j���+5�Iܕ�Ca�Ė}��c�����p��]��wP1-���c&����QP�1�@-��|d����cS�r������w���D(�Nb�<���Ͼ�мqR��Vi9�c\�����xe�)�&]��@�q�8�Jč���s��s�����[�nR �Q00r��A$42��p`�AAG�W{蜈`���@�744���/"CV���x�;�골�DDȍׄ�)D�+����9���uLK��}���1X�MD�2���e��������8
..._W즰��6dvG�>��v�(�����N�;�GP.;�/��˸�P�ڐ~,,PiNMqV&�8?~|���>�
�&��!q򘞀�}&����@��{�-�&���Ѹ��eè��� 
��܆�(~w����>�VM%B%��:��1���01�?�����{jD���|�ѨPC�Ͱ�䃬�D��>���~l}���"�\w�L��k��L$����f��b�i(jK�x|J֗2���%'#5�%�d����-�v���DX2[�~@�EL�}����n��m޾��EG�G,֎�.���:�������i:�'�cY$C\rr�j�o���Ȓ�`�T׋����{d�pU�=��&��ؽ{� �[[�R���t^A��D��C�{�������7\Rrr*H�'�_�^����Pf}Y����*���$�^~~���n�<
$4��~��o��8 z��|g����MK��G24�<-��.
�H��Ҭ�����q� Byoq�$&����8���pII���XYax��
�{��I/T/��6#4�f���gh��Q�k_�pwF���H� �{+W��H��PrM�zr��L���:�X>s�.Zu�q�`��
#dQ?=?�{�̠���{f�
X�NK�Rn:���zґZ������{"Xs��ۑ�;�33��Ƣ[���	�,�
�Y����Z�c8��D+���#��iO�Cv?@"��^�$t�掯�1�?�J�徊��FgfX�quE�"�Πz���K�j�����g+�ܧ��XH-�QO"UǺ�?������jq} Y@˝ �Tp��u����H��,��y�M5�4��7x��Ѽ� �m�T���PK~��w����<؛I.i,�+�z6�@Jj��I�o' �P��ٸ�OXũ;�Zq�4:1V>]�L�#��#iA��zt�ЭZ���ݔ&B^Y����A�+����������oYx
��c]�ӿ�&hik6J,���6 S���29�y�)~G�ŋ�����?U�{��.^e?3Q؋�cc�d���8�2��z-���b���+��V��z"n�--��x���lp�ԯomy�4��0R\)ل���=B)E��c�W>��b���xGI�(�ܘ)	�iॼ���>0H䖏��p���lgJh���r��j/_
ꭟ��9&�TT�	���H���m�e����zNM������CT����܎���i�<�������^��ZgW��
4t"V���9�S���»*,�/��!6�b����|�LF4�K�a%�"�^���!G��O��x�����\���;�(��)�+�Y׻��e1z�,��_��H���%�H�Jo i��0(=*��w�`���9����@}��~о�1���~��v�*RkO�ײV�]mw��z8D��W߼ޠ�"��apE�;ަ�Ĵ�X�7��FT��@ ��g�����	�T�ssfff2�HU�*����ֹ�d3���nPr La9/�ڦA���],|S�zH�����v��G1���I#��R�.''Ŀ�]Ϊ������h9�Z8C6a�; �Wvz�\��U�l1���m�� � &�n��Y�����������Q��:�c�[|��Yf��-�c��̃{�Qd��r�((y��Ϟ��V�W
��c�AP������������Q�}�Y*���ud[u�u���?��ؒ' y�|[��O:R@:ý�����R�tѥ��3Y&h��V�OJ�4'YK��ube�w��yy겖M;� ��mqݚ��o�V�4s[s��5�����*�f�"��[����ZOEHʟ!;K|A�X�յ��3ll���t�A��.'H�1�J˝�Q�9��<�A�6��"����V�߷o�f��Yܹ��mmm��tt����w�E_�s�sQ�(>���N8$�X"�}- y�w�ki/-��?�zN��7�])�]�{�ď�_X��� ��l�V�N�!��tq��IF��K����dS�utpwf{1�-f�`Z6f�W�Z�$��p;�Lr��|��e6���>#n���F�;�+
x_�7\,�J���L~�F8\��qؾ��q�O�O��hDD�~�"M7\�(�k���,
�׾��2�P��1ړ��`�Tb?�G��^b��on6�����Q�RS�_S�x��*���466r�Xd(w�V���R��k:/�
Y���_����=ϗ�a���	V3�2���c$Y��$��N!���aYR�������U�H��ಣEק�o$�z�G.���3W�r#�j^hNnn�v�6+�4P.[A�Fܒů3�/�y�^�#�O�M�hkh2��ږ���� [_�
$E[��9(/��5A�A~��j#�%B��d����ט-�Ĺ*������yT��/������ī�7��fhv��c[��s���ED�=}�H/��G�Z��&��^0%(,��;�ϑM�d��US�d@ڙ���g꠳���*DeV(*$�ߛ$2��K��脄U;��>BN��"{��#�������I�����H�����7u�Zd;q�t�L*j�LO��]{�b���U/ёt~I��HC)���$X1�Yĳ"{��}�G��F�H�|[���r�;�n:pPS蘗����m�&��1*7"R����o��Q5뇪��@���ǒ��P�rG���6s|ǩi�j���!@�x4����N�	�Q���� �i8;�2����g�w�+�J�k��TQ���4GC�f���6��7<�[h�����j܎h-���fHR�L�}���q��qH��#�g�D�g�2�Dt�6�J�"�;>Of�K��6��It8q ���=�K�!����UX�~�-�
�����Q)E`IY���"�0�8g(_�ɻ��+(�F���3]k
 Z��߬�M�3>r�;<>������o^�;<|�	�.ۡǚݿ�������e`�Q�.:3��_T�C
̟?�_��100�_���ԣ� NBF&����V��H���l+�W���	��^��F���I�
ṕ4g���~j��W����I��S5TO��  �rV��`���:�D���EԀC�r���Cǀ �[J
��%p]ꌸ��賄\��7ɖ4��w @ �`s[M�)&M��ڏL��KJ#�!y].�E��G��q�`\��)%�z��& $���x�����<�-��ޛ���Mo_S~Qi�_�5�t�^����s���W�
�_�J��'Z��p>��ɎWK�����
d�wYTf55Q�ѵ�9mj�%�ZF<��������@S~�oP��̅9!����.���O`�+#�z]r�mV�$��c$�NL���M_���cL���~yr���p�����%������ ���f A7��*�Rϟs@y�̈��/��<{]WN�L�Z��C��4����~��h|�'�f����2���	(��|��8`uc#(V���ҿ���_��ל�i���ۃ'��y� Ѯt}�cy�� Z���3̕Ax������	5��2*�F�����$��t����,�8�?DެEXN�dj�$%�1�% ��I��3g7�:N#��k��S�^�(V�020�f��a�T���AA�+����I�YV��(/R`�����Ŀj���)V\I0�m7;��L;� �)�"����`ɿ����g
�߶FRh�$X�0��qb�V����F�oF3W=_?��*�.	�J!��Ӻ�߷I����T��gR���X�@;F'!��؀f��'����!�!#+K��p��AE��ŗ @̋^�ߞ`SE��i�e��^�ln���K��,r�!2C[�e��ޑ���9̟%:�����l�g �RJ;r,&QIIq���h��Q;2�S��/�.I�c2�N�H��T�_��
�Z��05��u��?e�h��� ��X���?]�γ	Vv�/<<��������#�w^�������5��=c��'�T��?.z��)�'�u�T�H淬O��)?�X�p���O��D�peYYk]�T�H��pKtj��"a���-F��h�����o�\���$E�����p��N't뾔�:u�����Ɇe����<Xu��ϣ���h�oDJR8Y��>��(�����m�KȜE����kӆ�����Gs�!!�)��}q�=����L2��9*�����h'�C��� �k�n���3(&�26��Mu:A,ǋ$K����˟�w�p|��O7E-C��x,7������d%B�W��+J��$2)'�%$�����:G���c����ש9Oŧ�		���""��8I��&|}	������:�:�D<&� ULV���]�ps��5xu{�65����R�����Ǐ7E|�ױ�<�}=?�n�c�.��?~+\`�aU��Wr�uY�8<N��iP�H��$H¬��;���&H�ʯJ�:���,���.ڐÅ�<�?�3���T�E��/T�BsV駓`�GD�1؊QB�C t8��T�<c`u�����鲦k�i����W_�gG�a���K*i<D,����`;���.�z^z�l�MWV��3pu|�t�����C�{�������n
��f��8f��H!�;̣ۙ_�M��:��}��J�����k��O'�rU����6z	K�^^��z¿'p�"��l,�^�R� �N�G~��E��s�fPVy9>�ŵ�iU�\�p-�;2������ں#�U���lr	EU��M~R&f�������-'�������V����ͮ"�|�����v�P����zLk����J�&�H{JM����2ޒb{��{��VY]�HHH���J88p���;,C۽�L'��H���Ņ�z`s"��c"3+��R#�l9�g���Or�󈊼p>\U�8m�{�~ _^,+�?�mʪ�P��,�[��X ��-���5���s���\�8��u�C~?��]���X�@�n�e���	��H����bM�����22��ǰ'\֮���KGG���L]��y�1#�e��t��VVҳ�}6�6��&���#�ͭn�=����L9=3�:���gZX�5088��v��I4�
����}7/�_}h/��-|K?ЋzzvK�hGG44Hr��1�5�T���>{4y�}o:)-����G�8��Z�
q}�#Ԑd�l����� \IGb�J���t�nGo���g@��1��V$�
�L�.��οy�<��r�����H���S*��x�����U���G��W��k��LN0���)M�`ac�R��4�F�]�ܚ�f��o�5��+���;>��X��_�`�_�%��x<犅�E�c�!$�%��>l#���G��|�V�F�߿ӓs^�W4^A�b��>"`��@W9��v�ω�Gz�\����5�qh�<a��k��.`�jC3�;~�[��Z�D�>���ĔOc/]�P������J��r��[Y+Ϲ�SZ��@2:/�>]0�OUJ6R����<���<)Z�{{UV-tw2�2I��okR?��ea\����%�^�!�����������i��h�&���`w�V����L�����v����3���&��o�]�4z����+����E��iƓ�rL���*�Y�a|a�~��c
��8�����uh\7�����9L]�@ʜQ�C�F�����n@�ӯne7S�Q�/j x;��LG v�MG�
[j7����K��S�i��]JE⟲d6�s8�e�Դ�3�a�	�#�0@	~��}�tqi)��t%���"cߟ.������N���o�ν�gmfƴ�&�ǧ���M�R��[8�c���Ңy��?)�v��@q�M�H����Y�ϴ�����<���H�u�_����z0��W��^�w)�RW�
�a`p��G<�(o�Ͱ:�d�����=�,��0 2�o9�����?� *�H�!	+<ȉ��N..�@4�L�k���t��n�������j��)*y�B���h�����f[d�(���ʽF�P��9��4�}_�\)�>sL�	���O�t�ds3�x�]`D�]6�[x��ߐ,���o_s���������77�r��忋�1����������)� 6�M���L=��m��s2{�A-й�`G V��.&&��0��L�v;̺:;9I<�*�JTT.#�<H�C9���g_)���h��Ա�{bVH�����`������7���iؤ�h��l�h�
��gH_��G�x�"�Z\��-��㡀o@{�S�O+>��#EB��J��$���%��ɯZş
�Xdru��a�y��R0)�G����LS�GQ����祝2��
 ۿ�Ț�o����U:-��"l�Z��K�Ԫ������ĂP�z{�&9���U� �g8��^�����n����3?���1%Ȏ�k���T���ò$���1�� 	��V���x3`A��ס�\�0nj���]_
�c�g�R>~�������"D����l�c�8�oZ���nJB����8���D�?�o��#7�#n]Pln�:��L���ޒ���+FX��L�#"�?��?Z��S>I>]>8�,څ�	L_�5���~�pņ(;�2�Vӣ&�@+*2J��:V�H/l�>�58��������7C5�|l���8��zc���D��qQ���|���/����E�����ɼ^�&<��0i�����e&"7�����{`�kHD�������aݫ^=��etF��5?x�d��vV���c��
A�0=�Fx��V~z�Q��*q����vo��hF}�+-�*M����ʖ9ϼ��}�x=U}�賈�N6-��//?��f*��k���f -C��795��&Q?���,��f�6�<X�n��.Q�3])Ȣ�3_E��/��x��/_�XVV̫w�%����I�s��K���&���LP)���N�x�y�,˹���Pn��Ryc�FTtN.1��{��qۀY��J-M��C���-��_X	=<=Mf�ҵ�Vb*�q:����[�/�n9?�d�}F���<NG�h��ae2>ckuub�6���)Q���?��5�Љ�S��^{���5[Ue�%�A��E4N&��n6�W�-К����;A��O�O� {X`�$H�D����q����T<���%��X���!�;>����rG�c�cs
~���/d�Z��<0��R��7����o'7�����ѱ���N�$�<���_2��#ظJ��z<����A�	@k�t��Z�b��ed}���S����ńVU^�R���Č���T�S���L]�CB$�yO�M�yz�6{�+�	!O�L�au�Uس&�m{�q�/k������LN7T��ӼCϼ�g�7��C�{|����$�E�&���/�6�xM���cx�+�D6�>隶uX:������#��<�;[\�隧�{B3��0����D�)��G�R��W��5�L�o��Ӿ�/���`Q�n� �/٠`a��q�m�@�|M`cz8�1n�b LJA!++���'E���jQx��N�����i�׊�?Eǁ�^�o��E�vqٝB�ɱ���T���MO�
���$�<�Q�����? o�� ��lc�h�1�GAC��M����F����@E�\+}��ܜ�A��k]�7������:R��9����Dk@��ɻ�]U'a����-��[C�*��ծ�����l#��|�V���9%���c��97����Zbu��z�z]:9��������bŽq|\���~R��u���#lr,�(��C@�4�Q��@� ìh�5�*�%}4՚��kuqÒ�o����v],,-_1��'�US�}�d���aF:Ǣ�=R���I����*u�qD�i�)����HT��~"#�Q+��� �WBvC,�D8����=v�'��?M��~(4��6+u�v�{L��F����l��C�[�E�}����4�-� ]J#%��CI+!J3tK�)� 3t9H7�w����{��g����}��{��9w,	z���������{Z�F�������\ hMM�g���8,��_�@NN>�<$|�[�p����Kr{�ތ��߿̴���y�ȷ����?>ʮ�A[��d|�s��]�& �u3��v`��߬!���WF��)���u&�?�BR�S��o��/F�X���ϗ~����A������ruq��,F>4DݏY#>�E�m����l0��N���C��ơ�<�&�s��
߁_��&y�P�o�J<���!���e���˛^��s4k�5$=�\2�>�ll�%^����8x�����@�+��孲2����}���Dd)$��	����E���������s������𛡹�.%���I�4��P��&��EߙJ���쪭u�lfw��߂�b�9N�]��[Uن��bxM=�ؕ�{@CI���?�2{ޝ�D�K���Ej�ő$ ��p|fK�<O��K_���8�>��)VgT<�ᴀ�Qd5�6�$4�l��b��D9 �1�ސW%�b@s�I�tnS(z�7T������LT�szҖ�*t�T@��vڌ�=ʣ�l���� [��~�����n �X%L�k�>��Ǌsq�H\�.�D8?Nūl�8R��8[�?���3��	��c->���5y��\9�7�ʙӭ��IW�u@�}ʺ.�� �iUU��e'��>���$����b8B��;���5$����_+��u��(��#�[?G���@���h�0&�m�E_t)n�廊I�D]w�4Geů���ƨo=<�B+�]�H#�1�D'ZmkCa���^8,��D�M,m@ɫ�{��:�k}.�}�?m��d�]�6�����|�հ��3<��dj�on��E�ft&R�.ܩ�w��:�Pm 5��Y�/�rC�l�j�	;[K��^<[�)O��_�)3̝����O�����;.9&�eL��dd^�s�9;�[�`�S����Vx-�@� �f��>��/+�\ϗ��������PL(u����Tp(	�P�D#*L~�G{<���շ��,�^��@�Ɔ��i��M��RE	��̛t��I� ��[���h8�Ԧ���ͥ�s����v�]����8ݶ5G�ϱ���<c���T����1�l&����Lo!ks�L��Ӽgu�ߨ&�RR��ɷ6����[���?��P7s�\��\���rgtz4�I��E(�&�����Í6�/��[W��}�X����z����-�?�"���̘�{���<h� �+�YЧ�)�����جM��_f�&�����"����su����(k7흁���5�i�Z�8]Í� �Z�`1\���fj1�n��D���}8����+�<���q����h��h}��9��oϹv�bkro	�Uw��n�\�,>�����U�#�Y;j�,��8�����kv٦���$����Y�����i�T�ǁ���9���^�������s��OO�ȁ!���[_��?�y���&|�f�u�m�4r��t?��?%�KiFi�)ji����}���a��C�9o����7�)�����t��i8���^�+����ogƌ�"+����m����6�-��W��8��!��H�[W���Ƅ��k����y0_�,��.����Υ�߂i�N�N��_�=I��N���g��x�kGFn.��G��=�������(���g��#�U��Ͽq��3s����Q0�Ԟ�~����.�}߼�$+eZ�򤢒 ��>���\���QW�(��5�����B�fO#�ѯ���&]ߊ5�9��Fi�P�E}<v"�z��3\����B�k���J3
�)S�����Z��E*,R���dȲ���v?I%��g��K�ou���X���VA+vӼT�L9���?�b���'!A�;_6�2Z�奏�>.sZ�L�;�3Q�T�^!eFf��h�"�i��^0����~N^���ԝO��B3ߵ���@��4"����]��.-�5}�6����>G̗6_����:�
ǳh����&eH�j�<���5�M�\N�����T�O�8.c��Ɔ�����I�&�)C �s(�L�󁝱�2��|���h�*�p?��4�%�o�<r�\�܈Q����%5��4�m�^���(�����Iq2�
�s�̴��###
yQf7Y�yh����0����!S$��fd���M�ƛ��v�3�@O������\,���P-��響M]!{�ſH�V�Q���E�3r���,�jlb���@>ʓ�`���65�������i����'�Cy��v�H�M���!����������WT�VF��-��y�}�=J��u��&W�6.!���%f�J���f�QPPP�ps�(K8���~>n;�&��Yf�"�m]�_���7A�=?�/�
K��Į�����	��%��	Pe�@�#iC	0�ڙe�����m���©i�8��f��͓J���}�_��Ԅ���!�qݖK�/ɥ�8�D�X�ȫk�'��m��S��u�^s�%��.���%�'�K�s�s���U��؞:⛲8B�@���������3��~���s����B;Z"q�X	�Ӷz��]�����諝���� � ��+H�br�^����Q4oO��":K�%�|�o��kY�c���]ݏIi�l���fl,�ߧ�E{2��ߟ�ٵC����U�I�"�o@&,�s%�LM��q⺦�b	�ͱ0]�ڪ{ ��W����׼�M�,�޹ JӉ�3��>>�꾛[Rߣ����D�����KG���Z��c��� h���ς*�k�07�w���,��G���!
!����=C}K9�0Ix���#sl2W�CT,7�07]o��x&��_e~7�#�#�Xqx��� �O�	퇼A�x��C	��*�ʢ����<���Y&YS?چ^L)�;{��?C�u��H �JM-���}�\�~�A�&���ˑ�k����񗍈��#��"�X\w�hJ:�/�}����꒞�/��(�H�C[������R�x�B}jH�� ��6ss��trrµe����/������7�m�l��x-.� _���BJa�In-�!+�33����|�N�4�}}}�������a�����~{���T*7�~�f;?�1U�Aݷ`�<�â\qo�q����;
����;v_MU�;wE(��@I�����>������Vݯ-�܄P�\P�}��S��uCc����������>�o2��0�.j�H��6N�iu�k��PMyy4^_<�N�rn9(2�z��:U�31yr��J��ح\��}��P�����=�΂p���Ĉ�~R/wC���]k�MLS��
0����ٺ�UB;0����X0V����� ��֫	��x�0�<{D�Q-�cu5�L��8�h�p%�È;���^s~II,UW2�L"PACGDD�\�3ti)Kau���S�A����e���@+�y&�,K�=��m�������_k������ƾ�X���-Qed���G���%ѩ��(,Y�<����{$U�q��:X���gj2#��j��.m>�!�un�z��ʊ��>�eq�xM����9�fc�n,�_��T�#�?!����X,Q��k��7�UF��˔�$��%����Q�Ғ�w|pljQ�"	���26��nK5�kT�g�p{�~��A0�I_TL�5��)0��`m�0�^*��K�h��9�f��
��M}0�6��(~���)�z�n��Bo�آP����:�H�3�WPP�h��?��aA����F'��-�������n@��ӗ�aI�Ӎ6�y4'Vz��P:Z��]
FN����&�� g?c��z<J*U53�D���$�Ǿi��F�]1����w��5�m�����>kDM<��Vvv����\����Hأ��uѕ�|J�J�|����[�S��'3 ���������un���Ŵ6���ݾyu5Q�><�(@�P|�W���S����� �z1HD�B�Rn������Iv_�M���`-��f��Z�7���a�>����Ҹ����^<� ��uYP���ۤ���M۳��X��S'ee=�gD�{�]�V��,�o��y���:=�5w$�v�j�`$0�y`u��4�\���ɋಁ��NI�3����dd�X%�Js%%�d��j�A�f'�J��<㽭�b�����r�&X�MO�z;��h08�bW���93�]V=����=|����-�ѩ��U����!��L��Ѱj�����Jn�h�j�
��S���5�Қֲ�2۝�O8� RME����u���DӜ�W��<yhQ
�߫����A�5������u���Eǿ)��^�:��1�;�h�%���8��;;6Y>�ӹ�J7�N蜍� ����"c������nH�B �zJ-�����ʙ�D��9�'��ƈe����nR�����~/?�H5�&W���1�((W$�2��pc����f���D���i����KZ�e\\\�P�����1��L}R�9���+�:C`�eT�� �-�E�b��>ꚓ�&�ZB	j^���%Xe�I>�d�ߘQP����>~xܦ�φTvIMDFe���r,{�p�>���
D(�p��o3Վ��ݏ���"���1u
N��椢��7*1�'�)SX�(��B�|���u���gM�� 	��ܗ����¢���J�ޤ��,"$��j�N�N!y��}"���Ç��&R�7M&]�&������-2��S��%]]�i��l|����&�o��iNz{�����������NII�_��k{~hc4o6]1�� �kw<��
vV�3�;����Ť�^����sfH �{IQ%e�js�z?�iw�hH�7���V��+R�\ A�>�����;Pia!5O0{v׺������SHH�Y�C����p���{��"��/�^��X����a� ��99��W\He��h��f}k;�_�|�pܣ2^6v��/.63:�����*7�򑱟l����� 0xND$�"�g�`7�d-33�X�."2� �8[�9�]�Ƭ�2q"��)=�P/i!6Oe�c�h��cB,44�����r[M�m��4x��eV9��0X/Ǫ��s7�n�Eז\��L�B�����3����jj���M;hf�JEO�gPppLll���̬��D*��_�ѕ'�9kNM�3�Y�(�/�A�� �jc�d��`�?kw���X�=A���Z����ن�lD��ۥ��f���m��[��Z?��(l�ث�R����ԔF6��d��JiZ�+c�t���9� ܞ��4���(��
�P�E'rq�3<Gv���\���Ż���կ3�!�㠉56�]����-�*��2� ��r�*��f]�H��,~z��sx�:"5��k��ōI-Q3]�#�g���r�ځ��TS� 
�>�����&�W�'"�5/���v�1�̮����q@��\��`��$�E��K��[�(JIJ��9����� �[r�!Hk�0kx���h�?c�p����+����'=j�0�ag]"Wߠ0��x?�����ۋi�ǀcf��a������,�:[jɈ�?� O�����)l�������!�IC}�eU�*	�-��1��Yd��V2v����r	!i����7�F����Y,������r��cm�1c>}J�5,����R���ӕ%�1����R5�ç����ݯ$/�h�yy�+�Fc��w ��O*�H�%���� �8=�DG�~�ݖzg���?1�.d�.!Ϣ},I	�(!�p�H��Dg�<���ӽe��=�o�k����
GTk��x��~<�}� ai�j�t�p�
�����.Nb�"�Ζ����Ӻ�<zM+**�eT�1�U~���?T[�a� ���� ggt�Qf���K@����mj�r�D��<-"#l�X(����x�����f���9��~J>8b&�?~�;I o G ���w97@���>�Np�+��&k�Iu��.��7�6v�O�����O�3�4��z� ��������^oO�IHt����)Ni	�d��b������)�R�>{=�%�{�ġi��n�/������$!�j.�lk�� +�ߟy0�O#@a�z� /���ms�՛Z(���#:�j(�V���l��AD���{��մ?�]�K�v�a��1~�!�q�іSWd���D��3����%(d%����^>��v�����J�c��x��tE�g<& v�4±䠵%���Z\J
��`Ҽj\�$i�!�-]�!�y|���� N��@xxxbRb���i���`�� �bҪ�����nhH�:T_@؟g�Q��?�\���~9��B�����;h~i��ͅz�QC�v���_�������i��h2����q�e�mr����euu���y�Y_�}ds���-j\ i��*�4Uk����6������nf�%��Ĭ��<w�Ҭ���J ����m�h�������,��{��պ�h�V�3jd�v�gR����Օ�̣$H��I�3�KSD}�~wS�EbF4��h�?_t\�� �磕p������kh�I_<3��za��uo�I�?ѧ�{��"�	IfN�)پ��MMM�N�:8�&K��AaSeFLzMa�b_������ª\�HA�{ey���������@f}�:�т����N�$++KZ��mG���)�����#�;�q��F{m�aY�:@��@�߾�g����aL麩�Б��4���x[��)��B�w1{��s��$�s�t��/z�A�E�oE���k��<f7Y�s۝H�`9��M�_ژ����Lh���P�Gޢ 2L��T�;R�b��1��k��?~\A��ze�^�Y��N���tK/��=�B�r��8d�

K�߭=8-z��#-K�?P�ڷ� ��cfV�9�1��"�G����f��[�z{�gVp�K`%�:`/����̳�H�� ����o]���6^�c,¿%�9"y��kaʖ{�G}�ۇG��C�]7WH�zg?�(8ӺaGmpd?���"�/���I��-�{s�H����j��^�!@����WTt}� ddm��UGl��)��"�����z4��|md��� ��LJ��b+KKÅ����m���u{ۖ����9> g��ق%�A�A���lv3oXH�}�y�M�S��_�#汧���l�J�#�:|kL�I�LG����5�a��\I�o5�C�
���d������]��ze�5�Ch�!jm�L�4�p��t��&����y�����w� ��Sb��"|�Q	]���'~�SH�*-e�"ڀ7e�f�zR8�ݑqsJ���Q��d���pG��X:-f�A�^!��A�-HM��GǤ�M��z��YL�&�
뵔�tʊ<�/�ِjC�A�S�a�����|�m��a���Z����\ua��C­�88IVv6�y�u5�ϹK�C���ЅU-�`�~��?�*7��2���7*v��fq�jt
bBo1�Nh��"9�MY�W���|��<N:�~p�{%A��ђ��* �^<1��L��x%F��)��K���a��,�`�Z��m��.�|�� Ӟ�9�|Q�$/	֜��n�I�ش���������Z�	���КpN5���*�A aʎt��SN˚c�o
q����g��S��U�v;�g�� �W�V�̷5?#��'DB"�WJJ�q�}τ.��ԝ���x�w�|pnS�������~gxV8&�5�O*��.
<�/�$K��6���� e�M��}�����?D��/
6����� 4]cZ+*.^��"&n?A�
�"���,k ���z�և��gԤA�C�ƃ9+9�*][߾~5�Y�$�;i�i>����@k����w��;n��D��Ԓa�t�
������,�E�l�vJ^.q�>ݫ `���qr�v5e�6���kĝ�8����ʘ �%������<:5�D2�D���4e��1|1 �(��w�YYt���_TJ^��VR.���+)�I�Ø��V���F�+=1�sUI��� Q�%���$]8����0gB�Ϛ�DIt��5�����B2	��PX��ݻ������lR2�A@�#.�|�0�ݜ^�{�ϣ����@��	�	
���|ך�%���� ���%,����A0��ۋIS����0V#8M�,�%W�߯h�ס[�柝٭�G�޼ys�ڽ3B�r�.G�ܐ0B��U�Te������Rd>�ŚS��K����G	���C>�@�$CR_cROY��5�I�n�+h{�)����;��3��6D��(Yy"[���1���5��a��)�3�����B�X+u$Rx�����# �^�sr�$k(r0X�f� Ar�Ŷ`/s2�#5`�,�n*�s���O}����md�5�#�|����&di{�f�m�{�v�w�_�6��/̈́p���v�.���7ɋ������I�NMEq�ջ����.|��;�:�'#7���Z��#��S<�ʮS&����73�0�G^V���N�P� �Ѓ�8�_QQQj�i-U�GO =����:xai��p��
|�H��T�0���)T�[z�N���I��ӫo�b���䑑���ҋuQ�R���TYEeT����:Z^���.��K8�]���WW;�GK;˜OfO��䩛&&���Q���n����}[�!  P�U��Q�_���uqqq��Ɖ�����-GԹ��"=�q��&�5Q�69\��	���OZI}�S�?�]/bih�ڽ�&̈́8��o�Fj��h� �R���э��6޼��B� b�e�d�|"�@����@aAo<��nI��W�>����`�M>��JŜ*�r���Y�lȢ�� �g��f��������Ȥ"Iv~t��6&���kO�L��o��?�v8;;���^6���6;#J�S�nS8��	jaT�
|�O�}���I����C6�0��S�o�!��-�Y�tp�z�M_Zf���T�;+ǚ
�c?�!�m"�IS$y
���i^�5���}z���-��ȸ��[[;, ��R\��QFAfX/��1����W,,���V�B.���*�<���@�z���׻W�B��PQ���QdF�����2�K�	g�>DU]�M�D����M��S�P�aƎ|�Y�G���]�.�K�� ៥���u/��e�q��?$��������܉ ���\����aZ&Љb&\��_�>�Χ������eނ����U��?���~S涣}����(##3l�p�G͜V������cW�A��0��P
4Y����k\9�K�܁���Pc���6���_D��r�,_4g���'ge���G���U�ǿ�?�?�n�$em�*��*bH��xX��,�ʽ���|�Β��ם�e�q��z�[GH�KU�Ϯ��i�,�d��=NN��:��K@�(������-� 1���阵z�)wu��
pL��d٥��A��.wޯ(�w�}\�����|=�yG��Ԧ�}P����m:É���g�pq��:�_V��WJ�fm/;;f>>"N�0{g�aT{X�9P���f/�1�����90�&cf5v�'
zp�{� k�I%����@.��&��j�D�S�K�:]c��㓞z/��ЍR���]Z���sk�c����R�h�� �Ƕ�	��.��km�1c!Tr�W�N�V]�A-����9] Rv���_n8 mӜ �l�� Rt�F'������bk��i�H�� �f�`6bح�x���+�)L�A��s� e�E|p� ��񔊼TVl�5��խ�"u�Nm��@�燨Ҳ��EE�TۄW�@I^�W��!�'�#-��� �u"����~T�A�_�+��L�W7,���B��@
<�?��T9��X{BJ9N�<��� mSH�t�p�J^T��$����K��PAA�&��}����u~I�����an�����5�P�}���P☋�5A��Ky�Z:�'r�f�B�>~w� �&��&Y�׾��s��h��sr�_]�p��M�/���np�~���f`*�x�<D��������bğ(D4�~��|w�`�F	y��O /a��	������-1�/
o�z6I ���OCwxC��<{��|�Q��݉���M-�<�`�wZ�UP��1���08k��J�|����Q{{###Lr�����8�t��!���2�+@j���\��D�7Y/ܥ��
��KH���_[)++?
97�튡�<'��4Bh9�2z�p��Lm�Ti1t�lJ0:�*�B�Mq�-�1���fXcJ]�6�b҈��2q@*���Xc>�2�O�6Xt�T/)�#W���cl�~+�q��V��'I�|���naT#�O��W8���<vW�q�"�j�����J�Y����;Ѭ�,�o��QdH1�>�F&��m2���GMM�v?�"��y�?�G���
��w����Z��?qtA�F(Mkk� gڳHG�*\499Y��%���*�s��v���Um/i����w�&�]�5S�����A��k�+���ԨMG^ͣ	���9/d<0݆� ��T�ed����I�ӯ���׵�������!��}��m.v���������n�U��ycm�₻��^�}lF�J��a�� �NWdLl�H���j)0Ď��Ё��%�U�S��3$@{@�\	em��� [�d]�����]r�ς��Ε�PS�n7��B"�t_�
X�M˓��V��#E��ݾZ���Z˺�_��ඖ���y?[����+N��a���90���;w+�z�"�9�.\�e-B����z��>��<��V�)��bzLj�̯�D�;�R���^0���zԻ��!�@�bg����3��zq9*+g��Dn���� ʉU�w����7�S�( ]�
Y�� ��qh�1�>�X����-{v">���<�?��:QVW���!�镃o�Ȣ�^ܺA�+3	�-���8D�m(]�_����?�ho ���GmAء��,�:YS�����{4�v����܇���R�lO��r�S�z+#�	��nGOI-������ǫ���~�o�Ó0����K�#M-�w���s��Ðξ���3�c|�z��Whooo��Q�R��;9���6��(���_1��.=���
����=��쥧G���A��Z������w�h�5Xb�������gR�~v���q���\c���\-��5��|�:�a:���}}�LLaF;+��T�#�>�>�Yk+��	p�-&���+��s455�u��^�6v��RxC1��h·�_�`4�=dџƃ���P^�ayIm~��������{��7,�X���p�3B~��{g.�;~0�;���b����>�:]�۶�:�/j:bVn��: |��������醤�"�E��Ǥ�H���)0���P'�׌��l��)�H�f�� ioK�:H6?op���W�\9
����çtDx/����y�'��z�xtmm��&�~U�<�~z��f�1P.�KZ�`��iJ�{��J�*y�v�@&b�}	��<��	Y�]� A9U�m����u>Gp� ��z|k��'(����T�.U����N����I���#�} �))[��(�>V��<�7=zJ�ܵ�F��4S3s�Z?�����=��U8�J���-���$���̌�)��J��2�-������2��H�m�p�j#��(��z�d4F���ͰN`�p���Q�W���1�ߙ��&U����rw���ٙ��f��cYST�\���Qה�
Y��W�gF���y�������VI}��O�3v�i�������/�|�� �I��QiI��՟�X;��$�\�9���!AH�0]�_t�{w�����t:%�LE۠�|� �)(P��L���F��0l�^�-%�8���J�m �������'�>Tl+���*k[�3��v�4����W
�Vw��	�a��߾�ƃ##|��e��u��mr �>���w�*;�'��6��>tvX�v� ���;PŖ� ����������� ����'+wrb9 �����0F�%Y۬o���ԁZ�5$����}�54���6�ܖq}ڥ�n,p	�ĳ���C(��&�����ڮ�m����hK9�|�uq����>���% T���U���|�k#!�B�mKĖ�����p6���sr�]����"!������jq"7CW��.�t�2R��d�]��?m~-��h1?�� �y������_�~Muf����l�������%�x����_�NNL�Ӓ:�RP$����{���������8�~E����"�y䞶�ړ'�c�Jp�f$�BC�������0ߞ���zx𡠠������ f� �8Z��
��²^�%��h��$\N���9��**b��d��a�K@ :��2���#�s��t[����YF�hXK�����9��P��`�5�>���|:���)I[ML�= �v��h�������~�@<0����h��� H��D�3���$
��٪9ښ�N��O[�i-gB G�CP���m����{�$�')wD��}F��j�j�<�^4"1늤��=��ha��w��͞W��.��ڛ6����Vg��[��PW���\ZZF�R�|{��ξ�:=R��e�О 	yt�f�(^��Y #&Ќ_�������7�,�����K�)��< %F?4�B�=U��Z�E����<���9���B����������a� vX~�Jx��'***+�?�|,�M��U� ��썄��F����K�eߔ������-@��!7��{�c��4�
��ߡ�֮�`d�M���o����!����67l33���N+�/�3=����{���U n�xI����g�%�4�;�ZR�Z�	��������qS��G�pwխ፹u_R���Hy�md�
ZY+K��/���o��h���陙��H�&�<�m���r�)�r�Rtq�k���8O!�`3��_16d��p���a�m��}�oFJ�"�������F&�I������������L1����<Gr"�����d�{�<ݚ�4{�z;���K���g�=}:���9r�f�b�R5��b0���~��`���]�TOO�z~z�|��v�c1�<������ifΔV���u���O}&��	��G�<�k�*'Y|V�k��*w���&]��TUx���Q&Z��Kvi�P��[ ��4y�]�o�
��?Y�bݻcwf��6y͒��[�w`o�L�3���R.�0_�#�׊7�I�D&1s��l&kr�.	�|�Hž9�N2��6��Q��9TRNSXXx{��)%��֠�N+�*s�9��O42��\1@c�S��R��������VBS4h�ipc�	�Ȝ5w������)5Mi=��������Ղ4n&Z��	M�I((�>MM�r�����U^;�;pȱ���eP�{NSr�|}(��K}����Xi��E㗦e����8�ց	����L/lܻ���\�����8�B�f�i�X��+����=�y����h��*�zu���S~A����n��ay{��v�s�3�����&[q��v9:,�.��P����M���L�q�������K̟?�K�'�	�Z���L�s�9p�� ��Ɠ��w���1UW$ivE��˫\�Z�um��Z�_iմm��<-�TC�m�N	���٠C2C)v�X$)Oėsϐ�����_����y���'q�pB�����x���G�o7�(
��N�]�=<�	��o��m�s|�A%W���Jԅ�x;�"�b�Rw���#W	?��^���'33����u	��/U�BkՌ7al�+yl1ٺ��>��
,".�����;��0�]����c���Zb���_�`�/_�bd�!��P[��2�2}��C�R� p���ڪ���L��*��!c���w۟��$���KB"��B��7d_?~�վ�DZ��	pY�������K�M$=T����!dYY�W';��́(%7 >x#ɐZ�Ѷ�C�tf;̦L�<������NGʻ��/�s,p���H*F��\��V�&	�c����3Kj�Lr �#4�m@�� �9�婓�/f���͕t~W�<�_��(\�¾�a�<�� �~�"����
�H����r���yV�|.�i ��=k�'Ӑa�&�和�I �zN�"��+��R�G��,v�Ywl����Ʌ�D<c8T/��;e@<|����ȳ�Rו<$��o~�狭���!M�,�&s�'���I�,;x��+N���S��3G.����� m!;�������Php�\�`�EBB����p���� �$60�Ft$�ӟ�U�Ľ�̓+�%I��i�^c�n2�������# ~��ܽ�w�;c�����=|1y�^���h:���h���&�-���q��M,�3����t���3r\z��K`�����y�C6Zw��W�+@���"��Zd�u�M��]�,�?����f/����FC���h�s�*.�T�c��Kx�ɦil[%���0!�Z2�k�
���{�D�E�P�H
���{�t�O]�������~2e}��\��^&�v\H[��ޒΨ�Y��A�E���M�.���;��KW�mc��LȦ��2=����3����u �00���"َ;h��d��1r���۞���2a��@?xwe�H~�4�?q��>����$h��:��������i)6��f�j�ouR�����.��/_n�W��(����$�|��T��+��g�O}%i|?���ԩ��xH%����}������w,�������߄��Ne}(~�d��VTYG������n�A~��n�����Wa�Cz�-svX�������GD!�x߬���]~�zR���s��8���o5׼}��W��׺�	L?�۔�%3��ŪOr`�9��mɬ�c�t^It|�BiS`��K�����JW��3_Ҽj}�.qT��QT�Rq��YO猡���첣Z9p!;ѷOP���Nr���5u6G��Ε�ᩡH��%h�~Κ���j��ӳ$i�\q�~6�@b�[��[@K�қ9DUK�E.e�8�v*O�^��M�L,IE�o���r������Z��?��4c����=
Шч������$�Y�SE�l_5e+�HfyJ}�:��z
�y��MB���l�،�
�����b��dT��Mu�՜�?�O���m��Xn[w8�[�����);����CB�z�MBz�Ǎ!�R��;o9_	8[��۲JY�HZ���
�r*��;�����H����W����=�H��wG�	bU����յl�o��^��X��Z��x� �3����=F�Ѹ��Ϡ�&�@3E��3�^�l�B̞�q���)Ҳ�Y���"�(r�Y�/_0t3b~��䛄��̜�� ��O������:
�rč)�c�~�~�yA�+0�c�-'��7(|.BU��gO ʣJ:��
�=�7�	��٩`-���%��aYA��?6R��x���V�����rz9�T�=;�Bv?�c���x��/YvHH����k�St.,���}B����a�G!J?UgYů3�_|?�Y�������S7���CA�o���-\g8�L��/�?	���΅��<�9���X�����=�t!�׭�b�"��hSNa�͞��ZJ�j����R^E�4������?�_��ؠ~�	ѭ%=��]a�3�ښuQ���f|=ğ��B����#��+Gr��oX������cBeТoZ����O���`[W�`�"�{QW�)��Y�0lAZ��!'j���r���� �$
f�c�Q]���a����|�N٦F@8`ў�$��1t�2�������},��x��&:9ԓ_.��2=7BgLz\k�F���B�ޱz�̙�QP}�}��W�wG���RE�_�aD�Mv:�zD,�v&y�x��p��YC�`��H�lԵ���g�kc�����e]�.A4-C����TAm��K�v��+a���Z҅�>�:t���;d_���8�3��\J��U2|���W���j�k6�>c{3��3�s���ߋ5_9g��t?��#f�\'�'aQ�>��X;T�%���-����_+��9�@��)h@�h����Ňs���:��_�>,�~*����ֱ�Mt�w��Tɼ���}aU�C�&�~�&�����C) z�{)�؂"覓_J��K?Y�<��n�+<�JV��nN-Ϝ#6t��"��O������~ې��k��p��5�I{܉u:���������_�I�~*a�٧a��E\lG��Ov��n�(׿��a�-���)�(�`��iqNg��7¡���}���x@t���˛`������It�"����C�=���i��g���-tey���!�.O#~�~��Civ����l�A���5lrԨN�0m��]2*�nv��]u�c�6,8��p W��?�
�NV4�K	��& ����@ڊ*�s3�bаN�wXy��۽RG�w�>��6%�!��@?=%�����6E$LJ��s7�ps��'�P3ܛ��#�'
H�������κ�̓�;x�8�G�����ߕ��ޕ-{��S�Rs<F�s\�}7`e}-����y�]�����9�e�2�ݼT���q��sx�ﮗ��pd�NV�J��Eo�{�&xo���ܧ�Yp���]&C��:�u,��~�y���$N�?`���뷀c�\�n�}َ`Q����Eb�z]��_�D,ظ�R���>\.+].G���.���c͙r�P����g�ν2�uҟM��n��<l
2�= �
-W�V�LN�s&u�x���9a�`�Y�'���[V�i�Cv5���r�w��t*��ldMFE9<�Z�+��)ص$y�+��5��p�P*��D��D>��,�屋s�u_�I:tk^�G��2�
�t�'-�#�(3�}<�{�_p���N�a^d#ᣗL㜏�Qv����Gt�
$j2)H��F�y�Ȯ�Gmոx��RN�5��4]TT�Ӧ�[��[��E��nX@B���s��k��NAr���k������s���}ߙg��y��g}�$��	�w<;�z��l�j̆���[x&�P���q�"h�Q�lV�-���i��zD�� �8�TD�~>3-J�N$���=���ر1)���A�$�SX ��˿�$���-6���@���e`Չ�l�_GI�L
p�)�+y���-C�
3Ņ<��.�����m���Jmp/-8K��m��~ȧ��aL�X����sH�؋�m���P�
��p�oLw&[�2�`��);'儓H}OB[
�ے�/G+��&tXc����d���ݹ�Bf٨|�C&M-;��ь4V׾�A��%Z[_��A�B�0��r�gf��b��݁�u��c��[޴�@�%ɡO���E>
��ʝ��j��I��PTC�>�oAR�		��ێ�����[È����(|��Zq|��Mz�~��?�՞�fм�U��"c���۟��)N(��_,h��cP��r�?�d�m���PӅ����q����=�a�^;��P#�̚7[YֵھW�`�8�]�h֊��p��վė���j�9%���N�|sZ2,���@�'��\�������n�����<��Q�+�D��;�7��$}�a;B�)�:ԡ�1��ykn?_N�A5���x��利gE)�>h��D2�P6;4�\�(�f6�����S�^r5!>-	 ������;�����P�'lb)�w`�������oú9��4��I,Do���K�D���t����ۂ�s�9�O<؂��+�\g��xl�Ɣ���#�Ka�-�^��Q^8/{��X�!;y�}�H��蹵��702"��]��^6�1ّ)Ϸ�h��1H�0�P��-�9n���PY��O�B�؆��U��|؏{-8�K�S�IYe��#���=5m�C�r�/��k~�Z�+Yi̦`����q��b�K6�ŏ�JnR�y�<�e����;�Z���R�T�*~�btn�:P��B�ō��`'CU�fJUu�Q��Y`y���0�H <B�-$C{9d��*���9�:����zU�(�_��j1�'O�0�����ե�+FOB2�b����o*����&Q����n��sL��c����7��C���8Em@ꦫ���#��H��.yd�%Cj%�R$��F����J�qg�%! �j��-��7�	=����(OC/_���b�`Q���W���߮$3�A�1P0+ի|�S�FW�L�xx��*�|$�"Z�,ZhC���	��C�%���y}�d'����-W������`-���R�6-Q��
9�{�:��	9����/������U�W}
��A{�H�5�]����#�|Y�%K[���(ӂ;����2)�|����2��$��Z�U [�_�" 匟<�v3�������^!�	t�Gx��8<L�D�}6��'�n�GC��������C|�0��|!��n'>��,ݵ�7��ѨY#������[j _��H�p�����Ve>�������0}�2A�({�_n]�(|��l�W���Nq�Z����t�7򃏧�æ���[�#��<{�I�t���S���J�z��_d�0��o�f����e��,�}?�+b�%&z����O�Qr�$��j��^�m�-)a:5�֩�%ke�G3:m��^���&GLsA	��0��~�rg3#}du】䴧����L�i���̘��Z���+��Y_vJKҏ�n���BD�Y0B���>��;��<���0'��AL���`�jN(��V������jO�?x
,�]0���������7��(��9U�i����'�s5?|fС*��Þ�������9.�5�=���^ujF��.�ӏd<l� �u2����'cIai����K	�˦�N�F��w"�����L�ʃ`��`����D�e�~ZC��W�`�IE��f������Z֫�~�7RG�R�)�L'n���f'�&h���s�%灑�u��x�Z�*웭+D�i�ƓP���\t���u5s5H�M��O���ػ_&�NW�5����O{��A��8?��K�s��ܲ8�"�!PT]��A_s?*��3u������P����ͯء��Q-a�����& /Џ:���s�ܮp��<���^������	^���"������,��c��s��vۤ���|�o^�E8�m�@b�|���j��>��8P�)b���ڨ�uk��1g:��nJ�-�L.�����m4@X]t�t����[Q���:���� P��~*Ȳ���O�o;�W�K]�V\ۮE7��n���( ���Q�:��S�k�ж���X�ʠھ��/�����(U�Gu�-�Z|�ߗF^X�'-f/g�������O.O|�,� x�����˲����tx�߰)���L_��Ը�<wG<�"p?}Q#@�C�l|�%hzg�Ӥ�v�7�����N����C���Mg69O�V7�o�����ȳ��4��8���k��hG��6�&�LH��D Su����=�F7���r���M*M���68v�TX��R��H�xZ�P����Qp�.�LG��1��� ��p�ì�?X��@�`�6Q�0Q�8Ii5���ȋ����-�En؎7&<_�`��u����1��Ca�Bm�h���[׹g���Q������Q��(_�o6 �mP�\bP1;eN~�c�#���d�w�s��_fV�J�6����[�ᦽֺm�*r03tϮ"j]��v�)�3jM��w��;�����)������P�*dؙd��-��  ��޸�7��\[9e�Z����;��%�d��I��ΕN��!�
�+P}��ƿ�s��ac��?�i���9���u��%w��C:�$�H��K��WK��	T�B:�bG�y�S��9��C_������~�*�{��=N���\�,T_��4��bG��)<��y�	�ge�'d�sf�gi��1���κvp'�WG:�(^Q��nۥ���8u���#ԁ�O� �R��;0&�X��2�!itüx@{�ite3�l�#%s����Ȱ��Q5��K.�94���h"vq��!scۆ�?�����(�����p2��D��i�"B�8�X�M���ػ�k����(�����\�G��L5�A����r,ύHD���T�{�MצB0��Ӯ{�����Jg�����zя���%$���L6;��p"�ruhx�x=�z4@�Jn�e�g�E�`m��_�o��b��L����9�?���C?-�Q�L�J�r����8��hŎ3}��"�dNi#�B�|��Ť.���l����`p�|�������Xg��n�#�|9�����2֢&��c�1��Z�,�?�Q(��-��ٳ����ܱt��ׯdN�q��[����K��������x����m��o��DH��)К��q�}{�\~�}�O5)T%v���烋,i�*qb{ͦ��VOD\Ju��k4B��=m�
�$��oj��*��<�k"x�M9���~@�<o�\>c�,��X���͠�E�/���Ƚ�ݘ�Psם�����g���C�xG��fsh��
ѥ��ޓ����D��i��H��"�G0~����IOL�������T�j22I��T��j?c�����$��p�H��r�A.�D�r(c�
��ӯ��b#I��=3Sx�vH��jB���*6��y� Nt6���UeI��[/�G=i{���bzumG(����t-�,a���gAhll��j� :US���K eR	LϞ�}��N���R���m��W���K�\�w���J6\�O-��ld�%:���N ���dIKm��^ r a���x�,Hy]�<��=W���Te�>-N<9C�&tv�*$��N#\�,`^\ZU�&D����� �>��H&C#_kGњ/�ueӥ�XyRE_�M�� ��Zǣ��j�S���>{8�+GU07���w�1��it��Te�����<�U�vF6���QxO�@�!5�M�[9F)�W_������mg1l�� ��2�7�X�z�n;��@t�le-�=8�baa!ۼ��:�?2IOI��=�\	S�ũ[KhE�:z��٘���2���R�nOo/JL_��~+���W�(A�/pw��W����8vQb�����S��w�] O>>��:���������`/,,X/��������x�KU�%j���mK��D���q۟��.h[89��^����ë�Vւ�НW�G��}ۏ-]]����c3�	�<�_�/-e� ]�>�7m�gK���&@����������h>3�%�|S�(Y�����S/��ΣwN}�����1�ww?����(�]�p\�`���-��8R{��`F�Q�G �����v�{�(�R����m�����x���'����r����J ���/��+B��gmW�B�o+�;��-\N�|�K{)�E�)��8�b��j &# }��jj����7T��fwӗn'��T!� ���;��n��r\�/���wq��m��^�ڙ	��Y���`b�N:o^��t�#��}��7� #+���⢠�}ݛ����OT�����v�\exV��$��|#��G.�1T?��V����B���r<'
Y���fiBo9Y���-99�s� �=8Y��y	�l����y#��t
�������苭�
��7��=ϧ��l�2F�/��U�!ɟ����{إ����� S�h��5H�E� ��g�(��b�W�9p*���+��$C��ͦ��?E]�_�)���K����>�c���{�.�ʳn�N�g�	*n�oLy�7�2��ddd�TƧ��ӣ�u��&@�I=�L��>���o
<sc��d��K���
������x�<��S�&�m���<��~1a�����f��CMʟ`�!�\��mh��	��� @-z޼'j����rӚ����3Q�m�=):��Iݛ7*ߣ}WCHם�H:�䤍��]^��O�N�~6��U�Zw���~K���X2W.�H��3��4#.�����ľ���`tÁ�x�tS�VFr������S�ɤB;!��D�D.s*0���e��y_J_O��z��c��F ������7]X�ptl�9�U5��. z�����b���-+��1�J���B�37I>�<����_��g����M�ŭ�7�sBQ�s�W�V�bg^�0�'Hk��7�l����͊N�UWp�߷�����p\�XdW.��M4��*�dN_��������w+2&4�5�X�+.v��n���^���XR����^q�D�0z���S�	��]�jo�7�2������/��ۧ`eJFf&�G+�����fw�}\�Ͳq���hoϑ�ٮ���*8��`�?��]]�8F͝ӣd>R���d��&z�&��&#x�a;q���xl|<�k��t@�E��k�튾I�^�oC�H�O����Z}��V��=SH�U��gzn�Xn�*�H���J������i0��?������9CB��<ʌ�2��'���]Ǧ�q9*a�O|'YG8Q���4$|���<�n��t�&R�fltt�� �Ǻ���?����$�k�F;Dk�w%�K��xuro��<+l��B��}/�fc�*�^�7XI���4*q��|`U+i�	T[v-x�O��h�4HU��&(.N�<]���4=� 3q�6L���q4����W���B�dz=��.*�:�<�Q������V=�T9�aX�kS��Da�g��h$����־݂2n���]�W�wzMC��Ԁ�XԪW�#��_6���?n5��,�5Q'���z���d(���m8�bW��l��OUk����"��:����]������Zx��|:�F�׵ϸ$]^��V�Ҭ�]���?�O�bn?�WDVN'}��Q���p/^
81��qj�j��>�B�rdzX͝���0m�?)�gǒ��3� �W�F��/�&I����%�E��h��p��ld8�����\l�6�����*#����L�4��	?#;{�l��j���;x�L��Z�u�/��^��gix^z�!����EEK S�������1n�U��7B�_����0ږm7���R|T��7a��z@x����%Z��(,B*���9W�.�d��/�+�m麑���Ҩ�YF��s��D)�D/��	̄z��͙ �%oD�~�~�B��aa��RR���Lĳ���* �>�̊�j �0�w����!�����;�&�)�t�����¨MO��m��r�-}�|�EhZ�C]��T����t��n�}�����~�j
�Q�@JZ�rr���������i�)>��	�� ��C���뻻�ȧ#ʢE��k�ޟ�̨s���rݴU�������+|X<`�2���W��F���Ȼ̘���5�k�o��O)S�����8�����+����R����L(�'�8\�\�sC��A��D�Tȶ7��-���UR��k�/��qE6,�[�����;���td��К�M�w��a�N�q`��=!%4dF��'��I�\��D��k�KC��pAm�	�N0�
���r���IQ�ׅ�Z��lR���7/�=i�%S���Vʎ�K�yz
L��c�٤m���
V���oE�ל��N�4��x��L$X�������dB�l�8a�k�0�:b����i`����VaI<"��d�1��!�3��Ƌ0��`/Za¤r	|WZ7z��AP� ��k���q���������'i�Y�B%dv-�^����5?�ͺv{w2A�m�����gM#�V�]Z�!�Z����@����$�����)ôP5o����N���X&���'��L{jI������8���`:C�
\�Bx �]f_W�U�C�q�P�EIҥ[S��>���+x���>؆��^��D�%3��T6�������"�LB;xpP����6*��PA��;��ቦ�2�y�|^�o����F�:ڞ�X/�<��Ѣ�!N��$�InE�p-=�	�}��6�+��f�d�;WV[�C��֛%^m��[���}B���y�n=�؃@�}ûR�?B\5����ִ��s������J�eM�A�ދ�= ��Ή����������q*�MG�vQ��W٣��e�`3,~�l�S�џC��%���_l%6nExb�����v*_ٮO���/�7�R11�q>}y� �(�0�.�����Z��(���_m�+�G6���H�/HUYL��iAXrЖ"�Yg�F���E�����&��7�v��B
:����r��R��V$��y�r0��Ɨ�}����E�
��a\�L��^��:��_P��X��˯��}��[Y2�W*L�.��F���<��VS[�T)�~� �/�f�� r��Ɲ�T��te��׵�)�(̘�+�䐡�O�8	����)L����Cz�`,P����)�F�/��7�������3s��,�����&g�� �V47�Ma1�E�i�B���m{{Ԡ�MB�^�:��4���]�Jrc��{یZ|C˴}"@��'��%���EX�~m�PaduNo�DL����3U�j�����!3
���7A��ږ�%�L	�Zo��i����ƕ3�I�i�o�~�����XĎ��^Ǩ¤�P;��A�i����A!CD����D�6��`�� ��&*BB���IP�F�_�eR�n��9�[�\2w����������.��,����MFͯ��^O�j�=�ɅL�M�4zEH�|����!ʪN&-
sK�*ˍ����k2�{7��h�<5I�cʛ�")��d��x��%�0�U�Wb�w�u��A���a��_�:T -ӯ�#�����#�c��G���@�B1�mY���1&�E��Z�z����2'�U� h���̯&2��B+UrA�*�����Ҟ�b����XRB	��'x��k�%���9�+��*�f���F�����;ftKR�7�b���'�DVɖ﬉�^'@���e[����hװK�wQ����W[2Ex�~<a�ƣ��>��̭UCdm�������]��G�.y����Ƽ-�����թ���Y���N���y��t`��`*a�0�c��
<Y+��6ֺ$F����߿l������a��=���Y��q�p�q�+-�r7�|�`�Ӽm��Y���7�=<^=��A�&����#>R�B�"7���"U�/�0�$�G�)5��hYK��@!Fڒ����ѕ�x���﨟��*uN���L���㽼��OO-j�|����Ќ�%(�� ƚ �ȬD� �>P?}NܰӓM�$ ��%���E�����E�+�ޗ���C��0��!] ����.�(d��hXNmv�F�\qc�3��h-�ַ[
b�Wx�:������O7�V�,�,5o��>����/���$�=?�����K�j��)��}��:�4�fqd�p~,͹KV�sbf�zG����)�Y������?�`��� ��PM?r-VR�z�%��/5��B��Vn�H��e�^Q��?�^ �Y�����;ȧM���I{c;�k=
�ڤ�U]��0t>�a���B��on��N�7��͇��F�~C }j7!@ �*k�B�V4&zT���oE����?�Z@%���̮<����?Z.�� ur�i~�q�i�d�љ!N7��^�RQF��>6��%�i�cN-w���d� ������ϭh�#�Ro��=�͘��^-7��]���Ҥ���E��ZJe*ޒ<�k]��9iu�z�8�޿VdD\��ή��U���aWZ���C��A�;�,��_�-20�A� ˘��	�>9󣠕��I�%L�c-���6쌸~���d�l��jL4`'�{��w�QL~�,)$�?OC��͵p�X�����d8S�D���03l�K�v�U^�|J�>E�&(�h�W�3>�r轓ϫ�B�q�J&o�Y6��`�%H�]����~!�����"�?
��ަNnu&����n��כ��p�b����y����_�*�ء�;� iQ����2)8l�lvĖ��#\	��(Bq���!�'V�%$�kЭ�����'��J����0�X�V���k,5UQ&���6�g�`H>�/����X�YԸ85,�}>*qCkm��`�?������/�bv[J�2�~�y�ٽ��I��_d�y0g݌�ݻ��Qz@H?����7�����ډ�����{&Z��Sǭ�#i�Gcfȶm��{B��_c�<z9��n>�,��e^ʹRL�ڛ����h}�0��JQw9#��~Id���kM��O��j��i�N��<�"�Г�oz�o�J�t}�ԜH����v��韩��h�*�M���RΡ�Zg%����p5�T;V96�1g����lVe��!���t�l�%|�1*<�2�����Cc��Q�!�Ez`R�:#PG&1�� ���'UdI�3�m ѕm���ӢD�M��2��QobG���&��������D^Q�5��~�P]Q�XS�i��q�;��[�y>� �_ ktV>���M�
n�*��UP����Y��ڵQ�H�$͵D9Ʈ������.C!XS��s���VQ681������}��o��o��-���;P��T���N�z)�5��[�	�h�O#U�Wo|�kl�Q�7J���#|Y��l�EIOB��1�oi"�g�� ȹ/��p��z��a��^R��>���I/��K�]�z���?J��$a�6�U�s>�Ȍ��j.δx�hP�m�Egk�ග`��5���0�ܤ�p͞�6�n�wO�/�Uxm�Q3ZZvk߆{���n6"���f�>sS�U1z�2ӢtYɼ���^:�2H�s��Zư?9�aWg,���D&P���H�8�pt����(��c�(�}�'�|��H�
a��c�(������n�a�����@�B�i���/��q�v�%#4 ]T7��[��i�r"u尴�B;/f�`��9�O-F�{�Ql��lt<R�2��=�H�4�	v���IT
��&�Y���OU1hTύ���춻2\UM|È���~�7ۧ�K��������Z&yI�#�`B=-A��Ĝb�u���CG�F�1�̘Y�dq���gn�#1�> �9o�}����l����&f� �K�cE�D=,���1> W�5;~Yy�L�k�k��J0��������/FlET��
[�cMF��ҍ5�
c`U��m�xb�W���x8��j�b��%܈=��H�$�%�|�ܭ9�~���l����8I�K"#�m��|�s&�;�k�k�x
������^�ۯ�%��1B��u۫v���$�_EӻE�)]�cx(���w�E���,S���o����-�JD͞��9|��tn�-�+�\�b���o9�Pe!�Xm�ޕT	,�%��6����Y��9�8����B*��u��UW4 ��s�{D4x�����v�ڞ�\���AM�8�/�-��^�M7]�*��(a$X�v�!��
P�b��O#H��1��M����șS�&?6lp�̝�g��9���?�n#ײ�{�{���͎E�A)BK�c+� ����%G���d����G�zz�}=�Wf[��i)b�� ���A�4�_!�� ����dΉ������]*�lU�
B�:�$����?I0fx�6<Y����n��L�w�l�:*|��0u�{=w�����<6i,T��`�F��b����d[�Ҁe=8���mRYY9��(���+�/L��Ok��m/�mE�Ǭ�Й��9oȊ�b���Y�W���-��]Ss�P��M^�V��4��^�M�k�3i,X���:f��w�����'M��<��Ļe���l��i6��G���B�(�E���5|�����M,]#�����/����E�e�_��43���Y@{�t�L�����u��
b�+r��Hp���&�bm��E����.�,��áj��C?^P��u��3Hb��-���[��������"���џv�\s$�(O'y|��>��=N���Ekr�p����ɼlr�{�l�0��<�����L�	?����Pk���l+Z�&��H>Q+r]c�n����j�22�y��ݗj��b�tl�iNMqy��Y�X	eǁ���qh�ם�OF��oҚ�+`�j�@*���1թ��)�b����qRT�������.mg�G�8٪,ߥ���3�_QG�uq�#���p���⨂�e{	}C!���u�ȉ���m �xbJ�i�a[��);��h�a۵i��m�c7�K���"fTV�N'`8����Wr��"�I�����9���������U�> �P��
@��s�¬��n���]�&ڮi��YzN��P^1�ɸvX��Ȏٍ��LK$v���g��m�k��Co�Nc@
�b��>�_�;:r�]H)mi��}G�$׋ͻ���&h��L&'so���6`I�<������C%�o�R��L�1��4�=�g� 
˝�]����̲�w��'��oI̿����13Y���.�i�܌p��0������N��t}J�lȐբ�;H����(�Ȑ�7�*����Iw7����&z�����jJVe�v)��� ��w�	fAO4[/%=wD�\V�Ҷ`��)�����~��$�C@��a�Μ���4d�q	�c�c!FЭ���Q���_fe�_L�]&��HM��������q�����6������|�a�����+pbӉ=&�:.����j�DHLw�/0E��	����X�3͘�VH�_�ǅv���3�,�\}���~Pg4)_W&6j�0�_��qd��Xr�����L���#��-�F���WD_��u<��h�3�Iq"`\��C?�k=�e��%��I�/��7����&�3n���ND��cKH�+�n����иl%�>�di������ޒ�c���饥
2�(���	�O���%��Y��\��B��6�Ԭ�J�3�?���,�ޅ~&�t�g@�h'!���ˣ��������kQ[�����R��u$��Ie2JYM�v����" ��(=����j��?4�lA�|�!��k�4��:{�D���������N���"�#f/���e�����t�~G�C��I�j�aKcgq��{���'O�>Hs0�ӿs�Sf�j`8an��U[�r�f�1�a~��Y_��a�u��y��#n%D�=E0U�>�2N��)������Kͬ%嶩i�S��e=R�.c=�ﳃ��!7�G=��uP�|w$�q1�L���B��(t�^񼔔��M�X`�R�I�����Rx��[z�̥�!������f��]l)M��J�������j!L�.]Ꭓzqc����?�k+��m��^��As�YNK�2���%Q4�}��{XiOmWu�x��'�qC-"'d�Ax�<����2�����Y�Ʒ�*�5���ɕ���Jay`�_��R� �0m�陙�f����%�ڷ��`\��Q1)���+X�������a��0��j��b�x�]�G�T�dU���^Y��C���!��@�g3c��s8�6�uo榺�u�$qաE)&��N������o�������Tq�\9<6;���}�c 'U5�#�M``�����l��l/>�
�	�����5צ��L߳� i����<�P���輦�O�$��D�CǑb����43d��g���vķ��ʡ��֯?}w���km�x/$�� �ʏWC'~y��?XS�?^7z�~>9��Ox�iW^�H�/j@�,llԫ��6O���٩��W|��T�P��5���ð/�j��� ���FR�*}E��8�Zi����N��8�;>�% q�W#J:�g4��.̏o(��+B�e����\|'��������r������T�^O�֛�5�h�������H�*�4-����IB�6^-�������f�u��zt]X�aH����;+&�=�6!0.�g �'C��u��"H��"�V{ǳ�g-����Ӌ(�n��Eh\p0b��h�M�6�J2�Ѵz�iطɈ��i�4v���؛Y��&��j�㢀}r���!�[�f��d�i�NY��u�%i`�e�JU޵t������F2a� �Uۮz"�,#�-�{`�q��PrgLk�ɓa�Nۀ�V��>����s����ݘ�8�Q^!c|,�n��Ϟ�����~[OrT�vȗK�,
�f�f�"�]]�`�J��0��w�(n3jt�--I����M��uͭ��,l�Wfx���\#�|||Y�pj�_�_�͒�+��WC�	�]�:AQ����R3u�E2�s�O�M��e.4o�2!-Ɔ7�������
��]��֛ogʂ5Q�$�6�L�>�`L�voљ���V<MAMm��za��FJ���"
�90=���4�^#E����*�d:6me�/�0|�}����<3�읜��i~r�������<�.�d���G"wƘ��<R�OT��v}g�W;۲�Ϸ,��� gy"��ZZ(�8MF�"�Ap�V������h��%���k)vz�Vs��d�#@��쪱悁�_�S����ԍ\����������<V3E�:�ǳr��r��w2�al����"z��]���O�x�~	P^���oL��������VQ���t��vfR���nD��4�af��G��>�p�J~��M�ϳ�}�CVD��ȋ�jL�O	�Ґ(<_x6 ]S�C�����d���l�f�%(�F���=�K��Vw��5(�� ��H[��|�yI������c Zwʱ���*5���^kw�q�����e�$� {�X�P��Cd������m\|'�=ҽ����f%�������[O�Q�s��8�X��'-������Jgk�u�,�J��,0��,gL��R���������=�&�m�`�s�u�\�r�:���߁���`��^��9����x�oP���H�fT���D���}é7Y��ρH8.�f���X�|�w���A�,��=7]c�?��OTe��J�[�4�� k�C*�Vh�y��c��g��)2ν���1;��9���ά�r�hM�Igo<믧wg+#��:����2LmAi%]��|����,�2X���?bۅ�?���+O��r?S���>�y��Sk�/^�{ڐ�{�o�&�X�>>>i)���%%%��g��;�ai�n�x�O���2޼G@1dL�[��^qHe�mP\;xD*�t��\����6XS���9<��a��Y練�l�` �[�����H|j��/�*��E�� �]8��B���c��yqi���[�/D����P�Q`��WG�m�&#�e�� �=W�p�t	gFڛ�׫��rY�3'&���V�9P6���;�6n�e�Rcd:��������ȯ�Q���I+�,s���I�J��$��P�ҙ݁1 0�I�90&��֥	j�?_D��&�F ��*=�� %�8T��t$W����J�{ӗ"쏚.3��u?�&Bh������3�������S���ot�innN#�/�޽������
g�j2���N���(N?3f725]�ja�e��i�9��^�|2u��'L�?�GÜ4����ndl��~p �q���I'�oQ7�#���2��!f��h��8 ���+'��r�Gx��R��w�2�ne->��cnZ�#\�u�Z�BW�jn�^*����<0F�����d��L��OG���ռ��>R����ٹ`�X�I�w���v|�M��1'6K��q�o�O4��hv|C�w	zw�	:���oXx~����!$�R���m�L0��&
�M�u�E�h'$���e|�`p����s����!��,��}��?e�\�8��9�Gkܶ,���%L�T
A�����͉����V"J�D��r�g�@�$)����Q�����7"�暍Z	Z	�H���{,;�>�פ�Y�U��p4T���$MP<��EZi�#��#9�-��||��#�<�^z���P���Kp�g �����f���Ϗ!������^y��秜����D��RY��!�͑3(,l�B0(Q���>���-
ɶԞ�w񛳔�z�zQ��������0�i�cZ�  ֹ�<��=�[k;nB1��Iy+]�z��Z�Q+Xks	V��-ϥ`Lį-vԶe��' ��.����8|�ԉǍ���7��>I��|�hfp7Q�:��gR����������ᴙ�6��ZЙ��O�y~:c�~S	�uu���0�p{��(؋��t�4m����#�٘�A�U<ͬ�KR��,�����]�#G���Q ��`���LJj;C$i�O-�$}B��㰶s$�����ťq���#������z�
�'�6,����f�x�kQ@GV��"�@-�� N���׹��Pu ,�ϓd<>�kɋ�l3���N���nĘ$�:?���p��>D�&>;� �E������F+.]P�}=���A*���N��iܖ�������/-`�T&u-og��+S=bPS�d�h�8�.���;�'���n>�>���|��<�I���UK�M�	��I�R�ژ�X���0�wՍ���v�%��4$��Fԓ;b���a��4X�64([��^P�N�#��T�)k�����y򽡦m�O"�8A�r�� }���<����Dĥ� P�/�#L0qho��B��rR�`Xϯ�}�����N���D�����nXA|�s�y�?y#���c/M�����fNO.��y=�ۦ��2����N����4�hD����\����I�`@Z]����6��fݱ���϶�ֆ��I`���BMH�E�0�,�^q��� �a1m
\�ȋf��lb0ye$���\��]�`9Ј�cW����iA��l�`��Da�e@� 1n��7�Gԝw�\A��\�@����`���"���#ğ�����s�8~���S�Wd�`���m�е�5�VVl��=0����=�a����6Ogiq�=�Yuu���s�h�Wl9(��2˛i��)@��^��9k��9h�1IL���6��(��z�}�0x��Qmr냭���bg�4�k䚱�P���Sd��{�q�-W`�%��f������z�sp���s����'�b&�jOc���uK:��?|�c8@Mj]o���=Z�z`nh�Uޯ�5��X��������^6��od�=�\�1�*mc�{����
�R*�����ͤX�W�R�
�;���A�	���ڱ��'<f��1\���_"x�]x�k+���U��YB �U�D⯶�Bqʦ�E�C��Њ:����7>՟��f��5�A�x���N�.���P���K/���'*�ZD`��>7�*����)�]^{� t(��P �N��`\��I���zaaA^t~x����W㽼���Q�OОЪ}{�+/���f�=%FY�v�t ^0x!;��ɕ5�G�:ŭ��Y�H���
o��%�Z�o+�.ܟJ\��dtf�aK���?D����*xǛ�Sˣ�0�#�%41W� ��zöS�������|ɬԣ�W���t��e�X��CW��k
U�y{��d7�<w#�Um�o�l�({v���Ū����х4ls��F_�
�1����$t�������<���������x�F���G�[�E���t�t��tww
(�� ����%%-�ݠ�twKw�߃�s�y?��e~��}�ֵ�u�Q��nr���7� ky?��\��%����y �ҝ�3�'�׳{�n�l��"�K�5��>���Hl@�8\8�dpݠ�a!�i��@��³��s��Z��|�]#��Y��	�;��vt����\m��{)M`=r�ѦKMS�}��,��5LVOVQ
!i��\n�-���i.th�F��T�x�G<K��+Wړ��v7�b�'MSk�� z;f�aӟ������n>Z��8+�8��{|t�@i��d��v|��I/���y��� �;�f�<��e ~ ��;��]�@H �����z� 鰻����&��$��1|��+R1D�6Ȉ�ʳ��5ނA��6��s8Mu���d��=3:�ϗ����2��E,��5ɺzZ/êl��'z���U�X�S�x���!�R�������_�����ta;o9��uH��vc���gG��1t�j~�m C�
[p��Qff�M����D�0�	5"�ᙡ���Q���H�	�A��Ѯ�vB��������F�Μ9dL<a��*!*rǟ�����ɻ,��XV:A��,!?A��Դ� ���&������r����ԛK���X�$+�r��!��m�@�8po��;@a9��V���n[e?��#������ʇ?�B6���M��J3��:�޸�w�7�w������B��,�����@{7�B���OjȤ����� �7��L��{bn$�է,�SaF�Al���,�,RNѽ3� ʢ�< ��͉]u`��G�1I��a���z.KԶ�ky%f�砤���t��7���LX�[$aw�R�Ik��GB��� ��q4�`���*�}S�^l�i|a��T:�Ss�H\m��B���KL��y�����8�c*Հ�Y�l��H�	���cY�aq֛�}1�\q��۷툚hx�X�]+���"�@�[.Z�$�3���mD��"���?R�%ی{�N�u��at���y�⾛t��?Z1�B܊B�Mi:g>��2�Bu<C
�b˲�����F�}T�HS���c��cd[��2E}�Ix�a��H��M×�0�(�U`����w"ht����h�㲪Fڍ!Uu�klHE�j/��/�ҼU3�=Љ� DZp�;4��> ��?�ܾ��	�N$�7)��� ��^��d�D.��	sW0]@n��6
�8(��R����e��� <�X=E��\�h�j��EWwދa���(K�I�G���Ҏ���_05�`5V��}��/��Ҿ��ju���p��a�ڕ�)��e� �e��[�ŧ��$
�A��ᆑ�"�؉3��6ı�[�P���j�}�i�=
��`]\��n���(J�U���vD���^�{᳋�n�����~�c�J�=j?�ή\���eBH�W�v՟P����^Pk~�v��J��h�w7�ج���v�����㒼�&�����E���f���⍊5�љy׻�Ӥܨ[�~�SM?d�ǿh�,Bl�gOX�	Ap�'�&%�G�O"�P����nE����=���� �K��2"a�G/�8.��j��8���l�F��?2,���3��;ٝ���h{��IK�{�g�x�
���{��h�����k���@�����OA)~��d���ͤg��s���q>G9ؚkdE��w����6^]�[�Ā����*l���3�Θ'�pxR<�lM���oA[>�_J����edn�C�ꋌtp�����H��@��|�@��&�5>:&�|�ו�[�����"����k9t�QID%�Wq��q�*}�Fc׃����q^� ��,�K�-�O`6��R g� �9%p)\��ئNT�ֺmeޖ�C�3��uA�����v�g�o^��%�2�'.�;����&�?��Y�7�hn���)��fZ���|F�s��T��PH+z�k��ċ�����儋�`�=�k��	^:w>�5��l����g_�l$G�P0u��	�y��1(o	�͍ ���������$��@�zl������'��V�c<�1�e6z������,��9��?TGfv?^i|��Y�hw�k;�Fl[��
|�i������\Ʌ���^p�vZ�5(۸��6d[�s%����j烶�☞ǯ�����L�K(�֞v����������lN��Zd�#��=m�p��L�S|�n8�	g� a++c�5�؋����1�.C�ސSE#^��V����)m-�x��-7�8��a��4����Y8B��+j���O�Q��PL��q{�pT��ݖ>�:��,�{oG2�8�"� ߢ��{7H���̓{*'@��S��C%���dbx�xP�櫸9���+C�ВS&��� ����*;���}�t��5o5o��sg���Ep��D�@��Z"��-Ǔ���c�#���U��p	�`���C]��jtX�^�ٴ^)gZ��\n��۠��2�����\X�|��bw�p���ƶ�����}���������^q���	��G��g5Tt;�(خ�ܾ�S{�[{tq�'Q���_E�x!{8����	�oQ��lx��7C�5x{��l�Av��G$mMDdo4`N�/��ԡ��o�g9A�|(�@���@SR��k����j@-/�kk�7�vA掐u]DiƱ����r����|�[=>�����xЌ�j���wV�������b-S��*��]���1�IR,1�1(��� 4Y��_�[P�j�}G��2�![A��L��
�Ɣ��/�Y0֭��E��s-w�plފ��ў��e��&��]�✸�2<�^}�"h�/�;d�x>�4I���#��{�ăM$;/jL�m�3n�-\����\ف��=L����r��%i�z˟U�ߙ��B�9�8��;M����^�b�%&�]$��۫�˗5]U=1C��r�h��N<�*~塇��t� ���>0�,P�h��*�m�o��Lj=���{��D�$�.��r7|yԂ)j	:����#pQ�Њ��&�.�o��"�e�׋b�{d^(�RU|t��Ⳡv�Ŷ��ا��O,��!�4TLO���T���/��Fh� �x�8/���>��Hp�KЊo�ݡ�1���n����D�9��6���c?� CR��?:����G0�9ZI��Wr�oP���Z��b���wLnϙr�m_�Z;�O��+��]/5�z�P����Jp��H>������nYv/��yܘG!Yj�n���?�v5�����P�ٿ���Y���V�y��T�p�ݽ0��X�=�	�pX�<B�<���7V�p^�������[X��@�ȸ%�&�QK���J��_L�0���f��GzsU&�n���y��Ih��n���c�y�������v�md�v�l��(խ�o_�X��!��ڌ���Н�}�*!�aS}|^���-��a���T�=n礁%v�󼲇��� [��I� �W��aթ3ε�XeE����k$��[0�̟LQyz�n��ߒκ�mN��~����!�)�=l�@�F6ț e��/���|�K"!���s1�2$V3K���d�m�Vf�f`�P;��V�!�#����cch߱�(��l|��?�B��S��k�GR��T弪Ry��g��m�X�q��_0K���}&�49Ό8J�Aod�����pC�-k����၁:V� �X�����AF XE���8ᖹ��f#�(r�zÌ.��؅ľt��F��^c���5��Ӟ{�_H�f��P#�3)[	������Hl�qQ;}���s��*`�����4�h�)�?�ЧnYy������q�5�9T<<�J�ؚql�UW$����
��R}��<�E��&��$��Y2Ȉe��'�o�E&;�Tf��O��fE���O_-������'K�B�08ܤ���IQ�SR��N��/�`9�� 3x��ۼ�E@��?G�X�±]��mQ�n�؍X���݊�XA�����<9X?q?�Ò�dU_fg�{��r�AtT����:}1�)L2Ձ��?�����NE&D���|��^6���f5�b������7$���cy3i�;�œ���r<�����sN���
J_�S۱ٞ0�∥��1P#���\��IY�u@�oa�NC��\D��I� nn睱��O����g�,g+��e6詾�حu�S_�����/f������6��6]�:?��.?'����o�,(}�ى��s|W��͖��0�UQ7.Ξ�ʜT�e�[�n\1�
����p�zP*Ĩ,x��T���":rs@����峙�+���^q�'4�t��{ǡ{P$6��q�v���Z���ߎ�R�F�Q�0Y�a�����8��7	�Nd�m/��7CJO�^vǪo��!3��ĭM��&�qA���`��#T����A�0�S[���F��6���>���Jt��			g��9R0�ښ����f�������CH��Hi����`�=8i�S�B��"�������Դ^'e��|{9Q��~Ym굾KnG�T�|�oo���g�{�mgR,}I9W�ľ#Mǳ:��3��x�N<����/��𜮻�/�_ &�(��#@�R,c�AZ��Y,.���g��yX�,f~<� �,w�^K�u[M�Y9q3�hpkp�J����h��a��%E^ ����"'�줚�%�$�´G�i����w	z6V�Ї�U\��:�9��J�.䒴���{�\��q$GAN�V����:������,�Ɉ�����&�$����ki��EE1���e��Y���d������=!�����k�KĤ/�܉�>m#�T�&XZJ'9(�;7����G�r��5]���:���NZ���ņ�_tt������z�+�78�4�4���԰zz{1qqъ�"���O+��{�:.++�c�m�Cg7K�'%�6�'+��.R�"���ז������*��Јw��/�ID��q8WVWO[Yi0N�.�SY������N=�����Ǯ������E��$ՙ��Bl��?�a��^���q�`�p/l;�����)��$� �Ä�TQ�2)#v��?lOOO<�Lܠ��2.�,�Q�}���@TO��}��H�x��%�^�]Ɓ�A���m?`g���U��CQ'&�##{�|O�1yz�+�mf~�r�����n������ީ���rN��CǷv-x�GK6�Y�C��@�Q_E4h����)�Z/���Vw�������mX�͇5Fݢԓ�gá�3�;��$�
������J�	�+�eH�?����⡠��[ �sW:�kT2wq	�a~{�����;�}}�����d�ݭ���1V�¾���t��ǘ��T��|�|�/�6��B�y��V����BR݄��?*Kϩ$syl�R����zؓ)�Я1i��f�tP��t�o���J�k����yy�R�./�}��[��y��rSA��g�D":�?~��Y[�C��q���%%�������#''�q-�|Q⤹�E��mc݂��u]��TINK��߿���Ѹ�Yc��SJv����555@���8�j�D�t��.��ٱN�ٰ���֮'���v��2gg0
�@���l�wU.޸`�����ߦ�B>���6����q��1;�����8�w�L�����G�w*t�?):�='7�����<z����H 揊�޹�|f�ƅ�\D(S3���ff�L�zuQ��h��c�+�2�B�̸4N|U��[ Uj6�1%�Ә[��Z�C����=NQ���6���ƅU���S.��< �?�k�ܥ�R�l�k�~��tff�p��ݠ74����G��m�֓�KG�xs�x*M�z�����i�9�f��^p@hs�O���C�`\�s�Gv���PNLLHW{{x�Sq@gg����m�u����6>�G�ӕ�3��z�3RQ�i'�~�9c-�S�t2���5�l�(z�͍����A�d�-0)�R�w�ζs�O��10`��[:Č�Q����;O������=j�u�������"B�5J�0F����U�E���斗��铌�|��_o�i~�%���<���C����� &B��/c �ȠىF^~GVV����~w9����T�L���uX�^�p��>�N�6��²����&o��{;��Cã�ţ��U��Y'''�Et��]Z���h���憻iwc#�*�%���0R1K]U���Ĥ��8�CgUUU]ؔȌiq��s��#X����uWIKs_B
�g����R�tBGF���-�Vf�{��q��, H��M%����2�
vv�������.��J�y�3��N	��m7 /%���Y������瓩�����U�#��/n�پ����[�dx���oED����&Nwu�RSS�}0���u���^�VQr��6�a9��p��{O`ʡA+l� T����q��#q���	+5#rw�\��'=h���떶67���vx�F�ץ�й����>�MX�������7q"�Mb����O�����6<���Ԑ����Y&8�%��x���.#*0���^�?�֣A�d��ajΗ*�b�:�c�k�
j��'i���YNi��Gd(`�b)�x�����(����|�..&�{X���{�?��ҩ���av�o�1��AE�3��n/<-i�����^Nz΁��[q�ᆢw��L��	�����d<z577Ҵ�j��J`�0�`(��忷tA���VoBґ���3q�3Ӽ�3�@�)�F���nK�t��D�@�E�����8�}Z(�:;� ��{xH�yׅ�5� ���Z�d�XG<�EZ�EAE-��x8|���6.9��ve}<@�|y�#�ܑz]{|�B��c�_x?#""�14{f�T:4뚚������2=�@񇧢7�9^���3Z^��؎��#2�zw)�g����6aFF����A�⍧,%����2R���~���;�wA��vrb�Q/��D�'���ښ�kө�!̓f,��tީU�i�A�����%�Jc�Hz�F�1���2T���7ὊWTV���W��ڃ�P�� Q�o;~��G	�	�{!!!
�*n�}BܨI9ʢ[&� ������=<�I�[��f]�۞fu���+��Q�R qO�l�XYYy����y�ԃ�� $ģ�
%�өo;��6V�J���b���<����!/~�Lb󣣣��Y��,DLL����ЍQ7���ߴs)Ee�S2�0
.\�yIIa���}��>���ɹ�-���,�^�?z{y|��V�i;���W��g�X�\��x�S��i��&���e���Ayj�YETV,V	^.�m���*u�Ƥ��ڱ*����=��['�ks뽮��T�����\m޸m��ٿw��N�<��Ej��g��F���#sNH��-�#�FD) ��O:?��U��PtQ�B���_�P���y8�����1)f�6��^��<��r�3�����'�b�Fަ��%"++ �g�%[�E�t��8CP4�LIۭ�0C�_��I�~hĈ������*?�fF[���W�
���\�af��;�t��n������G���C�q��?8��,5aއ�j����ʆ�R��W��=Ɍ�������A$�)Hz�sԻb�j�$e7cGA��ʴ�=?A�P8�T�����H��eӚQ�/�}�l����=�Y $-���wM����^�.�${^v�$���2��4BDK/ ���ƭċ�̃���*��+f����T�iL��p��I{�r��F�ʡ�@��l��/b�l尖E���
�_����z8+^��z���v����q��)�
iq 1/444>-)*�y�*��r��Цf`t5���9VW�޾:�ݖ�"~�b���xbU�	��і����W�����?������0��87�t� ��ʬ=Qs&�5�RPP�U�'7�u�����J�����C̉K��c$ߨ~(Q`#Q��g xl �����R�E��^�T��5�;�X�⽢�k�`�G���^�	���u���T?|��m{{�A�;3p�2�H^urNFFd�&%���i&���	�	,�m
�-0A�����[��:�_�Q��f��>�L��=��)���$�~�����5^{KZ�أ����1e��bPD9/��do��4l�<FH�pD!����b���(-��fO��^�;�A�>���Fx��y�@@.Ϟ��mn��^ݼ���{�����~�K����a枢r%/>V�|
�:6�sџ!�0�2��O=��L��ouuu�srоg�eK��?~(hpke��tGNÅS����+��b�c���
��ć��+`��9��RaaR)�~\�%xx*Jv��R�&G��Y���\2ldaS�O��Rr�l�����:o�����!�m�p_L5��]��><*���P ���b��o���ݖ�I�e�?|�( R(l�R�}�J�Ϥ�X��J��`tL���9��Ǐ��H���W׉�j]ƵVW�����e�y\[Mg�닯 0�i�1h:9�W��t9TD����t��?�'[�����X8�����5'�;������dyE%��rsG�W����9=�}����Č��-�,!������𩪪�A��K���[�k���5Tb��V~f�kH`&$�qP>�kttt[�vl	��<�M����|m��#`6/i~��������ָ2���n��o'�|��w8��k��T!H�������b�,��^�&dΏXri�.5/V
T�F$D�ԥ�?���,+�f,q`��EX�Qg^Rj���O�&��:\QT�Y������:ӽ݆S�|�#���: ���XXDW:Fx���
���@;��D�(�\^^Ҏ�� �O6Y�O��*�GIO7R
H[�lX��>>��;�S��v"���z"sp�Jh�Mω��H�a�(���琽�^2��r�O-�Lr�5þy�a�v�XMtB��/��Zݘ�A�j�g�m�XB���t]9�[ʆOF�b�*ggQ����Be��4��}|ؔ�ŵ�ѱ�����`��13S��۸v�:B����E��ƞ��c���oy(�q^�&;.���xQQP@�%=/2�������!=��l�;;�rN�M�q�h�ƮZ*��ߗ����J2pݟ� L�������NN�Mr���}X[�T���G@\P����)�ޔOM�fk�?.�O�q��E]v��JRF�����$�U,C3�S.qu��8ͤ���ދ�hs^f��/;��$���($?|7c�I�&O7���1U��t�}�q�«���/g7KOL`"�&���t�Bk��A�}�;�]Z�^�&c�@��|jLr.8y�&���������	��fK�eK37> G�C
�T�=K�����a���+���R]\\�厍)o-�׷ ��M�N~2:�8NHYH,-x��?-3�¶W,�?��V�D0|}ݰM��E���JBJ����w�&�o����=55����N~q��x�-'��8���hK\���e��iށw���-`M��V�-h��'	G롤�~j��P��,|�JJu���Q�wo�;�s��Y�¶��j0uH���-��1�L�D��^]]=s�kr��-�795�C��-d�����n���0�}�FoO��	�S�UJ]�Ow[d��_�'�3��K"M7G�9���gRc~@�O�{�}q\o�df"��q�[�D+ێ?&������KL�8<f�/�4Z���9��/��,��,�5�>3GG���N02k���=kkk�6L� @��+���lH��l�� �!*�,DC+�� 7��ҚP��4:OK��y]����$x=�?/�;��45���<�����[?ܳp�^���TK���i,����"�?2����rrGG�\hXXBnfX�_k�"��͋�3�	��6�. �+;	`�^���+z	�=�"!#��#%�C�ُ��<0�ϸ��~�7J�����NHR�I6n���X˝�5j���(�+V�ޞ�_�?>+��b}w,����\�ݗü ��Ή8�;�t�|q���}�f��	�͚s�����/��WY�o��^ E�\p_�a�C���ݏ~�	Qz����E��M��M���W D�|���ح���o5�=��JPM��B�ioo����}�V��l�,��^� )�F��q#�޶޵�7��m)��c3�m�����f�����h����g����m&��Do9�$qV:�*����`l�P�8Z����(�x��}�͍�n��ǔ���H���ך JRRm�������q���=v,d;�Z[[�ѽ��a)�!��`~�2qܷ "�D�J�ݺ�8���D���0&B��${G�r}C����*���Z�{R23����_g�J2S�����mR�a��=b�B���J	[ݬ�� ���))L��|^���|��=#CπK���=.�0}���K����!�8	������9���F��������
�F�%%��͞�H�ډ�]*�>����9�aZJ&���)'�.	2v^�7��2q����X�B`��������*���(�j&Q�z&j��> �%%e�{:|C��x�����2�52�>e��n�{�����>x��e)9��ޣ��6܉,��G���I'����o���qd��a�BB1'՝�:6� �����5.� /��c��G�- z�hMT�m�99�l�\(�nfV֗6���V����`��[�8&�3G�k���"0�0����	�Q���-	~i��g��IQY�����&�N����||V�I����HEE%95�R��u~����㸫�n;I��'��%�8��w�ei����%!!!��}[�#�x��  
����eff&<"�[^���3����[pc?ձve_�R���j�!y�F��S+c�0yn5[�a644�R���	��g�F�5o���%7k�@�Ji1�)W�w�'�������]]]�����yE�r�ôQj��D����$0�bN�z]�앶6i@�/�@�1���$[v��|�i�x$1yrb������/�J:�CtmvQz`���F;��G���~"�&(2�o,��ӥ�v����$"��,��2pn��Lʕ{p��<W������WP�Wò���S=W��pi����Ftq		9���~X�)5�}Z�_����wK�nj,�����O��h1�j�ד��q���^*B��=�EV3�����)���,,D�-뢠�����29�0 ��O���-�&����x�ӢV�O�D<���.o&2	i��ĕ\���ka�Bx�wQ8���B)���ZN�H$X��p�-��q�����L�*�;��3�/`���̈��O����]����@�?uM&����+���K�W���w �:~�4�|�C�(���{�����Qy&��`oo<W&�y��l��CL����꽁�˴xPѫ�\{8�h;ی��rR__Oǔ���#�#w���_铌lm��V�4�Z���u5*ϐB����ݿ!v~'�q���die(� 7�q� ��x �E��A��͵����`yP�y9�1ȇq/I��ﾨ�_�R�����{g��,���<��CGY��JQ�:^����n�qa�|���JՁhL�n}M�� }b���!�=7��tSVfig7 ��g]�.�ʎ��I��e�����A�B�o
h[��}~��ebd�!����OH
�:rp�Q< �:��W��I��<G`���|0�cy���'��{y��;��Wѝ�7@J�~�f
����������Ⅸ�a�"� cJ�;V�t���|Ej�
��%)$�$+�8b�7Z@5w���������9ơ>W����(µ�� d,h觻Р�\��������_7��;��w�w���u�3��Z��m����~6�+�@�>x�/���_�1�R�S���"4��Ma�Y�$Z8�WՀ�(9�fE����!e����l�i���Tgj��ǩD�N�z��v!�o��m'������X8�
#�-�I'��tr������>h����+i�+'��@gq�o~��į�w��{�T� �n.����&��ާh*��7R!$ґH0����s���4@�ۘ.S�E^����;�SD�|�sc�uR�ow{y+��s����8���	W����W!XXX&��Np��B^�g��oܶ6��ᓇ���Ƃ����t໑�"T)(l��Ծ�y5���7W�#����~��:���0�O��f�
��������粐��WIXR\\P�~��l������~��ЯHN�\9D<_��8^HN);@h���Ӆ�d��Է�e���m�da�:�r��L�Y��ڿ��bD�SMU���'��E]�%=?�V����Eε�����ͽ(ToX��������:��	����ɖw�n999bѼ��FN�H;�Y
��0b��v�,�Q��Q��!��蕙�3���8,����W����q{>�d�#Bf����C�k�Q/��S!����"+7���LNn��va.T��1	���V31��������-��g$�;���o�u���V�,MO�Wgj�'&��k�>�
��W�"VA���̕�"�k�'���� ��u�7��~x����%6�!a��ɓ��]*Kv�N���b�͙[X8n�P�]��%�����{�����)pU�no�*)����z����[i����b ���-�/���-�����X��8�G�#�@�i:�e�k5� �i��"��\r_�ig�Q�D�􉹠�@�#.*�w��(��t[e��0�
�	p�43j,Vyr���$T{%"y;閉����kN���L�̍���Sc�rUu�1��3���� 8�>'a. 
�N�|fs{�0�߸�|('Omim��rVY`���v�/o�}αaЯ_-,��R��[a���BQ�$}%�~^K�*ԓ�C2To����! >9ك�H�^�	���J#"��i�0�g�����$$\�ڀ�~�l���$������G �tm����������5#��?��쟞�}`��`D���|��U�)�U���޽��w���������`�����BK����$�kAL^s6~������	cB�m6M�������ӗ�1�����8 &^��A$̤�:U�D��N��Wy#k���׾u�V#��N)��gZՊ��hD�utl���V�������f�P����a�����;Q�ps`�,����`Ak`bd�����mB�:���V-U�Q�g^^��C%Z\�v�b~���/M��)o("1f�p�0�Ђ]蝙�)f�����I���_�t�P���s�%)1��ʗD2Ҽ6o��(��4i�(S���vu�}��w��ґ>4-��
��S������Q�>������ �*�2����p��[���ĵ��C����jT�M�P��6����mp?sre4'��%�}G3��U�?)���#���u7W�(�:8��l=1c�b>���_��&�p`0Htj7�Y������OH(,>_Ke��b�� !K�����U(S'�?O�4QEM���)�^�u%`��u���W%��\x?���bF*EZ�4L�`�UYY�&$���U�#�k����64�����p���|%5��'J!��D�+0-G-3c D+׵�=��9@���m�022�57lm����T�O�`�d�z]�Ł��wCoQ��y��}�\����'9��K��VW��,
h�k�)�E���OϤ���4��5?P��~w6@��U���������i�
vGϬ���N�Iփ���M:3�O�̹ffE�gߝ����������/�lM�א�^����h�2�fkP<�d	OA��/wWd�/��JJZW��\m����-������]�d����#?������%�M-J�������c444�|�e��!@���I0��N<�h�(��fh6=��D�D���X`����y�!yDO�2jN�	��+{����f��0'd��k�$l�~S+�oUR˴��ի��7f����m����;!-�F�AK�[�H�E_���
�QY��4Xÿ|�v��}�7���"k~�FK����J����:��3}��+�p Zd�A��TGH@*��/�`���lR��̲I�hǵ���eap`�B!�s2�|���=���{y�|�xv}]/X�M	����>��z雩�!�-pI�!m�C�ՁX�[Z|�d�r�E@B���%.R�J}��<y�t���Q�����DMb5��:��ښ������
b�ތ��?�Vc��z=�c`f��{��{L�͖��Q���t�Q�ʞ��58(w�S @���{�)v�U��>���������G�	AEE�۞Z�!,�_\ <7_�'6_����?�?�I;[�@'ԝ:p��v?���7t256�Jy�LN�(�i���X�:H�Yi�����M>��IPkH������`9ͬͅ-g�^���<zIr� ����k�1��i��}�յN�{=�`�;;��*\-���/��V�Դ�1���ɻ[�[Sb,+w����g6�@����pVj��e����C��ӹ?������WA��_�8��Kk�?OD�6 *;�!V1��V���։�L;n@Tb5/k����ָ�L�<�~��>�vQ�/����F����vvv��'#���L�X��c���9���#������i����6m#�؎̎�m�Ě־p���QXM�D�YSG����(d�
p=}M�@�k�d�OϷ��������k5e���ǟ���Q8�rpL@� �e�/U���f���_e`���AZ�vcqy�G�5��k�ze���:}fM����n\�V����6��W��1�j��"�0�p����������%A{{��Ѿ�������������ە0!o������i,k7�n�����*"-�����{l\#��`�IV	Q�dF%����m�1ו����V�X�����ؘ2�\g:�D����������J��()e!O�
/�Dkū�fl��v�$7����*�����*K+���w�׋���P��(Yx�rE����&i���%\~.L��س��� (;)�qI�O���\M���.'����P��՞���nC��nF�H������).���1�t���)�F�Y�ʾEW���S{�JQ� E��fg=ܨ�Ycͺ dQmΧ�1p1�_U��?:�B òD�ܱ�y���~�,u�1���9A�H#��(?�`�}���F~V`;����#)Xe��w��>� �vYW���J���hj?	E<���E�C���z�w?\���JTu?���� *��U�$d� G3�&>�c>C�o&_Z䫲Ch�5���U*{��\N�ѿ��3)
��m��<�W�K�5p
R`<��d��5��y�5����g��0Y�^z�͖����]�����-*
��[h�o���M�x��z�5����n�ٚ�yy�1�9%q�WR��0�����|��"���6������f3glhh蠡Ɉ���Y0��k��]� U��N�:�P$��Qe�~�n �����{GD��`*��3��{�:�T--.6�m5���=XGaO8�k�ú٬� Iѫ�V�$�
&����y���O�Ԧ&�6X2�b� K����C#��?w�씂v�p{@�ܘ*s�`���i�/m����v��*�^qykk�V���|�����`f�:��\ms�aI9�ϼ�I���DƏ�bʱ��Ĺǒ��<?��SRR%���0|��[rJ��f�����`pH��G�=W�;Ч�&a�Ϙ�J�t��H;ǟ]���Y��i�W�����6��N���^V_��~��|:u��&�\inl4�G��E��o�ǈ�g[��l�6�
�OO�����>�覣g�?�|��ګ={��[�#yy?fd��uPRӄP.���I��K����Tp��B��g:����B:���-�"��6l�;���M()�����zDi��:]8���3)�1�зN���r5�����k��+���n��ֆ�>�7�F���V��]j�di�Z0e��ʝ0�c%��9p����z[�+*v���� ��O����.7�>,�r ��*�t�N�u߿�
�Ce��ʹA��T���^��K�2W�������2�ߓ�3:��.[�r�������}���P�L������"(�fd�i}�z�U�R����������ԡӇ�����ϝ]�脴�k�\"���$�c0�=f޴�����q�K �
sr<��n�/>'Ci���Z�^jk��?�Q����ǌU��;p��{���#���'��@�ӿB��:�%�,Qy�6��1\�?�����ډ��=� K
3'�#�٭lE�<��S͗�\:c�ָf�����ɬ�z���D����FZU��
���;H��-�޷F{�_Qt(y�yc;����g))���gdg#���G��=t.~&��|@
C'�8�! �}V�.��G��w-���A�5#١<�������xg	��2�}�O��B<k��I�89��]  nZ�ѥ���ɈZ�o���h�F����u�:s#�" "�ն�YnV�O��.�~66�̀؃�?2e��� $"<[,�VMd�=�]���~��ix��.���$#���E��UHR�]���I��b���;��)��'R�$%#
�e����͜�1%����^��Ԧ�«��@q���~�_}����f������_@}�ۍ(��(�t�
���k�0�QX����ck�ek�QvV֖�4�'��µy�,�������ghgX\�� ����ތ���ά�W�u�\�zx|�9����~M�Z���;�)�@��~A�4<.n��&����ֲ+�	��4ꗡN8�z��NC���S�ݎs��M�m�� �Iڟ�}��Qk����D�!!g����������E�ړ0�������[Fe�um�
�Hwwwwww�tw��"� ��tw��4HwH�t*�{]z?���1��w��������s�k�y��q¦��2=2�̾��h��!#�;a���g��Iֲ6�����M25;�R1�B4O١��TT4�U�w��I�"�Y��,���s9�ڻ�980"�ϾT�/IMܰ�����#�o��P�Zpk+_Y�Z$&}|zVد��tòIk*����,�FR!!��n�&�������T��go��6����#w:^ih<wm6`�<^E��0���T����-*.N�ThZ}�B�0�ۮ�.Y͢�ʪ�_��<�z�KJqg���ThX�e@a�����6�Y.��P���Y7��l�|����(�og #R��0w\[�� ��+���P`+4�5˴q�$������Z��^?܇"�5�		�nv�]\^�s�&ǊJHϒ�=���u1A���=�i��*��A�|�oFɋ�0HUh��{㠕̔o���FHD�R��=�(r��� ��	��&a`�y����K�h�G��� �B�)B�Pv�LnT._�ixx����~��;H���S�֒Gtt�����=D)~:A��O	��Vc"�B��`��j�~�o�q��-�z{Z�R(��O�|Y��0��룿�#�L�ng/���:����rrH�7�x1�a����~S�������> ߈ ����:��(��Md����@�Pk2�l�Q{d�W9	)�4lxxdqss���ca��KAAU5:j�*p�LCi�Z��--�������eʘ�V��?y��$y�"1k�bg����l��߼p��/�����p����}m�$��� �����W�?�{���w���ҁ��^�|/H��䉎�r�)�v�Q2=b���g.�01y9XZ��Gu� ���3
��v''����6-�}���͂S�L?��q22�ޜ
�g@doBJ�u�Ҡi$��̬������Q���R;�k����%x����n�"���s�*�	[*'��(+d���zຯ�U�w�Q����r-�	�7c�At����d�!]
��ϯoo�Tc=�p��$���L^\p�ҕA��8��R���!3,��Y�%�k5�zF����Y�`I�����>�X�䫝y$څ�������%k9��4��@=����M�/����*���픺i擴c5`���ŝPRbϱ�'_U�i���%3hu*=���#�g��O/@d�^o�@z�2@�Gy3r��h�ʗ'ߢ�L�rv��Ē^�y'��:Gs������l�X_j�8eE��(bEE�n�)Y�j!u&���JL[�A��+&�5H�N����Z����ԧV�n���W�Q�z�О@�f>3�=!ofgaa��_]5r�t'�������)?b(�5!����>SU�	��FH<�ۄ�ė�1%TD��dd2!���!K�L)Kh��	�� �ϳ�T�Tv�F�slm����CbK��������EXyڻc^@�o]��33�Ggf0���ߎߎX��������.����Æ������&7dn�T*E�paY|���l���#�|�e�hcP#!3���Q[���$1�BZzzO:P@aZLh###٥�p�eZ�4x����q3�&!]�n�Y�ed`��c�_�7ڦ���舘��3�p@Ɯh�j�)��Y�Z0�d��y�S;D�xuw�q�5°��"��G�d݄� ������F.k����.����*�x!�y`�4�f����[G�"d�)�Rn77�skre%
`�nH��v�"��Ʊ	��BJ?�F����T�&,1"$"&����#R�A��)\��^�>��yVV��Μ�%P��+�SK�C�p�)6B+�����C�PvI;DD�0��Omǈ>?�uY�;s��ߠ�����m硳Y}��9��o�{a�F3D���e(TJ5RL�xiI���
��9��R�t� U4���B��k���05�/�F˜T���,ϩӡ�}�������ݬ���M��pS��V	����Gd����O,"��]uwC�Ce
���ŋ�'V�҇-��~k nk���\u��fD��(�����ȇ䐱X�2%_�jee��a9Ttt3gH|mf~�����-�X&���3��}��I�����ɸ��3��v���>�I8��zZ��a�e#ߏ���	�f�<6��L��j����~tj#a^+E��'m�.%%51���m^�,���L�8����đ�x���p���F$!���аB�v�mk)\@��.�X��I�5aүq������إ��n�&��)f��7�����ĀDb�3����|ɗ�a��������V������[\�i��>��e��PY���?Y��#V���8�����v˟�a�5 �<T�h�PBp�Qլ�y��K��r�ߵ�C���a��	��
�T�XS���dč�(��^?-=!�c���//@�[�|YY[Rō��}!PD�@��+t��MV�Ww؇���b��s�x��?S�
�9�~��{w�X�@m������[���0��'�����4��T�����Bj_t�m?/U�33�>e���LO���`������������#��Sqa�HUK
(5	���XY�z꿄!Q��h$����la~n��������q���	���-�JE%%1#2��u����^:e2�)?�ݯ��	����i�Qױ�PA���'����3ǩW�`�S�[9��ķ�;��Rff��#6���tC��!5�y��He�߽;�$�����2��g�χ$�*)����h�2WwͿz�8�EAI���`�I\=���ď����(����}�Y2���%J�c��^� ��ar����w���cUh{g'w �crb�O��BM1J��E���д{�(��F+j�N��5�z�l��,!Rٕ���-��^|{.�o^G_��Lj#<Y����\!��dk����qL��:8D
jj��I.��jͲ41y���rz�,T�5�(�5�j�c��ؘ�B�%^j��g��w�+��i"V�i����r�s������z'݉D���{M��◨��^�C����bc��I������Ѿ����˂Y[��afR��]��e2�g��̿��9! ���P���n���/�z|�VE)f���3!�27���/±_a�4����%��}�)�V��g�F��6[�)��i�鵛g�P&s�5����,�G�)��g,t�hh��b��!m���$	2�6����Υc�S�O���������XJB.��Z$.]�".���}\"�)��4rq��Έ��*�-���u5@Y� �.k�fV�,U�0����L�h���.�ߐ�P1TZ�ښHY>��5��/jֳa<0��}���F�w����j��b���3 ���^%����d�p�ڞu?d}���%/?���p�C����)�D�s���m��q����f���t�}��GA\�WЂ�V��a��jbb)qO[(d���֮�e�!ȁ1�xiDBa�>?uzvpӏ̯�~��Ջ���-ſ�mN[���f
�ԟ�OT��-O�'q�bϕ��n@�t4��1~�h��ө�l�\�UW�9�W��!��+�?V�|ݎ�6)	#o�<--MEM�~^j("�eFyI�ͯÍ�~r������nn�L�:���!A�れ�o�4Ȯ����G?�ݯ�Gۦ���3	���>�OpXnn�)�z`�h��E:�S����� �����10a^�
,j�9 ��������;2RO��*�2E�1�|�(k�ŪRد��b�,,�Emm]��9��C�y����>���	3�<B�K�{k�:�\dD� )�D=kq���W*�j�e%%����w0����w��6L�=��ԣw[SĚ*��� ݞ��v:��G�Y������m��Q���y��<�v�xA�wA^�H�a�_� LZe�l�8�EX��ֹB�:��u�QD�퇭C�Yl��*���qL������*�q��^=#����2?��͏��Q�wY.�X�:b�$�����x�d�Ų�m�R�����w�&l,��G�m���X.{`�p�p�3]c6������Z������t�������_�"���������mξ��ێr~�twX����I��(+s7sy�,������Heg��gߍ��[.��XǷ���ل���ܾ;����<��6ʥ� �*2�H�b�Q��b ���?]��;N�������U\Y*��h��� �(/���h����� #)�

��935��
�I9�fff�E� �e�Ѥp�X������ђ^��E_ѵqa����+�7� �H%F$\pg�%$u	��W�h%��MK2gsI-�0jǓ+x_2����q�r]�[5b�������r�`��*��
;��1���i����2,͞߿b�����ӕ����)i�}]����3
8���d����yL�b�V_p�����rq���7{5�{8_��D��	U��K(hh��Ʌ��2�
B�=og�o��>?d%3K��i��Cj�lVRü�Ӓ2��be%�����v� ���{.���-,.���7(�d]���]�G��_ގؿ���wX_iPy020d�Ԡ~����M�>P�|����Ӛ��^�fo�А���V*�گ��sB߿�U�<�����E�<�b����!-+i�^3,]A$�<6n)s+����V�P�?��g��]i*�v `|C�&�|�6��8Z�����3b
�g�'D��!���>c������Jg�I�A����Y 2 �,�؜S����5�|<ᣃ�'U&#e~uqA����o�)l���(6!��jw����h����cMY�|5��SB67��Fl�:e�����C��߱������flg�&x���ó�k�nη\��I��C���|yB��h9�Ь���[R�P2��
y�Oq>�Z�����6�6��LV�=��h�捥��۲>�ь%N&#�4�
EH���$��ן�Z'������F�4s�
4Q�7��[&�Ƅ�;N����^��@Z���R��;%I�����f��g��<�'!��(40���|c��,�o�^��rk�$Q��v�9����}�4��IkN�x��N����������u�b�N���O�y��E٭��'&��n1e�ǣ���J@`�\QՄ��۲��S��Y&i�I9']A}������BF�j#��_u�v���N�7g��'Q�؛UԨ�����Zg���?��=%~288�Ң�7I"�L���!�.�x���'�!�3jCCC2���˿��2��8�8��q��сK����&%�i�������B�����8�$p�7M4geeu^6�j`�ᆛ�t�gw<+Lo%"�i�R �i(4���s�3���f3�c�ّH�}_ߒ̄��7�1�6���-v�hb.�%�OvU-R�FJK;�M�|�~k�4�ܳ��\�ʘ�R�η\�bM��3bZ����Ϧ���+b��c�_�8���ȃ ��{IHLLRԳ�w���͕�� i�>[@����c�2�I}��K�x��ᦗ:3�����0�hkg��G6�L�M��J
«�sʹ��t�O1���GD^��o�a%������3����� t����}�-�(�%Y�ߥ��W'��AA�U�.^XT�j���իW�_��f��l�jw����^B~��^�k❀$�������!E�)�`SK�ł�YP-�Bn�X�	XW���hN���?���$s�����F��k�2rik�s+ww���8��H<�	�����i:o_߃"ݾ^�?i�f;;�g���&&�J�w݀�)M� /*TL�OL��%�t�I�rN����Ͳ6���4���ȧ���Em���0FLL8��Ko̤�tƗLZ�}@Ȥ�5?pӢZ��(+,�J���6�=A(-+C���Q�
��-��۸���(cG5�����;������6�S������(�d9ˑ����l�����x+/���Y[�c�4ݙ��.{G��n]�"���g��3��w������@2��g�)��5[c#��� ܆K�MqJ�n������>��I|o{���7�]\��<�9�L���71��	
ƅ�mN$W_}���)Y�|�l''�JR����������7O�H����~|k����� �޴d�o�7ۨuh:��u�v����jɶL��)ͺq��3��=��iFt�����?_�'n�v�����B��J��n�GtB
��*�ˡ$�\���j4�;��};@�M������Ϻ~���Ç8�����RM��)�$|}VY�7�#3s{R]
N�������"$�,<<)�X�o�%.�a�BI�ȓ���˝Q�p_�'Zt�[v�A����o�dn^�KC�|�,u�;*XĂ�<�K���;���Σ��N�-��K���v&���ZZ�x���6Z��Y?w�lH��mmm㓓C�׍���͎6�m�����9����c����Ot�ޗ�����λ�b�A@����t����[�(�?^HI�4���|/���=��xc}]��L����E�&�|'���Sh<�f��B%�.B�Fn�ހ�
W�%>�b��7��b[�/�#N�z���Ғy�Ч�7�I�kl�&r`�Pb�c��p�RE&�M�)1-bLJ�@��&G͟����!��
���V��H�S_[+��;vL��n9]<~���ZFY>�!&f�Ti�a9���O=��*_����D�]p��T������a�p	K�"��!��m��(kjxy#zu�6���k��d �0b���l�Nb�0ɓ|4�
;;����5*��I��r��D��v�E���>#�~�TFN)���`f+2*3���Q�0�R�~uMMȰ3v� /?)	�]��b�R(�t8xlƤfY�����µ�+��{���)%%$GN.S�	�G, ����hs�𐕇�+�p핐̫�UJ*-z�??gʗ�T����r�;2�������d�C��ܜ2�a�a"���+`��/a_�L �<B_jzjc됼!O^y�����^�����yxl*?��6��oYi�������hACx���xICx���j&:��B�ß:��+)��I�t��ݭ�4���
o�;;�߫��S��*����b�5)��oav���q��蝉�,,l~	ܦ3���~���~�푝���F�÷�{�֏�S++1GG�˶�I����g�Mt;I�[,,,���涔��L�?������x��ǈ�G�����CE��n��S%�tEC�ds���m�h��q3@:�#"��,V2��.0܈��Oiw01ӭ��LD�:������~�g/4��=�qpg��-Ю��Ɂ*�˘A����C���ͰLN�g/�J������	�y_F����pX�$���;���7���h�}���>h/#�m*�/���"����YH@����s�������p�~�j�;��υ��^5>�T|�*�	��i#C�)�(���֎1��9p,7��]�4��C�����;%PF�T�3�r[���\���mc!,0�>y����?o�V:��{�j�
(I<=9q4����˃~x��6N���t���,�T��J}��/���R�R���Ж_�J(cbb�T6b�B��ېQyN#A�&�׃����_��[;8̪��N�9Pr��LM��S)��»�qX��IF'0N-ME"FD�$��%�V��������q���3�"�����!?�Ώq�=�<��67�F��o8XX<��֮P��ʎ!����h:���*�0�5�/.�'��#K���-2� ���n����&U�p�g�m�����1��*}�*�����~~y����d~b<zzz�)\���5:)�^L����M�^�YJ�9����o��s�ٳ98yzz�c�m\{Bur��	u1��dll��� ��ߦs;��P��`����&fd��9�̛i"_ز�ʄ��:ͦ� 	Ȥ��x��2�%ҥZ\Cu�pH	YY�vּ ���ŝ�ԑ��碠ڼ�]Q�ٯ �'هGQ�����a���1I^E%�u155U&Zy"J����Ɇ�/_yEE�ct6��M�o�>��Nu��e�Հ�D�n������*#�K?���2\�//�������o�tT�.��_����e�&�L����(Y�(1]n�}.Y��BDU��h~֋�6�"6eR�뚡�v^^�.�/ĺ�#���������+y�e_#�$$�r����ސ}�L�~SYW��̷V8��r�S����߸�=<@L����Iz���}�E��^Q��C���Ɨ�\e(h�4�t����4̀�,��W���++U�S�_�O�
'	���D!"�M�Uc�K SRb��4/f�c?u$	H��,�����-�\Q8S9|\�N�[���A���3v�k���v\q�	��#..��~8_y�$�����կ�e}MM��9I۶�?����c^u��~�GJS'��x���c���(����zt�����<D��s��剋O����c;��A�y�|��a �O���sp�	)�O�b�{G[�h%�!J�--��P��>��������ӪĎ�\�HQ�\#i&=���bp)�1�\֥)�6D!?w��N�ET�8{�ޛ�_<ݔ�KD��G�5���	��v�r���>P:��l����bM��.����*���Q#��tZ��Qߝ�:�����RPQܑ����rU�>2N�#M��6�ѫ������00H�+ �z�5MM�m��J|)��٪6��Z+�nI�W�5nt�"~=���^�:�*4_��GE�����^��k�b���
��8�[��+�6`��jpSTD^�$	Я%�-���� Q��V`�T?~��^����AE����`�`��@��P�S�	��RWW��'A��QH�p{��T��"&%�\���&>w��)�b_ ��������NZ��W�=�#5�%d#@l�G�� ���\�e��f�(�� 4>}x������$'8pw�?V�ё)-=�#��ǯ_�jrl���7��>�}����������$�S��������(~������A���њ�Vff�����Y��R��Tq�t,7�� w�mT<`	��`i�Sj�R9z�'��ZZd��ؤPO�>͘����m*�K����^U��6{A��\���	~�21��)-��u�$��C*2�RS]=(��Ö���Μ�b����Q`gHW'+⢁'J�S0\���ss� ��{ڇ?�4>;;K
V�cb��9�_Z~��j`��Yw�K����� ��Ii_�I��r��\Ձg�x����ږ@���1N,�
!���:Q�f�/�ݕ3X����m=U�����@Ǡ�&��Xx{uj6py|�ӹ�7�o�W��%� �n��KoŒ�2��ڞ�����(lk#�LP-.-�26/� m��{���h��J�ݬ�\�]os���pp%]`%W�~<�7O[V)�w�g��c���9�Ҟ�TC<��IC�%%���@ 0?Z��]���;ri�n�zj*,!,;;{� ?��;c��R�sD����^�:���X�|��3F�¶O�9��I�8�Ϙ�N�VT`�I�Ꮦ:����S��i����Ԟ�S5 �b	�3;Y��⇹����	eC״i�.��&�nO����}d�+-�#}�Rcg�
�T]�B���5��K���G�d)���������-��F�"��) H��lyD�Hc�V�t��+�FԺ�N� �T��O���T��������_����.�+D�*��o�;�=�PXM�a��u����İ7�J��	��Ȅ|�MM{�.I����N��yb�ُ�%dj 4�p9
v���
 |�{�(|m��{�:S%rrr�T$|tS���0�I�}=ؖ���88N���y:0��4C��'Q\Fv��"�p<�3d����HnV��r�7��NW�vӝ��E%��2!�ߜ"Qѩ�]��N��(@�dd1�GK�]����^�ŕ76b��� ��C��◊����U���vK�B���k^��QS�ws�]�]�(b7��f|�p�a���ي���5�3Dt��RJ�<7�����V����#^��D����)�����և��!�ԳP�=�E�����1�_�J��C �AM��ǀ	�^��wD���h��c�4��c��<G���Ev9MM�cj��B��ΟQ>�Ǒ	n�n?�� ��DA''Sy�ݢ�~r%�o" �9�����XCC#�Nph�a�����(�@�#�65I���-/���]�K]�9���!��g������b�2�.Z�wD+**xnvU����f�Y=�u��z��jRԇ����
Iww���!AJJJ:�w$������z4���/�#��=���~]�@u�����;����P�5.ݛ�����]Q��f��L֟���F�T�l,C�"dP���MWwV,_���@o�HB]�AD�48�_Z���[��ᅑ,�;�) Y�P��n{�M헢�|�.���?=������p~%�x��&�b�+�hi��֚��*-��E%@�Hz{����(�e���ٓ�p�6�����o'�����R������a*ŧļ���S;���$������� ����ڬKY������¯N�4��q��~���8\>��C.��G���q?v��?	�G�����~���?~��kk���'*]��/Sm4�0�d�i������N.,��t�f+�m����+Sx�vF��d��)�ǧ�gg���^î��4juz��q���9����o޼IM����
�m������� ��:9-F
<�'�h��|u/!�_^^f����:��I��V[F�.d��ߥngV������%9�2�0���|DF�@HO�^1M������Lp�.�*hXXX�q5u!"$"Jc����<b+BmV�� �ARZ���X$@���D<<8ar6����.��ӿ�CA"{�m�)��N!�����Nx��"�;�B~eH���[rZJݣ�<���/�o^�L� ���RX���)%O��K��a=]e��ԕ��V��,}!r0�k?to_YA�c��i�&&��yfB��-��!KJފ���u��a߭�Z��t��h-#,D��O��I��r���?\G��� B�C��ov���8�Љ��v�۷"itS���5��lk�� yu�1?k���s"��I�:�������M�yrffe���0��i���F��jk�Sj�\ �jg~��9	��Kց�鄌��ȃ��H�f�����J��
b\�:���z>W�t�02p#0PD�����y��E�T� #��iQ��� ��BZp�;��6uq�.'`�2J�bRd�v�3��:�*��%���`�j%t����Y�X�3E��]c2���Z�M���mu�p~���b)�Lm����X!:�����5�8��0�_e��`'8S��G�-����Y��m�"K��,�=1�|��`�oG?55���xg>���6�SV�Oޚ�I[[:`�8�Vk��ƀ&�=�&��Ѕe�n
<I.�f�%��qߢTI?�}�陟OA~�W�(��������!a�y��n�où���L�RgQ>����~������8=�t�~}�9�cr;��;��:�4�C�Mݐ'����Q�NX�l� NOaq��5�0�6җbl��g�q��V����d�3.��s��՛ig���㭠��DV�O<�@;y�`���@4��
��3FffiS?�ζ�����`�A���WL���K̭��̖đM�kXXX�~.<��4��4�7�Q#�����KLL1�g�&�-yEy3<�������]�t�,&&Ff)>�����-������
�|�:�����|�
²N�c�Bl�@�V��ڡv�w; F�>	�����
�*S��'c+ӌW�
�{����п�Z�Y�>שq�i`�p#?��b�a����Ib��xp��0p�g(KN��"�q�:U�T��':�LL���I2�}<�iZ����3���1k����l���8���G����+D��,?q��>;�&�*�x��LBDH��E�I��
A�#��p�rdU��H�I����ڊ:.$�:�})K�AywuXՀ�z���Lb�_�������m����t���vvv@�KQZ�p!>>��W9�{rۏv�����d��ۯ� ���sW�M���VY�t�� �3� �I�vw�QPS��k%>'�V B.�+������P��y.�4���E��� j�v��da:t5����C �(����"9������.��Bo�� �;���2��D�O����j+f����6RRRN֍.A����M�ֺSkB��˓`�)d\㾯�j�p��R��N���SLkt��~�$E�`ӷ3��\p��|�5��(�Ե�� +���06_��{���A��-2���w��➫Eo��Xٳ��'
.gMk�f���]h�-�X�^Etp���w�/Z����kӱ��Yhƨ���_��Y1�������{��{mh��a.���J�@������R�g> {ɅXEva��~M�;��Q���Y��s��β2xb�kR�sC�9�p��QQh~�(n�4���ʊ���sb���Cxtdp��Z~V�v������8%��\%jz�}6��}�i���������FG��$p�߱_�ߞv̫����l�U��(ʊjZ$�@O��SQA�u[���ީ�p���/W�d~_���B��v�+�Ht�h j��?��칰���-6����`z�Q8���Cj���#Vĉ������n	�
ۖ�2��b������=o�v��w�����[\v>�|4
��$��;'[)'������K�>������xlf���ǌ?��
 ���%
���P11)w�Ea'�O 	`�@�Z�t�;�C����݇}����xs�y��������o�D��}�����eЁ�]�����=��T��Iu�q_Za�
�i&i���v�%QGtv
�IJu3��=!�q~���7%˓�^j)��ܾ�[�ý����5���Λ�5�	|�����0s�׷��
���6���n�Ta�J.u�S��Aq�����S),�`��MF����ޗ����\F�F���l��o��!,WH?��D���KH��@FZT�S���M�1;:B\���l��"�6��)�1(��"e%%�b~���cPL�/G�?<�5;+��ȍNM��D��-����K��s�Ga1w��[��c�'�9�Ε��n�-�:�.������̮�X�B�ʊz��� �2���o
�k�)L,,2q����sK� ��WV#�P�l�����������zf���*rR!��`E]�4@e	#�7��M��X���
�����ϕz�A$���(�He�& Hx�~K��������C��%eˎ�'��/���Z�ՃW�u��>�\�����S������⢉�!!d��GG�a�~�yo.����_�� <������%��f�)��ѿG�^�*�_B�N�?�j1�:����/�(M|-���P����l��o�o�i�=���^�ݝ  �Cy�����$��>"LOD^��}�����t�t����;O��ƍ4�؝��98<&B�%[4��0�hpxTR�}��^�7}mml666cSS��-��2
��ѱ��ؙ���!���rS���ͯ���X��d4��+++�Cc]�R0�^LJq�C��ժ���Jʋ�;����F��Ս�s�E�Ԡ��oݵ��܊��T��}("Q�`A ,d<?�o�OޤUt\�6�S�Ϛ��9D\~��ɩ�����c253���27�ˉ�5VTT��3	���ym�������.�l��Ëvu��/%v��@%�98���[,�H9���5!�#�'�l++1�����`�=��-"[+V���J�d�5��JCC��������Cҟl�=!
��������������"�D��A�e���pT�jGF��"P�!d
�@E���6݌���>��������L��zVvs�η��?�=�oM멿�|��ԯ<i�������b`�t���M�͍���uq����O�:���SRx��ׯ�> ��^�f�2�A 7��,<vv_:�{��B��fd|
���ۿ��~NAE�7�£rP �%y�( =������k����޿G���E��s��B��$�����߯�Y[�!,o��ׯ(�1��t�8555�~�
'�	z�����gl�gϓ���h=~vH�&��ڠ�O ��x�2��ϧ�tC5�8��~}����ؗ�P__O�J�j����P'��>[��-,��bH����@�_eNJA�[�!����d X��;
��;���j�L_nRt��]�!�ܟ-k��B��{/��nl��A��
�)ꅑ? U���r� ���Z4��|���^nl�	Iik��\;�v�Ta�.%��M���EQ�zKR�Gx���w���Z�ݽ�7�?G���������e�b�AƢ��a��D.'m���tvv%��F����W�������ހe���IomB�x���[����bT��K��X�ͤ����45J�b���^?(2�7�����W����C!���Zp��#�y0�E����B��&';�%Z=�K�qJ"�`����)@�Y�[�^p6�: k�HH��p�p(��Q��|�<�v�p��x@�n ��@~�u�ݦ��VU��*+L����������#~�/�!�����X����^��f�o����Y/4���������Bhd�a\[� 䚹#��	��լ��^'˓���~�(B���d�����DH@Jd�\g����VlV\��.'˼�}[�6;LKK��<����7��( n�	noN������ٔƧ�GML� l��$˨����\�Cr��o����!·�����#���%��{Q<����v�c���Gm
t�uX�TR^,bd$u�6�/%�\���ɹ��c����9/��� ЏY;9���^W7�O�6p6��dO�ٔ�0�$�fAXS3d�Z���s$|�4��خ�ax������T����mQʮi?z��~��7r�����M78�s�O���I�z���A$Isc��±���r7��:��ؾU�<NY��P�_h����3�@��jż;�9p���1����Zg����=L����B-Ǻ���u�d_F�߆8���� �T�f>�$G��g��fAŹ�����@�B6���޽�ơ�7��nB�v{a8G<쌋��w�'�1�o*`mMNk����nR��mniIFCW���9`l|��E�5�T�'��\�i�a����mj薌2����H�Q���cf@���N㰚�]k�?>^���wp��چ�>@!����Uꙸ��o��%�/j�Y-f�@�7�4��j��Cj*�`.�'II}�Yobo�N��fn�����Rv��ޭ,��A@ן<�}�{������rMb�y���E���,�0ǉ��I3��ݬ%$q��E{���&8��	@B�h��LB,&#��h�ݱ�a[~��˅�TXx�YO���Ɉq�{���H�q�`�^�B�AX����K��[^J9T"��}�B;~�
t���k�1Th^��lRF�����Ez�.)�Q��AB��MC�h��+��|Y 9!���p��\�F'iy�(�����ݍ>���ޢ�R;�M�:����0`AXtn	��Sg�!��f>X�nJj��PY�^��ٲ�i�(��� z���c�VP�y�C��Oo���y��?��}Y����v�eҺ��]��Q �%#�O/����1�>~~�~�����3J�]WV��d�3M����VnnB�Ģ'��]��i�X>��뀠 hHw��'�R�@����_�I��|�or�)-�344��G�	lj�MC�>\;m�4]CSs�ހ������xp�Tn����0)99/���d��o?o_�w�)E��[-�^� 𣅅ɀ5Z5���V�x2���%%���]�m��女���@_�ô�tU��1��,������&Gn���ps���F�u�+++����a��/�ڊI��.}��=�#�������������ȃR��3�BX'bb���S���\S�q��������ߊ���YY���}�k2}�p�6K�����g/��KH��j������؃y�?�fh���Mx�9��"���V�:T�mB?���n����˗'!!!�U��\˂�&6&/��=	}ڑ���ks�rN�<6ν�..���)�bc����K'Zb�w{fG�:"�\�7m�4��7���onm��_Y������y�wpp�P�����ގ��I�ڡ���Ғ��;�$5uf���򶸢L\צdd���UT��m�@j�GYSk�p���@�/���[v(\����:::{}����	NNNX8�4��r��urޤ�M���5�g�\A\���M�����olj����S����|����g>�~\�����������M�?/�����K�!=���J&`Nzw��Dq/���pM�	�NW%ump����}����ֵ������k)!1���'���=�2rK�g���2�R�"n�0hff�����k�󕯤-$C��998�씭ht�o6{��}�O�AB�����k��"w=]L2���oҸL{o���T^���t�B����R���TP��]�!��@�dWOG�{tV3���?T
"�Nve���K\�e�ߵ�-w��[TU�K'<8�'+*�~���ᶅ�����H�%�:����O��a��|�dH�>�rkQ����<��e�5M��筻��׍1�U��h}r7����ZN��!5044$䌨]���8nE��7����4��P������^^�CW����_�'ff����[>�LuC@Ǫ����oJ~N�%�(~��<��O��[M]]O�IOR�"�Q�~M�Z���Fu]��u&c�5��6��C:MWw��-��Yox`���ȵ:��MP�Y������_ �'���ƭaKK��#��ׯ�.�Ay�O��~�k�e������.\���4d�`y�D��������洀?�7pr�f��*�H��5�6�*�Rd����d�n�b��z�>�'
�i��%�gZծ�7NN����vv�A�JZ:��t8���7�s+]��U�Ύ%0Ud1l\|���U���֔��Û�H�-n/<<�ڳb���ty��o)#AO�{���[���ꫠ����L��|U���: ��/�`~��ˢ�:�C�Z.	y�ϲg���$�O��(�>���I���tr��{�d��j��4x*wkOO����w�Z�Hb����[�E���è�  ݝ�ݡ��t�4,��*�R� �%�%��Jww�K��>�﹞?���Ù�����=sn�3U dRY�H=S������J���o����{�xH����h�����u�Sq�0����\?�d������%34���_,' ��ei0)))���4�ٱ����S��a�-��h�2��99q��~8��L������YN%"TD/���O'k2���l@9����ӈ������c>��
|x��ks�]b�1}�B�F� T��)���6����MW
p*���E{;I�˒)3�tC�� Q�.�� g>qjoi�[�QS_�������9�@�h�(6.iT��mS 9��]wώV�ѭ�=����'Mm�͸�@pnP�֊����U^�����Y�Y#�ǧ��	��[?:����"�~�Ʃ��d���Pu�1��&�}��X������y���Ay&�}�?3�zl���*:����а�-.���~�6�`��~�
lfaI\�p�V4��iGF�����W��0KI�MLJo0wF�3=	�B��{Ft��66hf]��@��=ȥ�vvv5��q���=���CW4 �/�d%�� )����_�������A��怽K�0�����U�FJ��Hs���梩�@�d+ς��I�\	М� ����f�� �~������~�1�)P�Zm�8��j7b�[����h� r�ѯ�w+z`c[��9�����c��F�[f&Z��J*�|�#��_���"����b�_B�n�,���5y�#b,���yR�� O�XU���Uc��V��p&LN�kc��zT�����-�}>9��D�p,��0���viN���
�2 c�=��o�o��f�V�???�ygP�	�d����zq����y׮ˏ�������� ipFZ���'t.�nD'�!�U1"�����J}���u41O��4@�c�cCҒ~m�|��^�gҵ���߳I���z `������<�c����u�%<_�66�����g���7�v�}��5S�o��Pu��>-v\�&x QY,�2�W��>�`�ޅi["�]D$$���/<����ۯ�[�o[II�Ք����V��$� 23�R$5��(��a���ܕW��\�G�ĜOs�]$2/� ?	&�E �m�୰Y�Q�R��JuUU��A+_�������1_��@��+�������oG���,yXQ`>`	Fp��+Q�J�^>[��˫In�-���t'sߊ�#	�l�7���+Z8����2=N��m�Ł�9ڨ�[�����!�T�7��`��h��B��fY�cnI���.סQ��qeii�3�j�ᥓE��Pc3��K[���n�[O��7>5g�X�|x
���x���5i�(}K��O�2l����a��c��Ӓв�f#
�LL�~����O�f�,�hb�^�&���'V��Z����=ɦ�+���F���O�˽qf�UO��5G��ەv�Ťљ�Y�=��'����k��2Pmһ��BY����?�knN�d~k�x��s�O&���/`���1������E'm�
�V��X��ӭy������ד/��{B�J�K���߽~�텋g�Y�<�7��ן��PQQ���E�a�s#R�?�0cF�I��I��cccsȾ��A�+����
���; Z�6��T��˧b�V�s��J���Q��^�(�5��8�++�$}씼B��' ���!�כ���-���>�^ns/�K�')(,|����r�
����gS���[?8���2�UVN����c�wTx!f���"�߭q��i}�}Ğ��Ȁ����}Z���$�ԤC�Pq
�4
Һ�O��'����i��#�������;&VV��D�u\��Po�R���nZ/����-9�#�sD�ĄZ�����$1���#MfV��S `G���~4cψ�3���;9���%� ::!;ӥp���oy�����eP̎��[�?�xO��߷��TQHx��,�ɨ�7F0��g�~�B�zPC�'䇇<�q��l\ �����ݐLL�m����s�a&u�gXg����[G>���Fӭ�x�玣}��Λ�u���i!���k�����dce��2�:I�(|�1<�6�_��hyL�Ƞ�G�A�P_8�����������u���$"Nӵ���J���!0��yq` ���_��r��E�/X�֕�zc0hhh���C2��곍 �QS�VWv�u��il4��~�ɨ��rly)f�� �7{#p
���0O[�4NS�}��2����H����ƵOBjj�߮�����b'i�9�tJ6Mju���?�襏XS!cH��0�ǒ��toho%�UH(����4�����C5
Ī��h�#�����ߢl�B�y<1R5̞���������ell���1�1<bnn�xbk��i=�;�'33�3��+��o�i��0*'P��|,�РE�>�~�eyH�$�^�=;o_`�5:�Au\~7g�U�<憭DDDT���K�Z16��]	Y�W������T��\ d~��6?�ti���H��ga� �:Y�U���JՄk?m���s��1�)?&�l���8�?�\���%�K:FR�`Vd$�z�bOz�-�^�`��9*�W��Niq��* �#�#�	ޏ)mmg71$�@ ����Q�Aq�4�h��ڣ��+#
KL�eP�WOK����҆
�	4d;TSWWWH|�����ɝ�v�����b!ѯ�����m���;��vF�h�������ɝ|�*��-�WBC?�m��VA��ވ����4%%%�������<<�b �!�ݵ�Y#�a<A@M ��	�IDtܐ�Y;�lQ�R��&L/��!H��M�df �GgJxV��b�	h�ExCD�CP3FC��)R�z	ǜ�m.���:���|��ab^�� Ep��G�Wf�^�,r*�R,�O�̽P�oS�b122&gA�!x)_��םor���߅:)�u��z��(�Z�)o2E����	D𒐐09�T�����-Q���ۖ~�$ʄD�����߶�]A(fS%�D�.�����Y@�ayby��ƻ�!"#o<<�tL&-��q�mZ�Xs�UM������g2@(�Ԩ���-���^�С$��q�z;7) ���}7�>45�a��^1fp:�|���vF��8���ٛ��Ԓ�w��	�֮7xMing]H�|��qr�h�59�ܬ�g7�ލ�(
KG������ո.˙�>��VU�/�;c�dkF6y�<g&���i���E뭝��xl�|���j2��y /XM��F������Lf?��h���Z�u��C�����iŗ�W�?���U�J���HN��qpe%�߯Z ϴ;3�B�FU�v �T��aT@�B/�إ2��{ʸ�Fd2����'�p�5���lVTTL�$��}�ԫ��ϯ:*���W9?�����&�$�jx�ʺ�_y3�UXz�g���|�1x����~�ޅ�tk?�*~N�{�X��1I�R����O�@�#nɬp����0lJ�y[M���T����>�����A �k�]�Fl�	����ѓ��������zj12�����Y� ���Z�}����ٱa���_���A'��y�Z����m�00:&֥קrޥ>��6Ϫ����6��.��+��/�
�Ɵ㷟f;�+*�G#�ڬ#��)?���	
��OQ̎��py�4g󌔞�NT���8;hǟ���1a1<%�>��DV�Um��Ic�@�dW�x���z_i����b��5�������U�����皘����J��DYYYkؙ��a�����N�G��1���*��q�4��A��!�A~�oD���A9-��,�V'��<��%����0���F-����y��_�j�psS���s���N(�����wsvrc� �AF1�ů
&�- �p�?�R��+.֋��ZX 8Ʀuumm�k�]a-��87��ނ�Y�����H�{g[�ty�'�8�7�aM_�~{[�#���@z�
3��s�b4Y#E�ߵh	5��tw����1��Q3o����C���7��E_U&xs=^�rZ����!Z�cz�fǲTw^8��T:��4����:o�M�Pbq���XX�ƒK���fx�a�4@����_\;6���+��HӖ���_py�}����Z�	� s�A��|���VͅπR_[/]�e�}S8��⭥�63ӑ�vLN�i{���ӳ.�Z���!S�@2��e�dl�+�ܞ-�{Վ���:e��BC�����GP�m�A�����mER�0p������k $QR2�qF��|h+���p�4�9�w�2?�3
͉σ���z܊���R�^�=2��j!�Fn�R��}���F��]Ԟ��j�83���`��4�����_�Tkiy��ܽ /�@ۅ(�69w?'� e�o$-�`xh���%`�'|����?��[X]�������mij�bb��=GDBf٨����q6+Mh�xx�협D�uO$��h��p��^�OkN�D�1�(_�:���,��;��}q=GsK�'��?1��I���&+���.�Qh��x/e
��U��e>2i6���T���ۢ��8Y\.���u.7�Z���Q�JAAA�_�D��{��&}C8���{S:`J
�3�J�Y��"�� yy�ɎS�O#���~�
mې0 �*W��|dg,�/�Cl8�] ���h��
�0�V������A�]�J'�?�����!���[�Ε��?���䌖�m-����u���Ù�����=�����*̈́���C69'��c��Z�x9O��#��R�D��N�3�Ǳ,�s�C�?��v�����@�·���||l
�KPc�}aG�B�j�~��恏WU�F��y�>�WV�‱�y~|��ް.�c�>SA%0�n�P�&i9���N��"�0x1�c�֎���9����NxS쓷ƑG�C��nc�[ÿ��f�NJa:���Sܜ��'xb]�6! /�&���Ma��S��ݺ�� �\��0� �1v�DK�ۜ�����]f�p������U�;��,r���u,~2;�Y���I9��ccJG�vq�8�
۷�����*�Y����]x��Y�O���%�0@D�Ku7GW�����Q�\b�N�52E������VҜ�'��=M���X�� vhS<�S�fd7�}�X�	ɼl�u.�q"Q~	J�E�0�����eMCG��MzL[��[
�����KA߂������d9j�]]'�<�|��'��C���+g`7��F���xf�����G�k�ߴ��%T�zjk��_��0L][�/�zEFERl��Wͼ~�uM\~�����.�Nw�[�����e������V�����ھ^>%��ż=��qT��_�m`��V-�װ} �<W�O�L�dc����7]��.�:����[~⠅���:��� ��x��,���ot�y4_G�z6�����C��gL���"��*pm %筈��3�ۘ���j��}���3'�$-�/����'Bi�d���'慦���
~��^[�zJ.fgZ�������Nj�������l �U��MY&��2�������c�)�i_~�������H>U���V�ue$�����P}x��&89�����=*�F�f��g2{}C�X\b��fu�u��UI�~�I�;��]�G'th�Ͼ���B��j�5�v
i��G}�c�"���#����@#D�����ݎ�O��ݒ!f6�چ}L��:zz_�3��s_�"~~�4
��G��4���j�C��R?��}���쯕N_�1�[�Q ;dcdD�"d�~�j�JT^խ�t����իW�Y���z��-�`����©�4Q��q�j}q���:������-�m�gM-��_��^I�җ�A�+1�9)�.;��OH��4�f��g�q�XM����~546n�
����UTVv�JAf�c+Jv��ܝ	��W�ܸ�JGG1��������|������[���1q%�g,�N�N9�'d-���A�m���nN��<<8��������U7��st�$�#�çܻ�蜦����E��^1����_���`4�~�����p�)baa)d��><�l��/B�)��������N�̜�qWW��@�n�S��3%h$uܲ��l�K�����>W��{h�5���AE��%�����r� �#��i��i���۠:l�G@ ��,�,q|��HN�vo;nO?��I��Y��� �T�ϻ?VNVZ�66X�=��҂�:�.��1������xn1o:s���D��8d��r�>���?�P ��͖U��w"��Eq%V��c7��a�B9 �q�IcɄ&&U�6d|\�v�ˏ@�f<�4bl������B��~27�Ce��~���[Ef2q��b��@�f�>=\l�+�@,sJ�Wz���ޞ]^tGh |�c>f;={U���r���?A/�G����X_o)z����1���z�G=�	����̗�������?���^r|Q��y��{�!(��Ůf�F��隐�����2AE;���5ZkH��Xj3���k�D�\}����,č����x����qr�|�l��1;�r�ĉ��7�����/�d��d���4G�O��[�n�c6՛M��K��T-�F��L��FKR,�������MM $�H�u,��ؼ�q=c4)V���\N
qE]����~"� ����1����{8���W��n�b�k0ך�ZƎ�E����v~���B\%��,�^r;��@B�d�ޥC+�.ʏxx�q���Z���B���=49[-T�N�/����x�����t�ƶyz{ݜ��E���Xli�}�h�ҝ.�ll@^�k�"!i��:�p���6���v��"���6f�G>������R�Y'���&��:s���<��ӄ��YJR��ĖB[�m�Ll�e��~�̿�_�Og�
p�<x��L%'��\�����VnLM]��l.L�?QӰ�7
\_j�+1Z%�ǧ�OMO3y>���<ٝ��t>�aK��g����HorJ�;���v���/H�`3k�~}�Bۛ���t�[���H���:�ퟚ��s7"����Ld�!��H�k3���+R�1�ax��.S�Ү>���i��>>5����]�S(���T[[+�ˠ��@U��(($�l��!�+�B�E����I�cl��7cׁ�Oa�0@��%���I��I�842�;�Z��fꏮ����2R��43n�7���s}g蘬��3����偷H�a��Yh�o�5*��6;\n�؍Zz�Ņ�d��#3�d���пR����%��ϲg��d�BV����S��4x�g�˵�Øz�	GFF�-.��TC;$7��v<5�!���C�}V��x�����F�hz�^������W�h��{)ă�r�I��߿/2��͒�5>�Œ�����i+*�L������(c\X �g;��׹b{����J0�9c�T[V�����P�o�5�v;�b��DiWy�<կ�є���j���`��bHJ@9�]�Yj�4���)�A�/�˞�|�����Z�����f�1dL䟆������1���[�Rwk�̑VǲT˵ؔ�W�Hvc�\�[q��D<��/,�-K�E�3��|a�,Oj��~��hQ�_Z=0V�����²�9[3�	f;{�q<��������I��!ss�$�����iks�[[[^@'��WF��ģ~��8�PS			H���Y]�:CSN�xy]�)��o:�����ZF��^��Ȉ���}9ܚ�>X� �j�f�ѕ��_V�d�'����˞��s����q� nA���xI��D�iV��j�����q4��P������;&�T/�Y�!f)��G�2�
FQߢ:��}wXd?;�Z�l/��<<�+��]ʇHm�Bw��˝��:O���K;�!c��o�cߑW0�t{�_O+;o�h*�����V��/ug�����w�e���o��f��4&f�&c�a�\�z����x��$(�u��mT�(�y����v+�����.�O&��|�X�	c�㶻qک�6�ދUI�}�֩���~��[�0s��L��$�t��<���:~(s�geaA�E�N�����3�6/?��,�����]�㢖 ���`o�ŲfA���kf&Y�fI?���޿��i��������>8�Dfgg�g��ɢ5/�f���P���>��I��*{m��IVk��=��Ӌ��F��H�t������8���Ɗ��Wo��7���[=�r>2�p�.��E�z������פ����[(wg��YzA%!A�]�8Ve����Fw7BL�p;�e��ap��-����d^��.��Ϣ	������M�^�	��1B���~�/<�&�������R�P�4�4 p�D�b�1�s��*�8¨���¨�Sj�w""���K��Q��a�ynZ�i�����F=�O]5�߇w�p��E8�3{w?85��AL��ʖ����7�����a�.��}ao�r�8
��ĵ��ӌYG�����A��'�Dt��su7�^�7i�������Q��q���a�Y�]�����o0>��y��nX��wy4�h�n8�'���̼4�YQp��8JU*���K��jy��ϟ?��︭6�[u�l�X?
�.�&n���T�\F�������C������1#����)TI���W��N*MoR���wed	�b>���Լ(2(����2q���4�!3�V{;C�:�C�v����L�Yi6�OZ(��wD[BN�gm<���&#��e����5�yvs��=L4��FG����()b�%*��'D䨕�=�]͖	����ei����0)�xX��}.�<M�h�m�+)Ezΰ�LI������Z���-V͵��Q�3�8�A!JĨ�9��"�T�d`�Go��:����/��a�%�#Js�����C�;ˮa�ۉ)�&
�������OV����0�׵��}i��NŽ}֘�y��$*���w��c�ii��<wP�H�n�^��=ۣi�Ȭ
���4ٹ����ѷ�4[?S옕)�g�U	����Lj��s��g	�x� P�YS��N���9;�~�C;Vb��}�nHh4}o)$��
>>��h漶����]H���k�+��FA�?�T�:��om����=%�&���Fi��EEE{�Έ�`�t`�w8PM��z"��8��r
��c),T3�ҸP6�+?���ɢφ=W8��\U5Y��{�M�Ǣ2�*�p7O��a��<h�m��^(n����b��KJ�4<���v�h=�QJ�N��
��O�F#H�g�G峮)�^�"����$�;��S8���IFX�Rsr�:+y��=VVtZ�]Zzv3j<F���_���]Lsَ���� ��j�[��m����G�dȌ��������s,��f���Q��~�+�y�_�2
͊cG�)(e�$��u�Ʋ���ķ���B��Q�;����j۶�/�~;?"� |+� ���z���������'�YrX.�,ax����WR��i-����v�.I(KJ5*~�r��3�]�p���UaJ��.�u�f�A!���縜WFF�^iM0'�ć��}��s�_��v��;2��x�2��U�А�Bbb4V�ϡw	~���1���ջ�����C�� {��y��� �G}�#}�����������k�Y:/�ϔ T\FGF���B�@K�{�a��W��J̝dP����ժ��������$��5�����w�'��PWux�wC*%Nw�SM���h�����9M�>����A����ʦO�?G��^�%��Kj�hJ�ã��&p;���\{ �UZBv�c9q �%�AYMpo�ؑrND�i
��Z@	����Іa�8��ۏ��3~0{W�����ޞ���eF�=ߏ��)����5ɞ2�T~it$=���	��4������a���h#U,��*��{��/ez0���>�e�SE�dy[�9E����<���?w��:少���/������D 0%�+w�����p\�AGG�=it1'T���0(xxxTiv�h���M4GE�x�onm5��'�����˱~���f��):?��8���S�Ⱥx�0-�+��n��;�n��IDH��q�Ǭ�����崀��v;Y&s�D )dEr���vt�I���ֻ��{��'������c��, �t�hۗ��p�����:	d�s$��{ͥ����zz$�9Ġ��$jj"+�A[I�Y�n;r"�B/|&f0�aL�qOD:S����5^h���[�U	��v��=�E.ͭ�]h�o��p�h����%jN�o��R =M.:�sIܻ��t�8����U#)�%_�\�H��m���pʍ�-Z�ݡ�Υ5HM��Ӑ�t���	�#"��W]��d�gkBAE��N��e�/,v�1^��ü�_D�a���ߌ����M TB��H���xx>v>i���|Tow��|��aR:����t)��ƥ��H����k}<<<+�2944�GH��SM����Y@�b�Ｉ� �l�I;���i�-<�'T�k���<"�@�j8J���}A4�%  ������t��;��~�:%[/g? ��;v��]�y? vV�8I=�����q]/w˭:`"��7$�����F���|%%�J����F�63�?00�o�611�U�s�g�v	qq�����f�X���b!���Q�c��ҹ�a���|L���FG�c�=Y�%wZ�W��wQ�S� d^<��3�qp`�7���w�%ܿ��i+
xEī|�Ⴃ�������Ԡ��C॔J�['!!�_Sɷ�f�_���+��l��*.�����E06���p2���p}X=�q0]nv�)D������
��j����U�Ez��"|no�3k�̹+tj�����Dp�����v;�����E�������u[u{�����Gy��(����>a ��� ��{w����!��M�x�a�5����j��
~#V���fE>��T����Iؘ��7F9<����j�q�\@'�~n���`����R�ن�,>3s$ڈG�S�Kr��\{�J��;JJ����?�I�(va��2��ن�q�|�Ng�\��W�Z0�7�4��� �N素�����Єc?mg�i�������Nj�+� qxu���

+���V��}���{�Xݹ1�/�RFS��	�k|��R&�������W&���x�Ϧ������]nP몛-]�PtW��UT6G��(]
��}��b��t���# =�!��/�	^�����*Jkk>]�1�'gdDʧp��D�&��}u],�ևI)�����]���ugb"�m^^^��8M�����@b ސ7?����j�}�E�^Q�~�v���PLu�o�L�j�����,-�,�xj|�t����+=�0����X��$x���=�o�戻kL̽�A/h��H�l�{��G:��S		L7���`�ؽ���1����F���� ź~h�9v=��C'�qvD\l�����Vә�b��I�Jg�?h�6_ƛQ*����T��Qڡ�6P���=�/�߽L��ݝ7E��7pE�:v>)��|]�� �/Ǟbf��*��)QQQ�[r��cX���V�n��>Fs�,�?
�B䴜p&��#⤤�#i�Uoӝ<<BSR���B$U���?>_-�W)��u��~�N�433C�%\@j��jm��};�V��{q�Q���ڞ�z�@����M��.�h�6��
�h���XVP\�r�@A�Ì�l ������+6��i�Wq/	8�Vp5RL���j˥Ye�{{g�Fԏ2�rl��J9�n���GPȏg��,���vw�Yܧ�𽺀��وh���,��qM�J����E��X@AA'I�ڞGN��q�vG�/��O��FFxߛ������a�A�|n�f�t�si&C���2W2zoL`�<��Z�ĞB����]R��������C�ۏ�\ ]F2$���ED�H��.-���dw50�)�}C9�.qxQ}�|��E�Y� ���c��v��{<��?�bg�4�܃T�c����J��98T�9�fO�.6�lll8q^�zA�n���yv
�g�Qȿ�{eV'K���!fm���
;��R{�����5`��p=N+o�[�����h"�			J�������e�o�Ym����.Q�ʠ5�F���"�#'q�[�/��� ��Ǟ��c�>��*�J��Q�ZJ�R�Q�#��[��0iV����ىrz???N��_�L�oaX{��?Ž_�E����d�����(�����������ⶏ���_~~/`?����,KGO�h;[����������3l�1�������xC1��|Q�p��\��]��QaPKZQ�uK{x��d׍��+�>���7�B�]�N�Ji�V���߬�H��V�Z��م��LL�}��>���.���EDD�c��F�L�J��U�u �n��(k����ZZZ��ܔН1��s#q �LLLREً989��L�.�i[q��Y�^|F�"�Ѝ(�s��uB
n��ƾ��;��fd�Xq�B;�� 8���G��oA��O��M.���f%���z������'��>�����'m�p�����h��d�jLH�v��6�2��~�@�	�L���[�=�a���Ó�X�B�*@8��n������@�~/U��p9t���<�58Ik��p۟)�_�� #�~�����RVR eR�?<x�o�a��
	��w��o��Yj%�U]:��s{��	����XGω�g�.~�"����a�Jo���,�q�T�����5�{��x��^<�b��EDD���Z�������v(��`��8 .km};�E��+�R9I��x^�&�$
�c���Tkb��s IQ�;iij�����D�4�^ZZ4XR��L��0���W�a��"�娤��~{���� �z�b�t���Xc}##��u�.�g��הkgP��^��"��Oڎ)��8#E�����{܈I}�ݬ��h.^=>��E������b,@ɶ�E1L��[�K������Uu�x�ؼ^%#�c �B������q^�01�1A�@���­8��� ��#^�@C�7���E�RG�������4�Ǎ>t2a���x�p��_��B|�^��/�Ȍ��vq�.n��.��l�|AC���n뤁K6������Y#�Ju�/L	������BFmm���6|*�fH4�9x� ��t2��Hv�DO�ty�?�e��f�4���3��99kO��>W��Ty������`�!���^� x�2\y�Ls|%LDB_Gg�5�ڻ����nwl�\�M�T�5���A�!P�`)��|L��V�}5f�^Jq�p}Gg��J]���D�4-=�t��7'OO�kFz4�����TU�3˅Tzz�s���rrh4ק��R�##��f�Tqr?��~��R�"e0���\�23���l��i\k�#,T͎Ȋ@�{��l��a�xg�����i�)��-�[��m��S�����i>|aH��[y?�3W���;��xz������f�΅�[qQ5���x竑���,�K�8X�q�-+/ov������-M,���=f�X_���^�&�~��)�}ɋg
�XY�Վ��Mp����N�8|%#WD2���p��N��e�c�8}�#S�1铭��� 6��w]IX�/KF@@�iIz��bS�z��HLNIdT�eYmHא-n��I
�==��}��7�_�0��V�rU���'��^���CjZ����4sM{�������xR��h�47��mhW�o�bFH�xy{�~���2��g�1�%|����ES^��s} Hҳ�@R)��i�·�K�3����R����!��R0@��Ԕo:� �rejji&f�Y��ڂ��Y)G��Ԭ�����3�3m=�@�5���u��]&���Ƥ��/姕��r�,b�@!L���󽒜)�����	��@E���Qt���7O�qq�� r�D��ŷ� hA��5�voj7��\V����_- ���j%�?a���v��
]b.��8�����e����P��{V�����ݱ�'tx��c��(3�K_e�(��r�Vl{G����)����{��sE�)%EEK�2!�ߌ��3��=�4�o8�x����\m�B��k�Z�ќ������b�ˋ;T��D�:�����*e	F �������J[�����y�1������6�$���|����ؙ�^V��b����AB�տ��֞^}�s��"$�����c��j(��
0\ݓ�����2�K���`/�1��J�:1ɾ�P*����$j|g>���
?ۣ`ʌ���ڿG�@s-�K������ Ƙ��a��;w<<<'dA2�in)�D}Z�f�܉`{z��#�k;^WǢI/ G��C��c(CJ�ʶˀ*)����<nb���!�k�u|/8����<5r��Af7hc2�8���s4Q�_�~��g�7����}�R5z��=��uF��0|�7o��#�g+{<W!"��I���Pc܅����,-����5*��u�Q�I��'a֪(��҉s܋t�����و�������gI*��~Xnq?��W�A,��<]�f`@�/�(UC�\>����|����S�\I$�B�mG���:��@�~x��*�^�۽E�TwkSĕ�� ��� �lv��w�i_0������tl/6�� �RbFݼ�-A�0U�S�ަ�>}k˜��� ����S0�pL6�>�����oΖ������8��i:33��)X���n�{k{{��c8`����, �#~��.����
N�nyd��A^k��q������<�H�e6�0��O�4�Jp�g)5S22r�?�.��Ў��Mako������sD�g�Q��r7+:��q��d�$�L�<����p�'H:�>`�z�;h�F|j�Wrr��W٩�?�Α.��]__��u�Y�]@���,J�-X��F�e�5g�՗�K���Y{��,ZR�E�n$��^�8=��0�u|Nd|�@�����x�o��^�Z�(;�|�)V>|$+�����E��&淛Dҁ�ҎRv�~*��������Rs�cG�[����
|=O���x��IUut���{��@��s2��GG��<�{b��y���{�7�#^�/���rL.�|%�,���,��0?��̈+{���\Q�����c��Z+�	�#Ɏ/�x�����Ft�I�H�񍾚�Z.7��7��	������0�:���P5d�+t�f��!��3�Z��y�:�ߍ�d���r\���>^�h�V�HM�ny⻋��D�y-l�%��+[��0���>+�wi�i��B�-����,�S�=��uji�����Ly���11���7��]�HP(Zh�%�����q����v��-d���
��_j�r>�D���ds�K�]�5�>� )Liׁ��4Ow��>��D�©:Wi���V�}}$���K�uX	���+�K^���u���H4l�>��V-s��!|���J.���d��9�7�sB��$0�6�\g�=�ߞ��' ~��7�˘�<&�qЫ�#�`+�zR��V���2���s����=--�j���>�e}�r�x��vL�vt4r�^7nYKe����1:Nwƀ�~�
ͥJ�T��e�}*�"Wq��	v�	����f��M�Z� � �Հ97H�ň�0o��v�mmҼv�����0`��t8�˙�u� �-4��[ZZ��Ձ�<����VN���A�ú>̫�cbpꆿB%�%0��O�)i�p��j����㠽^��"M<g�Q�O6���#���RW�cǸi�	��os��/�E�x[�[�T?ܚ���ip#65kQ�cN�s�}Ī �z�YeP�&I?�\Z:h�mDHw��]Yɞ������|����E��	P?\��nAo6��J@��=���6�+v)dl,v^)�(T�Y/TNk��)k�6wi��L.|Ua�(i��{�� ���
�XWA��~ZU�C_���	�A�>��9a�k.P{����C���Sr�k���V����n� ��Ӯ��NK-o�-�Q[T!ƏI�R6�:�h/eQǥ>jk��Jk��_�P��n�{�^o=���ڊN@�P��x�L������\9�M6�ə�B������1� ]��o���).[1VV��{udd�EL�4�*^P�u՚�3D�N_���n�'�r��]��cvo�0�ݘ��:݈��ϧK����w�c��W)�0Y��d�N ���QRk�Ze�$��f�w�Q���A�ջ�_#�ٹܘǿB0��X�"�# �s�|�k�pX�1�J�'!1a�ę����̰]�Y�j䈔Ӊ��_��A���\B�D��z�禽��	/�$˗�-�d�����|VT��p䍕Ѣ���A pW�d���z
	e9k9�,(���O���v�|r������_Bǯ!�0O ��S;Db �b��$n�S@���w:�D"�ݳ ��w��� 1��b����"0���^_��@������>	�6{"5����pq��+ܢ1��9��{Xp1N"�0�h����#ʛ�?��^ ����������^�4z\ʇW���+8�Z��Z�O./6�tz?��K2峷�r�@���d�:�l�8ɋ���Չ�����Ș���������@n��Sx���?�zG!6�L����c�i3s�61��[-b
u��{z{�b�� �M,�̦����?:�1��9�<�hhl��6>���R����)�v���L�u�xw?��̊��{��&���C�S��]	c�E��6q�]]]�Pʹ_jj��\����5�/��~_�l���,���Z�lº����� Ǒ����	�e-�4����W[M�?J]��(�B)nŽ��Vܡ��K�Fqh�x�R�-H�P�hpA����~��{�u���u��5$�g��#3���M,/é�K�9�f��u/J�0��Rj�8�?1�K�֣����òӄ�Dn/�\Sn+����HɗD�k��-럹)��y�՟jbb�A���[w��<E�+&�%ց�Y-\:`�k�W�y�z�l����PqoG��sy�3��Mϩ�D?�p�&Oc��ϟW���*V���&�z#������S0oS�2rP[��[r�zz�dnbw����e�GB^�Ł�%pޛ���1��,��-buX-_|@��>`�ٸ_�9r��d�odll����	�a��������޾I9�g{�_SSٜy��P�Zi򺌼FDtUF�"�Z4�	d��}��$�'��4s��.G��˭�z+�=��hJnOVSSǧ�Lr_up#�S�ی�=�H������@�\l5�/�~�:���[�yU&Ӹ�v��h�R̠�@��#){pc�;�Hd*짴u~~~���թ3(ǠQ�4>�IN�n���<�cc$T��e��c��mL��v�����Dt2�LL��]�j�����D���39����#�Gs$�/��!+����N$l���#�H9��(Z�
w�>��+Д�$�v���b���O�Z��R�_���"K<��Y\0��"��[~��9وhm�*��6D�vGQ7��Q���ׁ:>6�Ҙ��u2v>���G��y^�w�}�c&,y�dn:co%]���]y�ZV������2��Q�DQ+>jq�,U��K���C���*|͂�E�F��:V{���#���$�s��q��҃i���*�.��
�v�0b9Kx�tۭp��Y\��kِfS5mi�@��Y� ����mm��$��@��ᩐ?���Jo������V\�Bcb+_ )�E��.�occC��x�9�:Tu/W4�X<Sљc��N[�Ԉ
pWۜϣ���!O�3����=e`���V�)Ӎt+��+ϸIlF�vښ��]���>]�ݿruޡ�V��9������@����M�504,W��3҇�Z�'��@ z������s�c �;-���!x���6(W��O �A�����Z�Ee�p�
I����= W+�l7S������C��ϖ���x��B9���;D��J��Ik�������%�������'j;����f&�vzA��B�>��f
ʔ[|'S��/�o�EMS ���r�[W?��Z����
ת<7F��uz��e"Rd�L!��PB�a�u��U�b�*�ze��3���!�R�۷rI�`O�d���(W���33k�Q���Z5K�6{v����N�&sO�]���(A�q�Y�ȅ��T�YY�G2k���?KKUP�C[y��>X�Gj*�XɃ$r��Q9���D$������b�*�r�/�"���<96y9��B�!YK��~�zo���c�[p�գa�_�􅼡��r�����,S�X�@�rzhbDJ=��!:��SZ�����"+�yd������YGO����f^�Tx�y�x�آ���� ��˼��u�~Y��\��gٰ� ��+)��o&%Ój+>��2.
���&n�H�D�7�������}} V�D�������ҡ�E%��M��V%��f*��?��i��_$ke�ǁ�VU��M�.�����������f-'c����3����7Q𚧧�͐V�������y���zȯ}�}ހ��`�}�\9U�}�n�׍��I���8�y�ˋ:x��[���b�X�� �8-7t"�S�������f�*�R��7�/��n������T-����p�r�̓W�R��i���s�s���pi�>D�&!>�۞T}鶄;nR��篘sג��NM�� Wv1�~�j���*0��������_�U�<���3'9���7~���� �
��-�J3��<���^z�OD>e}�E����@G�v�C<0Mm�X�����dW������� �?+�ؓ�#�11�����9�2�Ͳ��l�K��!�E�7�j���'��\R@�|���f�������w�q��Ɔ������X�'�~�� �t���l=X����EWO��J��Y�T�b����>�������\~��YQ���|�Y�ʩB@�%�7ޒ����i��ȶ�6P�|���:`�W�@�0��7:���
7]X�MK{�ZG�`�+F�0ƖZW��"�ȗ��ގJ��0Ǚ�����q� �DY��E���\Щ ^���;B�m}�����J?�SZ��^�mm]�/`���ޱ�O�1V�
�+#��r�<��ܜ�!���<>�.����}���9�:YHJKH9`���:QN���)�)((x�07��3�+__!�:kZ�os|%U,HPDT�F�J/�����������p���"�߷=+m�K�~غv[YX��D�S*��&��~;�{���F���2�-��ܟ���V\�\y�tX%������I9�w���P	�_$E����M�f����2��:�u���y���O+��L�nި�L��ӳ�7Q�����N����Sz++{U��Vf�P�����O��=3U�bbi��?[Z$�k�ɴ.ι��7���|�ż/�aS��i�N�a8����ln>��"�,f���|�I�H�2F��,���Ȕ������Qu��5�gcl����9���G\���'n# l���ǳEX�3200@�;mz�n#�l���_�����mjoww�,��=�6�bFp�|��΢�ԣ���*GǨ��3γ����F��'�B�f��踱��~***.ˍ'��_e�d�8)>�_h���"�j<ܝ�Th�0f���n�</�k7�@��~�yp4��;�a��w��n `���9��ΐ�4_��W��:�Hq�5ɢ��?�ו�y��Z9��e-��x�_q�جQHn�7&"�O5��m
�s���f�)z3�=Z�+��UW6��c?�U7���Z�#�(J1����Q���\]˜h�_g�=/�;�^�O�L��B+��o<K��z�I_UV����V�IF�מ��2o�����$,N_�S��t-Ȫ�?�#���W�O�f෍�2Ne�����!mmo�Mǃ��K�f�p�h�Χ�\*?����A_���(�M�g��!���)��av��y�'�އ�޼q����������ba�Xiru��������lȱO�)���Պ�����pB������t�t]�bcc]������,v/�P����?}��[>[-��;y�K���J����ޡC������q k��Ύ���8!to��`�	8
W>�A����K�ջ� yܼ�<�r&�X[�ZYYљ��E��S�?��v����m���8)���X@XW��m���1��#4br�r�n159I��H$��{���jo�Z�=a�Dtu�1VL)tI���$��L�.�I@�7�u�LL��۪�-S&��wֺ	�����-\I�S�(���P�lq�;������v<̣=/ݥO@bnER	����A�y��(#Ϡ����^�m	NnnI'�*g��r�_R��E9n*M�)t���ǔ��B� ��S�2�N�����v��y�]\\|$_]��+����ׯ��v�L�j�&���	��!9���섄+��6�����**�~�_�h����{�	Lx*.���z�W������SP�VVJ���ϸ`�'q�/�cJ�YjLW�N�NK�`����][��.�-7,ӣ�	��,��P�EC(�� vȩ�i����^:���{��UTT�k��&8����9�����ot3�Y�jǞ����\>��d���m�䏎i��Í�x��:�̞�>^
����`�߸cVv��T��Z�A������e(�< ��!�: |�ѝ������fa,��4m���/_
l��c;U6M˟,2D��P�:L�'�����{z`j@K;񈼑��q4.ވm�w{���WX���%�$��V��4n6��j�0QkBWY*IN�m4�����&|kBK��Փ`��+b��:�#�S���n+�����Blw���=|�5#ؼ�Hhoo?��x-��_�ϒk��	����].��H� ���;%F�nR��߽���ř�D���S�Ne-��]��>�eH\��eD�y��c߃���BG���	t�2y�W����V�eấ1H��t+'L|BB0�~5癐��x,W�~w�s�޽i]G����v��~�^8�pK���(�6Z�ٳG_Ě`�<z�������#����?4��珬���]r�g_��҃pһ�V@ُ��k$O����T$|@�zt��+���r��ܪ+pg�%H�&@���	�DBb�9�p��b
�|���ٖ��Lh5�OOM7��L��}t�NI#(y�3����.�����,�ۨ?{
��f�|ߔt��=|�=���hq�~��
��P�"$��ݾ���e�^!1h�0�/��# �-�V�SqKIUѹ*`��=6��'���m��>a�����Hn��A�I�+�r�}L�߸-�F����ㅡl��@N6�i���&ץh�L�m��g�=�G����&��wQ~��d3�~�8��rz���@����5��yhnV�0B�M�HH�l�K����6w�~.o��NuP���n�ȕ$�Yg�ً�����=����;gn��z&�2��^>��+��V���B����}�����֘���rj�u��D�����C�dW�yWEA(�(b$q��Ʃo�7$:�����łO�β?�.o5������6�}C耽�\\\,��^-~i~���K�L��4��25�헖YǞ/��m^1>�B�f
7��B|��xU��3���H�ͩ|H/���X�M���U��MS��ZҚ�p�ٓ	�D��P�X�>S���.��#����s�]�����VW�&mJ�Ǚ+�#���~�%���̂Ov���\m��xw(E%��j�n̞`�O:�q����Z�ș�k�w�}�v����K���@���ɳ ��k��~��J(��5�
��d�%*;�4�ڽ���G�/������e��yp�k:"k�j�%No���HP�Tn}�eZ�q�i���H`�!��4������|��B�	�^K��ݒfSQ�QOB�J��M6���w;JpsD�v/���H��B�}~��NcQJ�[��TV��{a�ܻ��.;�� �;����S�9X�D��T��A���L�~�a����=����X�IH�O�zYY��ߧ�|?Y[P���S浢�b�Mv|�[�3e��&��z�՛S��T��~��SSS�;G�mD,�|�� ���Y�w��jfgĘ����%Y܆^5Ӈ�J��޽u.�负({6�R+��Ғ��[��X����~�,"3B��}�fX��>��A�����o<U>r3
<�,p.L���4��v`�Z̔����*乑��~��졿r�k��꠮G�fq��!l)5�g�~|��MMz�냕 �[mp�6'2ECH�֖���_�! �(���������KK&ꩅ��rr]��b�!�%�%�TM��qeF��?�]�]�v��{^	��)�0 &���y��Ը	��;���D���]�SQ���|w�����B������2 k|���yu ����Hޱ�0teY�{���i��6=������K5|�h���({����c����M�k�M��]vcE;.qD�퉻�V�w��� ���~C����;x<��QMŒ��^͊��Oܑ���~s���R��Z��C�2�'�����{���}�p�����l���3p;���� ϛ&��q���]��y��\5�e�h�v����c1u�͇�᜵�:��n�5�L®(*�\��AQ��E@%v����n��k�!��"߄L�(�w�	����+m����/��b*o��y���e�}5ğ'eg��&���iY����zR��i����ך:]�{yD����E(@��~Sgw�wդ��5/�����ϝ�21m	Է�v�6��J�}��4�����������'��KXH�+���fVM��Sh*j>��1�c�GC���1��ɬ��#c���Z;r�������o x���IH��杓S�,ė��b�Z�X�خ����kx�ٸ��<۴��0�"����+�5g�@q��njiiY��qQz��3�X*�=�$ �z�.$�s�WHh�늻w�z"f*P��o\�(�_:��Pu1���|�c:�6�v�;%Ν��Jd�k�'�FC1s��<l[�������E�V�������g?��W�!�Uz��	�����L�[+*�4n�_���I���{|�ɛR�W��~�?M���;��#"}�� ctTq.SP�l�0�̭`|����;�֬������Ӄ�ś30���be��T^{�޾ ����Ɔ}3IuTX�ܳO|�GhTvj����Tէ�FQ@t�����f�2
R�^���6�to���к��'�iI��y3�3`��1��b��������Jj��&f�g+/���V�[�lo{�5��!)9'΀�WX4����]�Ӱ`%9�Y|����==�������u�r��~���?`�`�c�ЯM\x7J���M�z��Jւ�Z,�^!}4��r�_��f��'�N>-��R���o�o�/�9o$^Ly����nA�����y���{4z�|k�*�9�|U�O�����LY���V�~��/�R���ϟ��a�bK�b?7P��鳥{`��+'��R��gʸ#O����/���g�_X�5و#��1PO�7�֧�eF�-�O1jn��zx�=a�S�N(f8�9==�i/�cF2��z����o?�L�1lڏ�yu|r��2n��/&o�T)z�^��?r+�e0\Ͷ6V\�ܛ��D��
-Fq��c
S^27^-@j'�xzzZO��jU�:������X��{����Hv{eNN�2���X�v!9q}U���c�����V����ҬW�
���y	���\D]�hi���G媤1F�����4�aO7�5�'u�Xր��Bm�����==�!����5W�+���}�AH�/���		��΢X4�\D��&�v�0�nih�����vs�7˼�r�c�1��8���ѷw' (Ŵ�7 c�S�3e�Ƽ$vI�x�2MC;M<����(�"2��}wk9?B�P��sl�!��_��>�zP�<�ՠ���Ӛ�TU8���f��%��s��E����o����z]������l�
��*��&!�
�����K�I2C����P��LP��9�XXu(%�N�Rc���8��b�)�&T��6��܄	��-�cK�D��J�
}#��y��4��N���G~��E� ��� 	\�,�כֿ�2�޿�)�{�$rQUS^��%"-����ͣ4.O�����p�K�6�v��y�͔���M�?���*�G��1�!)$�2W%�e�+3��:wz�6���
�t1�w��9̭6���5),�n�;�+����,��-����c�愻NQ�{"��]�V��66䍈�A�(�i~��%y�����-���`�/e��-�|{�l;�ВҰ_�-S���H�{Wgoi}�59A���Ʈ�~)�I��q́+kwW�B+-YR���m��V^$�r}��H�=�*�!��du�ʇ��HPp�=X���u��vgQ ��$���xHM���U�7Ml��*����no�)�	d�t3���ı�y��]����pg�M)uG��̹wA+*J%��2�$.N�+l8���ֻw|�-p�3�dW��p�)[�f��|�n��DU�aܛt=���RRH�N|>�7�%L��-B��䪻�{˼g�92j�Μ0|�9��gi�p2^^�}F��e��k���������^B>}�	(�r�?��qB�`/�|��7T�]W��>;dSN��ja��`ׇڇ���3�+YZ���m�_�=�Mq������0o��M���F?c~�^2� K�����م�RIQ��<��!<Ec~k����+U�biiy�^��s �Ԩ�8޹U�<��1��=�Aq�_���^_�˾���|�{��
8\K1��1:�����dŃVV����j$�����Tf~����7*����㢒�p��Osa\��BW_���Q�rT���̵pK��q��V�������e|F�E�#?�����#ǔվ��̑�SS�K���2-b��|o��z�W�=b�>{�X���pf�&<Uج����ɧq�F���jV��������j7Q��jý�Fw:�K��:F
�KKP�_,6*�[����"_�]jb�#��1�l����"�$����(�"��hss�G�<��o��O�]���
��ٜh6e�DP�b��[O�V��Q([������˱�cV��7P�������u�7k��g�jy]?��^��ʒ;GI���_��\���J8m7�/,�o3d�lg���E�7Q!m�y#��*`��Ru>z(�ON����UU���Xw_�$�/Ymo�J�����4������Em"+e
[� N�$Uo8�I�7TPPh�ԯ�j�a�z�'a��D�_1��W3�+M�����N]	(0�� �Q'�8R���'M�0����� ��+;aA��G������Q8��kV��^a����ޘ��^J���TJd3���;b��6�"^�. DZ��f�~9	���O__�X��A@ZO;W��`�������S�|�\B���I!س���\���5�!(����\��pI�(K�t^�Gn�en��y�W�i��w�g�޾}_������i�"FGQQ���<�_jP�})���*@�%-_�{�M��D�a_k���u��$�X������C=b��MM�RꯅO�w���[�B���ٍ��:�<٢�E���;G������x�t��)�#ja�.��t��Z�>rz8*���b�#�������ĸ�b$nt҅��k_{�BMD���0AN�/7����̶W����E�p����{.��B�QF%��0xH�i3�b��}��S��~�������d�a�_O��|u���G������O0��΅�v�vC~��ګ�K�ڲ�Էk�j���o� 7:3���F��ќg���W�cF\��0p�N�q��`sZ\��3h��b9���q����4�Y%���6������C3zx�c�:��i���b5dn:�ӊz�/�bkǙ�G�u�G���f�bf��xT��K��w��K�)�)�F�j�b�F���VM���V`��a7��Y&�5�4T�>|}�0�뫇CܱI(ְN/˭T����έ.��$�-ؑ�
e�פ}�G������B�R��F���˄�l��7��� �2��Ӓ�Vy!�ZĢY?�򑑫%�*5�C{睖 |}�
}��/���//�o�]��L�ͷ^�w�ח��nD�U�d�#�>Ym!�i^U�r����%�����h�O�3���.V�p�i,�+l�꿞<h����Z�7�I��ԕ�(s��M_svNTUUMAѫ0�Ȯ3��D90�U*���"?����}�ew#w8g���c�vY��í�c����}��>~#�t�6�^���u>���9�(�Gۿ������=KC�]��0��O7�{��T��P�;�C�{nM�/���Xґn�����$� ����N6K��v�������`��u�R?�E:B _�:w4�P��%�>>������Tl7�W<�8�V�r�j�r��nVi�c�=��j���ؔ��[�$�Nd0�Yhǟ]�A�f�)��x�gӯ���`Q_K�,q����LN2���me�5˩Z	w��/�o}�?��B+���ð���~]�c¸��oh��8M77W���+�_���#/0��,{p;EI.�T��פ��Tٳ�`E� �&�2E_�0zPh�ޓYrh�G�~��%((�u����oO�tǢ�]K����ϩ��\�����EMMM�B�P�u��i��h�����B�F���uɡ�����m����Rj�p��ZǖnLf���������s��
�L(:���Xob?�p��p;�����v$�^��KMAA-�91�O(��G!���S�G��|0z���Zr"m�@2�~�5�#�R�__<���%hnE�K����D������x�$o-��((,,��tZ��p�T�+���/��Q}�+��t�oTq���}������j��x�@�H���Ov�w��`n��?B�fՍ��]ؔa�=A[�]/�|N96:��$l4���7�i��fbh�*-�'ϝ�(�W��;����{4vg��r���tJ�����;���š�̮����,6s��z�`U>Ö�g���4Vc�IS�f�㮖Q�F�B�@b�E��ZZ��Q!I��ǯ�dT�u4��G_#�0���;����7��p����r��K	S�. �fwV7kfǲBc�E:��1��O�Ạ�(�e���V�=������ʢ�e�(���k��mt߇ܸq#�襺�^����g�2g���`D�g}\\�f�L���~W�l�)�)���c����/x���P���>_�)��%��bhRnRt/��AD��vQ��Ɠ��琤��k?�m��4O����n�[U���T���Q�H\\�Lm��m��<$�i�/6G2�������;�u��S��^�����}��G�/k�m��=�
�^r��V��ID*`��H�0yv�2�Όc��bzF��7�\�9q�XnC���ɉQO#�O��
fc�^) �"�s;�B��3S3N3^�N�g�VF�����)Ge�-غ��dE�ۓF���h�[p ��Ǆ؋�p�,�{��p�qݺ��[)I���7D ����]M�����Ҧ�);XQ��k�@��� "�r�n���]Z�������V;��OE�[N�PCU�[����u���G#����M#�����c�E�t�F+�W9ͽCQ*�γ�atb!k%&�a��+t��"[!~�&�>��A-}��/��)>gI�;8����f'��Ѯ�}q���Q v��$���0��KDW��}t�b�wKWCS3�O�	��	F��f�au��*=��qG�};=���e�(�7�����P�����H#��߿�{���mG<K�(w���|�� ��zN�[���-ȉ�uܻ�[[ۆ-ez�����%���m>[���x���/*)�� G��Hw����[�AL5�lEaA�P"��>�U�T����B��6q�H��;p�����J���oW|ǒg=��ӗ�O'�"�{�	FtM�1��a����=��"(TC%�z��K���e��Pt�EsVCCc5��>Ĩ��B�h�.�&&�O�>UVV~J�J6��^�mTeO	sn�h|�D,i�W{�4?p!j�MP��,�wj�n��nl�5[��D����s7�>ߠ'��_:�fq�������I��+M(���Q|��_�O����i�*֯�xrY�W�8 ����������0� K�����*�$��Ǣ��Mj4�I�1����A�J�L@��J��g��k
�b?9;\o���>үq%,��>����]��ʵ�dd��rC��j+˵�H��)����[��c��s��t�<�[�؁��2r�|[��CUw�JvnnJ���E�r �1"��nu9��r�w��lj':�"DT�܁���V|���w��:d�2�{|�Zl���ߕt���B��_���5��!}���t�%�G֞�S٠W�饘��r��v��������]-���M��7�Kt=�tb��ʼk��0�Znt C�-Z&��q&+�����ћã�f2r��L�8OnXP$z�ih�6�u]�v���V����w]��kp��I3Z�~G�!�Y.Yتd��̡�P�e���9�����f�ܖ�[jw�j��)|�c@���t���[Ǎ`�T�b�z�k��?���q�bTS�^��J��qq�fЇ8$ ��{�?v�H�F����Vl SS7�C�x�$Zi���Bt��A��

�z�fe�*|耬�d8�%f��wg�
������ٞ�/C_�*������<A�2����{��pT �t���^lڞ���X1��11�l����k:�5�qr'+-��t��̰FrМi���[����w׵���`̳M��[��>AP�'k��s�$6��������M��9s��]G����7'���r+;���_���h@F��e�E��f<�=|�Σhh*'�����l���@��d�P3�Ѿ�k6hy�{��<�	�F�#�ڥtp`om 5�$%%����N?�=�Ӯ��-��4��yy����P6�ZZ��30_��/4����ǟ�j���l�.���k�e=���I>=aga�!V���d�˓*ș��ƈ��tq�����Z�x��a���1�>bfgW�=sWG-��ٲ��5K�.l��/X1��R賷l��T!'T�OCa��ʊ����C�zN�* 
�EcJ�W��S���/��#O��}F�E��.[@���=b #_|�9S��==��:�G�q�\�e�ۚ�\�/�!yw���L��H��_�%�#[ ���R��<��4�3�Xc����jbMlze������e�~�Z	rv�n�1��}odt$�x� �
A�$��p�:A�F������yW�3��3]��З����p���ĔX�q@L�L�L�˳��3�J�i�P��@���)��hj=7������{�+��4ħ��8�!����a���K��tw�o�[�w��������;�E�>�
��$0��Υ	<W]L'˭������E5I>�^_T?N�ݧ/!
������Y)1��?��~"����==�8M�P,�x�8m@�e^������х)o��Zb9)5(�6
��H��Z ��������,j�ӌ���PL���X�R
��d�i@~��(��Qvl�����g�5U~�ᧂ��@�H�UTz�i*�dg�\���lgI���^�<mm�/�vy�>�3.�9����ߡ}$��y�$3����+����[�}��'~Z�(p�ͧ�3{���K��j����� nzČ���[w�л
P�������ɂP�aw��v+!>Go��4���������L����D��5ow���+UU��Cau7��-d!����vN�Ñ;��Sp�p��>KuWW�ߋJ�8r��H���~}��Ӻ��˶@�8�Z��-�C@Pp��~�U���)�{�3���Ji"��7eԿ��҇'乭���)i� �}	i��ʘu[�g]0D&�x%���qqq	�:wnF���B_������⩨z�`�M�R�X�䚸ryg\'((p�k��^PP�p�ƿ���47+�'̠�8��2���̮��\��_��A��R�?め���4DYN��R^P'��{~:+��c�Cr��sՄ�ܛ��c�g`�u�پ䚟����á�"�� ����,|�>����˗�	S�W4�B�Z���/8|����ǫ�^a���o�+�r'�=����<L2`O(((�
D������/MLL䕔FA���el�-��t�JA�杏�?a�����B=P/ꨩ�Q �Q���Ų�xWśO@N,--��Mnzҿx��P��&p̊��#"�����X@�8��l*'�/n�MU^ڜ|��&"bp�Ν�����x-K������~�"��]������p;̜J�����X�5vI���F��������zz`T��JZ�����N�"��7�\v.�<s133˃G��y�-��ʺ�t���۷o��%�-^ך���R)Mn֛��ʽ��s#2�����/����/��{�"8�A���wt0�ǇfE� ��q�w@�`�/�O
+*��������a��X4�4�\�d��bXɹ�'fG�r�b�&��/�HROAm�tc�>\����c���co_d����5�fd�4���к�Y�d������fv�b�$$$9@N��RG���k��-{q����}�'�fbg?�󂓰����ï�,���RV�	`6���e^��13�*��P�?M -%L1������M7wVV���z[;;��6p�j�Y�AR�W����A������K?�7n����t)tv���!"#ˇ�1lДXC��U��g�������.$`LuD�uu-�OӰ��ϟC�}W�UUU3��-F����7��"��N'`�zxT@/zJ�����~UT��̈�|��u�^�.?��3�ŀ-�U2��Gg��<�w,ث����z1h�z9�y��F���e �.�E�*+k����V�C�{�����	2��߭x���_>�����>m��w� ��9�7Z?�u���F���k������Ù+�n��zg��m�?��������H7���B�]-��Z�"z�/4��wE��xk��DSI�|��$r�[49���u�.��Ȥ���fC�Z�i�*���0� O�^��<��z�n�Y���`xEPSo~'_�7L�4m��l�6w���lJRy�q\��%�e�A�R��~�o���/J�g�z��Du6e�%�PSco�n�ȕIQ����>�K�2>۲�e.���	gO��v�Ք���6
£�7�r���(�4}7m2�B�=#�!�ɸ�E�r!�?���ذ�-hvR���n���iZ��U�������Ԋjk���N��+/�B�tiI0���[<f��׿���WJ����FU�w�%cЭ�]�fl�g����n���9��z�Vx��7�%�geF��W-�`e���5�똯�!�3Kn��L�����E}��Q��Ǌ�4S��ū�������&E�k�ݿHv��G6o��i��a��u��
6���|����/�k���W�1�W�ή�!�p�h������q�\@לs����W�m*IS����hy'��8�K$~9L�>$���/x}�2��M��ɿc��@�dA���\M�a�!�*��gM^�x�������q�տ���Y�;�ߛ����L��t����㬤V�O4��#[�Ő���$��_o "u��$�#�-��3}-;w½��ѷ��w֜������yo�����uV^^�b���O\�weeՐ���"��.9>���$$4U�Xk����t�u�1�cʨ�����
3x���Vȑg��kkkjj���6'�8ڍ��`��D[h�'���������T׫�͞��֜v��?
KSը��[�t|D�cܩLE�u��]~q�&p��F��_�T+//wJefcs�b����KCO���ttTT|����E�E�&���(G��?����[�		�MM���,���k�x��0H �����xV*В���b�L��oT��#�y�������77t۬"���k�Ne�/�ʏ;�ux��޽�O7�#�*���SF1��}3ouu���^E���
L�x<�>�``����д��S`5]�ܪD��q+�=	�99Cf��!)��}ܪ"Н��,���U��-#ҝNWāXG:7~���D�G�"&&f2�!��c����S��%��!J0�}��ɁBy����ڭ�[XX��G�LO�~*�q.|��V�M�� hubOP�g�����bI��םT^?6.{*
���F��S�򟊣"�^{HEUL�����MB-{��8��gx�R��tL����߿�~H��z��P�S�b��t�2_�߁�t}7��d
d�ӛSu�b��GX`���@�lr�kv%Z	�敓�!| hNw�S���q%kh��dJ�տ�ל�v`|�Fk��$�z(>���u��Y�1��n(B�w����\��q��5؄���^~�xo�m0F�"A�J�`�e�]Op��a�z����{��F���(�}�s;VCU����ys� IVkN�}���ͳ|ֲ�}�a,������t띅�g�,:-�����k#r�	#)� 8vY�?_䈪q2�Z���%t:g�c``Xo	g	"5̋cѶ�V���6^�� &��R�f7�K|�]�;���~J�zϭ��Gi#�>)�����U�j�S�D��%XaO�)X�� ��I�u��	�L�<���Y��{�]����B4�!��M_��(���ʖ�����zZ�k��OV�cTDĈ�Y�V�rjԱ��^�#|��cc�5Bɷ���Ql���1)�Qa�0%��R�cn�i�3�n�(V�u��v<���U�|%HC�nڔ�3�nx��CH���f|` �@@�H�-vDf��[�������S���/ܞq��^Z�0>�}�䭮n���y��ﯬ��T�y*ד�Fx��������NZ���^GC�����ҏ������̜�u`7WK��Ʈ�=��{oJ�~)�����!~����]HH/��έF�0e�%s�i�M�gڱ�����ʂR�^����ݜ[�6�}3X(�E.�E���)q�yy~��¦�X���-�ݕW�Y"N���y-����˳��ͣ��U~�*E %�[zMS�='M�M�[��1"[(����RaZ֙/E��ZIKG��E����"?h[�\7P+��3�,=����N�x,�s������tx����ȱ5��]�%B6�/j�.��.��2��
�V���;�������X�)L����R��'��3��58��j�)NB~p̘��/�B�"����߮X
���m�hܫ�G��R��^� �r�H���ڏ0z�Np���r_�'+�#������u�GM��JF߿��}�Ņ�7���#4��ϲ\xHs����/?k{4�K�^���4��,:�T�]�/�����?�������o��6��f�����SW�@:��'��s�����S$�0]��{��M��H�R�P��ՂX�4�PU�&z^�� -��7�a_Cr��{�"pPzg�n)ߖ��kd1u���@�7����d��y�rX=i_w��7n[)�^����y(������J�XV���K�Q���:�e��$!�d��Ծ��o�%�j�2��5�K$k�,#&<66��R���yh���褣n��K`k[�8PSW�M��zQY�T����,��Ʀ#Y����0����re_nj�F�o�$�{c��
��#Go�
*j��}���/�쥴����ŗ�Ń��cy��������{��� LJBAEZ��D��[��[�P���e%�ZVE@�^j�e%��v�=���=������9�3�\�̜sW�=�k�մ[�)^����4�X=d����-�\���������"��^V�]��V���H��17p�90T=��IK)��"��*ƽKW�N�sRNs�.���r���딞<	�����A|�{����� ^�)F�b}�]6�j'�/�ʟۜ����\c��o��t��7;���.�cm�8\�SJ+��>B��Z��0�>��t
�At|�X;F�'T��?�*���Vݑ!mFݑ�"�,�>��y���*H��7eAp|��+�J�����*f����v$�}\�@iu�X�lU����jC��������`�"�I�D�;޿�tyR�<Z� ϗ��Run����������.�Xo���E���t�;\h=T\��b|%�qyɧ�����}X�o=��X��W�}3.�*�
 ��V��w��0c������]�e�{�9���}�<�I��.\X?�S-w�>�B���n�ƪF�b�7%��/*a�f���M;�U�6�A*q�"b���>]`~�tc���I�0Y�	����Ө&�󴝄�Z�R����v.������on���哪$����c�ܲ���9!.G�B�{�h:xQ���w-��jO��5n� �xT컘��e�=&�2��JإW�z5��h�%O�Ǐ�����ܑ����%�L~Z�0�tp��+R+ ��E�wJ4W�����/�W����f��wE�j�kV�PO��-x�����C�v����@գ��Æ�[���/
��w�v`ݓ��5p���_^j��<N�����=w��_����"�������U(�X��^|��1X+yS�u%��Q�>�0����ݻw{��Hd�bu��_�ÊWѸS*��b�ݧ���jۅM/����L�*a}fW��6Us *櫄Q���YO�n���|�B�XX��2]'*�ܱZ�Lr�:�Į����.P�vM��B1my�~H�l�~����irn`�S�UDF�^�x4]�������f�fЮ�ha�:w�\�������F	�ۅ8Xqq�����W4n��1~����O YF;���[�L-���*F<p�0o�%��&7�ۻ ���Z��5��2��A �ൌ������	����������hDv�)�7�$�m�-���4ظc�bk`c�ڄLc�� Y�_C+ۺݿւs:����i�r�|�<U]2;7{���v�-#�j�*��jXgg��4Qa��:�&ő^X�c�,RL���q~g�Έ�,�S���u�8E �uuc��}f�ћ�P�fɳ��^�RR�d	�����u�cNM�&���k#�������(���d����v�T����n�묩6g1[`C���p-�;��{���U�h�§�[+H�){؀m]Vsh����c�O{�VY-{WbF]/�h�Э)W�$HW�6�S�`�7@�R�[��aecc#�ةf|�]A#��}r�����9�� ��h\S�by�Se�E�G7y:a%EZf�#�
�I1Skckejډ�'뛈��L�1����n��ڎ,��i� �'x�Y�'"G��~P�>�ဈ��Y�z��O�����2���+�$�uY<�3��#Ѝb[����/%�c_��M^�|wS�>��q��2õ�"����C�@b=��8���/=�O�|���|h"Z<pc�7���I�<��{>J��=R���sG��� ��d�
�DI�^�O�ub��8��g7�j�=����׋Y�I �/\��jny���o��{��E���i�a��VvV��e�?�rh�_Jf{W��(Ֆo:�����sܼ�x)-�)D�X�e���Zր�����ى���p�"��"��.s���U����G {�%:���������T�׷�]_H0ʯs],�����}�:���R���.���x�����s=���wn{�|����=�����(,��Z/P1�C��(�C]�B%}��ԉ���'
C41`��%��x
߭ly�*|>Iq���D���WN��2OY�gN�tϒܕ�/_r5aA>�##Ï%Y" y\u�p~,i1���F�����렊��\�&^&�bH�k�B�+�߯���xAw�c��k-��Ө���ps{�ٹ9����(�@��7�Nfdm�&�;چ�D���>��~�(�R���5�V�l�~���w�wl�4g�V�����\i���Y
��	<G�|0k]q���gfp�ɖc�]�ç��W�Q��w�|Z�<�o:z>��}�������>��oX�.iz>i���T�������B����>��􌜩�t�G�R��xU����@��2�g֚������Z�q�.Pse��;��	��g���l�\���Sa�Z�:�Q)aލ9i>��� ����(�����1�,����ѩ7+R^plZ��|#�j�<''��ch�|+�U;�sy�m>4dw����q���ȟZ��'�qW��6�j��P���]C����$&��==Z:I����dF�Ic�GT#�B�*u�.�.Ph��&GK���tw�U�8�!m�Qđ,�ͷ���@Lދ��H�Ў���5�V��a���-�~ncccN�N�K�p��u�;�55�N��A˵%L٢��B;��smXt3��+ζT}�,!�R]w#`<}��o�s@�l�],�w�'LjZ�iKF:~~��:���v�Ip��O:J=fτ[?��J�����ҹ�㿪�-�ʺ̴2H���ub��$������'��rNR��N��l\�X�L�����o��B,�Z$o�~*FU}����h�@�F�65�æ3C�(J��=4 I����+M ��yn�%?|��h�QIi�``����Ǐ�Do�:h�ok{�Û��7�������;���>̖Zj�QsYG�t@5�{D�X��}U�@b5�=t�߳ M{&��x\�-�A�H��&�(;�94��Ĭ���dUUU���������?�8Fd���R�[�6�EvA�}H��H]:MY���y���eX�/L9�&�$_ܡ��[�:�dA�l)��VV��P1j7�p�8��UTV�0g߲�m�ĸl�2>tʬg�z
�tqa!԰��Y����{BA�t��#��T�$H
���Р;2�*ك1|Ĺ���#��%Ƣ��%)(��CL���Q�ШS�R�4�}��T�g�i`��Y��ǭyr����9h��;1kW۬�?(l�+�d��*J+:�]XX�F��������@��d���R
�'h�;��z/� �h��n��N��1����]&��ZWqp��.�N�Dฑ�`���χX���Y��GAaA�m���W�]�r�& 3b�ԟ56�pZ׹����6U��г���K�#wv�$R�~c�����gg�X�7�w��X$�4rʤ���x`��*�,����Ezj��xɆi
�����7��Ao��/mak&&&;���pIHL��E1=2�R��'�z�/#>>��Gt��M�ju5�cb�@Q79$Z�GLL�7a��a�#\�LF��N���������Iϩ��L7�hڗ��y"Q����rC?.i]p^N_c3��!O�Q��R�'N��uzm3`��9e�⁺�ĵ�q������K�}�H_���j�N�LC#.��W�٭G>Wv?��]��81k�(l�w/��ȹ���=���x�zo�z�E���X�Ҹ��l�+�#��䙙s�����?+Mklxt���:��y\v���Ѷ��2�ƛ�%/���*xԸ��%���*�ق��C+�����@w�����Ý�P*}a~���V!r1�J.N)K����6�v,�dhd$���"��W��Z5�u%a�g"�eZ���ˇ�\�$��������/Q�y�fܖ�׌ �.���ўg˿��� �[T �Y���ٳ{�8y������'j�H�Jˮ�_%r\RR�*�%e�ϡ��ql��
SY9��T������D�4���F+Ջlⅲm�bY�gC;�F��V�W/]�ߨW{w�f���m�o�&0�65rqś^1�g���O�N������#�&C� �b΢�� ��[�S���p��u��^�{46U�	���z�~���Z��p�҃��4��V���j;;��{����BB��03?����Ǘ#�7����K�mk��(K�?!���sM�!�N�0�����e-��Ζ)ф�3X�y/���$�4G�'�,{X����V�||J4�[_�=qZ�	y�{�� >A������׵��ߧ��tH�lj��S�-�6�V��U�F�&���'�"�z�5�S��&�]���'��	2��p��:G��u���b�;����n�����M푆��"�]�h��u��GVh�����Ǐnã�{Ҿ�뙰�I���NmT�xGG>C��v3���q�9p���2���V����1$e0�:���"%�՘i���hӧH΍�����N��{�:����<R�&����@}�a�4��[/gAj�ޞ�������q�V8�V�*�5�����ʄ	�0����h�ѭ��6��q��(�o��7�I�DݑW��]�,�B��N�]�����*v�ƭ��-�o�\����sj�@�3[�a�T���3�e���[ZZh�\{W
2���$��E�:�6�&��\\]#/P8�ꢐJ4��0r�fΏ��u��=�Æ.>�v�������e��q�$�KTt��/'�>�>y򤰙B�1�#��l����������Ӫ�h? ��S.��	s�W��I���^����*��4�������WH���[����yF���C����nP|�ߚ�Y^`t����f�I���,��T(�v��lW<c%���:�����@�g����qB��z��cm�9�
��(��{�0~N�vR�w>���zm�� �q�-D4����ڃ�b�t �Sܺ]�SyeRU��'�rU�l;�_R���6_+{��q� f�a��o�0�^_�2���%x]��X*v��@�J�d�{<q}�(���hg����oMO*qnp}�,�,��%e;�^�'c>�x�K/��Ȅ,uW�V����p<��SZ�mZ3�����E�uo�����c����ߝ�6
��e��u��E��3�c�W��e�O��z��Yz���[�N4�l�G1��J�V19�B�O���a{�SF��]�i&}����쇜����c�׶����w׷�p"���9+Z������ ���WgrB�'��c�Ͳb�ˡ�@{?���ĩ�֘����c��)�4Z�0��s��5�L�x��wo+��mt!�����8����sW���T���^���H/�8�23�[��hWC 9 jƷ��2X.�!�H�,� ;�E�6d�� A=��؊�Q����b7e$�Ř��F�H&S�-��
²c�H�c+}]��j*YC$䝘*��fo� jA�yu����e��Mw��i�K�;��t]�t�]�<t/r]�rW^�s����0V�.�h�˻>�`��A��EFI�|A��4����'Zl֛a�.�d�T��J�Id��I�:-����u_]{����Q���J6���1,am��;@���]�mP�4^��0��g���b���k����k�+�>�AK�|��5�^vf�����������_䞩2
{��n��p���M���5r�w�8i�aR�kH�6�+-{9�w��l���~�f[v6�#ïb� ��r��7�Vm#�E�쓈�%��5c��Q-���-z��~'~�������J��P�>!ꪡ�~��ϗ`�P�؝v}��Lq��xS�/n5CՄ�(-tY�gT\��ަ�"o��g��\���~h�2e�����
g�h�Nw/e���C>���6���by�d@z�e�P`G���N�n�V���Y.Ȕ�IS�>L�>�*;��>,@����wBǼ ��q��+b+�ؘ(�ʸ@&B�`�ϟ?W74,��re������������^U� 3u��$�䫂������������
�W�Z��������@��Bzz��Mu>(A=3N��8�!3#���O+7�V�q����~����ԩ��q!�U���ٍ;�bi�d�_3��u��G��`��ůs��C\�s\5*�� �|�$�0(�xP�iyz��I���/�N{I���y�,����#����ֽ���x�P<TZy�;��u���߻��Rs��SAPW+�s7U+Fϼ�P+.�q	�K_�����ɫ�rk3���������=��<3��\k�@�[ݣ�����3�?����"�5TU�������Sg*���h�\rkkB�;v<r���dW�~�%����-�b?�ز�EM��P(^HX��O���6��WZZ	�΂�! ��ӑI&�D�6%�/_r���:f����>ZR�j�!:V��;�$ǝ�|��,Sy�X�@՜�ӧ�ߡ�&�Qe�b؅��24�;�̑�A��$Ҕ�YS�� ���b斖���@�w~�Um= 'z�~�LsX�����)bab��g�G&���W��V�o���8�6�O0����~�д?�W<��);�}x�@����B*�8���|�44�_��Y�yu(��hYӢM�;4�%�Ѩ�����%���rr���M]�$6.��ZF�ݒ�����M4���b�����
�qP����M6�?�<֬PR�PzU�ĭ����+�=ǫ�$m=��MO,��Ľ�I�5^��IW��=�G�>}� U�T���CW�Ej�⤤w���we�!BG��)��0��f[r���2W�+����������a�%e\�,�Z?1|��
�3,��G�/�y���B�(b����8�#��I3PBx��]Z�8�Á k�	{b(�D�/e��*��E3g0ee��a,�	�:����qȂ����bPKj̇��4�Nu��r�K���p������m�f4pi��ߒ�_-d���O�ϼt�*ԹtN�0����A�N��7��y�l���y��a�3��b����Yɢ^*\�L��]]Jgk6+����ǩ�C�{��;ѭRD��X��{fC���.����n4����EF]L�
4b�����~1��A�G�����&/�]�Z2%� �~�\~jP�$^��ߢTlD���:=Li/B\��Wc}e����|�H������:�<���(�F�ՅE8���^r������t|.�T�Tem�ׯ����!�|gg�ۉ�o��+d���T9`u����1]�o n�Ǳ�ո�t����\���?[Z���Pu����Tn^��J5ow>� ���k����{�QD��'�,�I���C��2̯���`�b�(FI���p�L�K/���SN�;S|��Pm�4�)^q��/HD��߂&�~{V��'�B���NS�	'.����@gۚ��=6����/_Vݫ����f��!�b������Is��gmf�(��C*�YR`�����rQc��i��&���Ҋ�z�Zy�2a��B=�Cu�c�z7 ƛ{�{��Q_��N)W�fQ��X�SWW�4����+����Ա5��la�K��NeXu����3�x�t�@�y�Z!|����F�?�����)!q�>#l4*]�e�=�,�Ze������P~iR��*'�f��x��)����\��ЩW�.�Pv������ֈf��F��f�Ռϙ��!��n&4Ϩ����h}-gggw��艥�,�6Vu;�T^�������{9��r>Չ�C��s,Wt��,����G��n���'����Аm����'�e��c� �@v�����j�|!Nr%7�*++|v�e	��F�+UB��o�Tۃ��ea���U���K�N�zzk����)�g[pqs9�>�`���������xb��'j���>	 �z���"w$�oc�J�,X� m;�!��5_i�щћ3� *;'��W�i�ʵ�X&1>�̓���r� slq����� g;�`!T3t��gg9��[��)mC�g�L:�D>0��T`�.�Ǒe�����3�,ϒӤ �=}B�~���KMY݆ns�-M�F�[ ee�O�hjZꛅ��ʛ49�ϭ�R�VxWB���wJ�^��ZZ����=�:����뇚�b-��2����g�;Y�=���j7�'7*�ggg�`K�+����ᇴ�	��q���u��_,�D���<ë��$?���*'O�_�v��(���+�u��]s��W���9)��/��3�����+3�a�k'�����<����oJ�
y�4��W|�U'5%X�s�+_1en$�qPd��d3Tl�{��A�PW7�0��������cWr������;Al�;=�֭&Q�8�¼��w�G>C�A������Y�,��U�em^9���D_���l��_:���T���טcѕ\�{G��� ���}M�נ�Y]���J��.!nQ��v�i�_�$Хޮ���mR�R��~	Ȁbk��A���0%]βGX�4�#�j�����iq������'%��^g����/p9�
�zL��hi�j���\C�:�sm�K[�;o���罜*�+qJ��R�5a
>��/y����W~�ut�m�g_�zu�� 0�W�"/_6�k�(m-t@I��b��6����QoC�+޲o�.fj3뎹���FE4ڢ��9���5���-ù��e^��*��5a�*�����'�m���	�vF^���Q�$w�^ڰ|��?��#�%}�������p���[��{C�kCA�e�Pc�hMĔs؝ ��7[�e�VM��z�5A����9��O�۠w�S�i��OUU��G���u�:d�Si����Y�9r��W�^M�E0H.u����$e�@r(�+(3�_�8Z
���ǯ,�
:+-�>[;���G}�5G$)氾j��d��a��*��p =+s��uu����S1<xG�ꎤ��6dd�qM����g���Wi��8�<����5mX?t����c}�H���B|�߂z������TvSY��4���èb^NN��L'~kkk�%,?8 �~������6o�S�N�|�%���9�L~�b*W���?���bs�P\%��W}5}��b��A��b�Pc��/���ϵ`5�`Ǫ5����GkjK������0����[�
S�I��,�pHLB��N̗��2�}���w��"�MS�f�b��Eĩ)n�215mޚ:�%%�[��X-�М�Ä�Z�W���uJ�ǹ�y@�/��'�jo\�š�M ��Q$�j���e�����7N>+{�؟��u�顎�}�	\�GYi�,�D���z?U�ÝI����o�O�!�;3gX�o���W�X�;qzOb	Ҩ�4ҥh��xtGiϦ��m��C x/��{�,�J��?v�!]x�\�y����)QU+贩N���e���`�����,�荋wΦa��"�1��ܺ~W*Eڱ��������?Ohy����m�xo/�,�Z�;M%�1����V�P�m�c[����4[��d���vݮd�)��)N͘*�߯��O���Q�smk�K"���z��H���$��ƺQ�lW�Q�J���))>7�����42�s�(������ޠ�AG7bmnTI���{BC) �)_1���]2���%:K6,(��Q�hݵڮ�9����'P�j�����k�5]�Y�l��� �Ve���p���$�f��������~�I��!���!�k_�!g���ye��k�_���t������<q�66\ƒ�-�%��Q$v\6Q�9��~ۖd��fˍ��������빯�1K�i�y�&��h��׻�0
��&�����.�ހѭ�%Ts��W����U�����~�m.���Xf�[x\ ����pwhge`(K�L�܍�w��ۧ����klb�����
/}�`��q��U�)�����O5���.Jb����Ue*��(Ƭ9d;�����8��	�В7�v�u��>��n�����T֥�w�)��mNu+��&�e�X�[Rܯ�����+4��T��:��szx�ڵ����O#�@*�,����a�v�N ׻��x�Θ^�^�[$V3����dtj#���=\*��Xڴpz����ӑGj/�CTG����ٻ34å:������Y$
��je@� "�+��nҕs�ʸ��:��I���|�s/�PM;���H��z*��l��y�]������c�֭����͖ұ��k,!p���E����.Wk�ז
b�஬��<*��f�h+�A��ѵuC�a�b��BV��
�UUUWG;A	�ۋ��/iß�����s)�p��Ez�ȸ�]��@3'C)+�Fη�ՂSL|���5�����i�cu�N�ᾣ�����R��t�X��ZQ��o����+ �[P|�D�H]x�����Ze;�~�B����)W.vչZf���[�P�f~�j�Ѫ�Ck0�� ��YX2;;��軳�
3�.(������G�o���˘>4�C6��e�m��� t�۱�>�����=7�� ���ID(�x���sa�&�z
��F97%�"bbb�������zWu�a�Q-���ﶌ�2qrV�i��k�����vp!�W_fW�/ħ��_%{�L-,.ڸ��^��7"��C�kڎ
�B��u�~����x����9HDk��+s����t�E����8ڿgD,�(}utt��������Փg-��&tJ1�����{��N����/��6:V��6F�Z�53���i�JmE��/_���	@E}�
�.g^�K���V0R:���]W��1tk{+.)��Ǐ�7�j�6�G���;�:���F�Kz�I+� �B�]"U�,<|�d�HhecG8`wq��6���RX,�G(�pޣ�n"�C��%Z�O��R���r�I茼t��U�Tϡ�i8��	�����B6s]-k5&]�#�SB��]�r�m1��������y��~ɦ��;r���m�w
��VTV|i4~7z��T�M���/��8�a<�Y袂CӾE�X���>�J˰��H�.uUV32T�{6ArR�y� 7��m=��N+	�r�i���E2w�Zp��|�J㍉:l5lǙ�7G#�7�.��s����R*�o@x�a@�+$3��oq�`�A����n��W&	�J ��t
�ܽs�Γ������s��uFK��Z���g!�e?�Xצ�2�[��{J�q�_��g��ԅ��T���ܐ�h��hip�XWDd��W���}6ȅ���1�8䖏�胋P�@��gZi���4�%ߣQZESw�k�����,X�!S|�#5z�ޛ"�=R����r�F�|���-,��N��ӡ~�N����H��??���US�����k�����h|�[�x������B��g\[U�}��������1��چi�l4-9`<��R�F�¿�)�!���F���}.�rv&*��⟰��;N��������쾊�#��+�>�S�d^�ɏ�MI?�p����0����N��Z*ҭ}v���Ҙ�Ib��� ">^i��V�?��@3O0�R=��6��Y�L�ɣ��� �{tW�|���1z��p���G�97���T��
F�}ݫ��v����mr
�;��_�/A�IXFTT4��_F� /z��)���|=����񧾀���T
��1�\��X��(�\���<��K��Co��Oui�>[
̒.�2���=���K0���N�|-s2��_i��]Հk���p�?4SA�A��j��x�����z�wb ����D��6��|+����=?�����J�\�F�=��%qE�~��Nk��|<"�Pw�g�<	Cj�?FF�Zo�H�X�J�|w���$Y�������<�\4�~�ڀ�ٛ	3�$R�Ac��E�#������x-=�p�2uK�vP��D����&�B�&I��tTn�-�u��`���2���a�

�E�Ƙ��`�*k`�N���ʑ����=29p�<a_���� ��w��t,mۢ�`�9�%�	��3�l_RS�<>=/��|%��8z�"�$��ߋ5���,G�����g�S�D�L�_#`#��v�w9�G�]����P�u�e�T��*�/{��jr��Y��'+�n�"z�����
7�4�5��Qx��8���|�"��V}�*���`��#M��{42�M�!j0D.��g�����?N���ԃ�~�G��GP�r�����>1����D{4�'�{n�O�^��w�R�>���r��AG��l���^m�5�O�%�[p��z�Wﰘ�=x�b}<CoCH�AT׺��i�����w��9��a���k�{.��m~�tW�e�uvL���?��We����_�L�u|o>�`h�mm�[<���v�%I㆓#��!2**�'�2���{��e֡H��e�.>\]��V^y��=hK7�w�`�6�}��5%���L�̨gr,�ZY�1��=kq����)�5B��E<J'�y���ږ�E&�b=즲 ���P|�@Oy5+`�/L�C�.�>�3t�^po�T���*d�`׶�TCC3��M���!mF?& �I����Pb�, �k�N�p��-����7��	����o`����� b��&1��:Ԇ����h���qO����_aJRf�_��G/�PRJ_��b�ԭuz*J-w�S���e�ip�ƚW/ugA{'��K��'�<�?�3S��/�j��Z�|�1Q�4��V*��� ����A/'�
i��j���vm��FIl=!��r�7rE+,���(�����A@�M柍b�����T��NcK������y����� `A*ʨƭ��ߋ,��s�@�ُ��Q\��zX�K?I���{6�f�t���{����SL��>�M^�}�T}>�{�((�57�
����uXh��m�w_"f��^����B��6QÎ��������J��U��>�H�O���b�_Z,z�7	�%��啕�U���\����a*4�HN�E777}�~s�U��SQD��_/#T�*(]QYY������օ��qh��Qe���Yw��.|��7�#/e�։�M�C�{F������ �p�d���E�[������:�_���PL����
J�][�?��"�n�¥/�4���m��rw0P{��3{u�~�G<(a3_<�}A��U��HN9�hE$�<QL�R��$%� b�`ѕ�g�"a_� ض~aXO�%���$~ݳ�ّ���D����س��8��`�qo]TLٙ��|��܋M��ń��D���X@>2WVV���z
R��mo��j�����f�ٴٓ�x�[V��V,���>Y����dZѮɪ���YGw�ir;*{�`X�>ǜX��׌��g�+��rq=G��=�nX��,��9�t-f��|Ui�uĥ�0�z"z�)�t�o�L�L^��F[�/�A�R��F��{o�h�[��cx�k�Y�%���**K����ju�mG����G�}�CZ��ۋo��a>a2C�L��63��;/��`儮b+PJ댜��
x��D����z�%V��j�ݡ2bhh�V�.BS>A�Q1x^�qxF1T�g�zA�A�Az�#m���6O���rE��`�]�<tI��K��=V�֑�4�;A��@����GVC���Z��y=sZ<FYȢ��/��fD��C`4w_�޾}[c���j=ԾrQ���|��l��6�(t�)1���w �w�HZ�e�P��)�8�H� �9�}JA�������K�j ��Ǯ�Z,�H�����X�&g������8����l�&�-O�`��P$�<#���Y��QQ��'������n񀮺���������x���������5����zDX%P�	�3�׺Ώ���\q�����,jj�h��:������kNR	�ͷ�4q�34,��rq�@��\���'�(2�$6��ம΍*]���Qo��U�Nh/��8�J�>u�,v���e1�d��s��r����>����^���w�"X��A�*I*�l�r�Q��C+����c��r��g�^����k�PL3(�~��6�4&��͍bw��o�
���*��D<�B�Ϳ�h�ݤ3?�������ܱ�Ŭ�Жz�5��1���S�����L���R�z7o��V¯pdX�b���e�&��Z*�\��ٷݬ!���n�ݟtt�1�4kY�ь<򠝛��]J+R^�A1�Q�����_�H��Y���R7HUqB�$?�Փ�O�g�Sg�F�J����3�����)�L�bY�΋fi��F�|A�������6�ϸ]�V��ʤԈb�j_*��8f�N�/⺸&_BG�&� �3e�Ŕ©kD?P��I�x���<%�eꚚ�u��.Ȟ��|��!f]J�����#��3����5�u�����/����Ӆ�ۧ�o��3qÎ+�G�b�T����𜋫���a�d��m���'�4.I^�#� +^��j����[��L�!ʠz���pF+y���^�����W��-����a���>��?(�18%�Og裪�"�� JUhC�V{��n[����&���v�\��cn��#��UΝ����cyg��t��[0?�j�-7mk7�X��0?_�_5���*��d������T���_k4T����6�6D���2�GM�*Gx��ǧX���W}}?mI~�Ь�	����BEqxT����'�Pӵ<����T��ٹ�kz�d�%(ر���e*~x54�B��X�kBϜ,/ƥ����Y��C/�Nwe���Om��_�)=h����n����������@��H�,վ4h�Y���M_Ǳ-R��5<??��>���S3���,�1�C��ܼ��5����}%�2� ���~K`�eO��������C��'����7d�p�M�M�㧩^-�]����H}8x����~��_�xttt@)��OIL̬'�l{a�� ;���Y���ocT������H�-��9����ffh��k��`PM�T�c�8��C�K{�"��Ze����t��*��ޛ����bb��a�0hz�Ҳ��3��T���s�5�n���5�B���R��Q��GǖLXcd�؍f	) �_()oεA�2'��L_�?ۿ=PhP��w�1R+E��������o��i4z9����q� /L�)�h�<Ͻ�L�0XX8��XZ�:X�#2�'j%�3���{&3���liY�
HX�i+QJ�h뛨�>������
��q����Y����%=�&��d�����E�g4��M���:�sO9�p� �������H��.�57C�b������ u�8-gɳ�wY��"k�TIKJ�*�,/>�Y��_2T,��^>d�y���P����=�n�����$"ު��T�t4+m���aA�G��)ɑuz�&��s[DiR�ss�9�j�����Ȯ�OH}�ׄ�Bmp�j9�����SY������B��7��w*٧Q�O~a� W��j��f {!�֫�|Opy���*�����F����l���f�^iz2�c��uެ�4�L7i!�^:W8V]B`�e��g�����xy�JM��իV+�y]� y������P���>T����~?^��B� 8�Y+�Zk ,�"��0��G`�G�a���7@P�{;�H��T�Uzj{��}ŖÃ�¦Wg�rF! n�:@8�;�+Ҹ^.��_�q�-a��Cvڨ��� ���n��l�q�+E���>�n�qD:���nr�M;�Z��B�?�tp���r����� uf)/�z^�ؿ���w��׻�3�YJ���-��=>q5;x~�%�����E\�D�����5�Seu�d�?~Qm؁����2�>~| .���8��h�</����~����n^'�	��B9���ǻ�(i��j�����ȧ�����:V�|ɥޏE/�.������Κ�^BO����Uh�d��r�/���: ���1ٓ%� ��tu׉�����S���j�ό�tz,���:�Fk4�|�*3��9��j��ϯB&�Ӓ��/%����u����.mDj�ДH�������y���/l!�]#��,�V��X��X��3g�7�H_[�շ�T:��`�a���t>�St�z}P�q�4��s��\7���a+Ia+�m�Z�rlz<m�ԅ8X!�~Sz)�T�����7�t�n�{��?��9>�NT{J��W߹��J�nb���.�؄���P��k�A��v�鐙	�6�4i��p���U�:{������Z%��6�6z�mx�9��qJ���j���g�C[s�E��H9��e�*'�$:Mo	�o���{�ѯv�2�k�ðk����^��+ዸ+�;��Y�Ǻ��+��Ȥ����8����5�@�J~ˈd�v�8���/�P�����(�\y��੷��cnii��O����{f2K�����,���bn�kĝ�.�Nh#~�[.�ke�����P�s�e�� �+�`��嫪�J�_�=�����O��}���:Ѻ|������Hf�#C�Wa�_H~B�cn@t��	�I�(�[0]s]��{;�M�%�F��)Y�d��k:j��*�5�F$���*P$X?�w.��.I��.�|#��ť3�j��Y#����р�ٍ����/��+�?t����|Ŵ����3�������|ԝ67�������
2-ny���`���u���W�/��r_����NBAA���hs�����;�1���=#�S��[��d)�|d"3���=�VnI^���K�����=w�g_�	趈�,��@�"��m���v�,W�g����PU�0�4r�x��J�c}�x����䚵�x��?�կP��\`bb�T��o�%)^�I������3���`��a��x�k�\$�N�CB�|�_G����U�YGL'N��ŋ�ѥt�U�j\/��ṭ�;+wEEG�~��(ƴ��2⍟e�Ũӆ���[���8?}1:���+ ����!<��NQo�g���Y�S|���+�,a�+��J.��{��j���5�ī`�����˗�M��E�6���^ĚaD����~cEe%t���
���v8�M˄�<�0Ub�Yl�J_��s`UV��h�-
��z��q,�ؘz�b�p��PcH[DLl�_YE��>kLB�����Ǒ�X�Z�]]q�M���JJ�E����N�3kG������^����#���ں��F�ѓ � z%щ^F	�轌2j		ѣ�:����DD���F�1|g�����w���$����Z�Yϳ��k{�>�i�����rp3\�CMM���(v\�V�$}Shi:,�Ǝq	h?R�,a����<@�w+��˞^~�Y��y�u�c}�8|3����"�������&��u��b�����EBڙ�[��&���6��q�0�
u M�������OK��d���)�E:S����������H��T���T�rn$���&3������A��r'_2�f�;����E@	ol��i��H*?�ϵ�8<c�C@�Q^"�r�e��� /mO��լr)��T�>��K��cb*��F� ��iF��b3˨��$ٿ7�l�>O��(����e�"��){�8��u
g̘;7&oʝ����Өes�FE�I�<$�[�?VQ�ˆ�ݕE#KF0��Ύ��ܥ��J��ٖU� � [�@5���1�~���9r��x����WZ��3�5Q�����3|�j�����>��,u������Z��q�B��d�\�ݬ�]3��-���x��kxs����!k�U�P���hy�����F�п-u���~�)옱IS�Qhm�6n�@y��n$�8� Y��v�&HO/ �'/��]���c���w`)g�ʉ��i���Κ=����2��mZ?��� �������i@Df�2���Ӏ;ry��z���$g�X���-�W��:"�h#�&?ߙ�������;K�}*�%���خ9��F�9`c��ژ[�� �Gt�<��,���jp�[�:B�bW	6�&��������"�Z�����U��r�	�[OB��	NǛ�%٦�l�������V����,O��	W��u�W�S���v�X=_�UsLYe���i�/}2���j3�+�UW��лL:f�Ժ=�dՠ�����z������b�!���:cG��5��೏P��~�a3 ���.Vb;@Ѱ��ү`������b��ť���:���ve�����]7N�3ڞpl�+K.�sZ������rle�cڱGH�ja�H5�z�f՝����Dӊd����>w �� �hkk�T��r6�`g��|*�w�&D����l���O��r��񟞤��PZ_�+X����!d+ۂ����Aɉ��r4BD"����u@{�'����D�k� ���.F�HA>2����#�wL���fL����2!6eRP����b/�gܸ���J`����W?����F�p�/C�=����o��-W�!6�ӗP�p-L��UW;9�w�LG��ГXXl�W�F���wܢ��'�li�6{���Ue�욫ty�yi����0'vu���*AVzF@"��L�|.�^|�_O)�b�.
��ֱ/�@*��ꪏ�;�/-�������D��`�3C{ŎP�:U7��������ғ��yv)�9T�/��~1��p��Q� �o@W�Q������L]�C�g�˥u��{�����:y�Z[��MA6��??;�-~O�	�o�xC��|Wu���fZ����h\0��r;Gެ����� eJ:?o�o[���r��5FFGo�@)��}F�{���9�����/��բi��N�	R>X�K�TD�t�� ����⺳M��O��Awc�_dOW��~�1x#����2B[��E�	�RM鞤b|/�^'�v�4��y!�n� E���	����t^F:�D��;`���)�=�'��6r1�ɘ�
5ߕ-��\7���%��}z�����]C��s.�2�@�:"�R��U��J��g5��������1R��s>���~;�����;uq��������C�X5h�1P�g�IE����X�>@P;#O�h�7sŉ�IT~6�)]�?y���Z�1�Il��n�����e�_H�=��k��Baς����u(��R�`�~r���֫�����j盓�c(.���B��>~���Eb(���8�(����!� ��O�j�Z� ����"� �_=���G��Fyl6�L�Uz�R�F6��M����͗+���j!2��
2��#��u�����S'~�_?-��q3�qӕ@���^�]�|<�G�&]
�C�WG�P��@��Bb����Pc�Zm:
"u�[�~����8o���t�$�b�![_H��-�!z�=�H����\��l�U�`"9���m/�4�E�!y���i�3i�;<
6��y�ɛKy`\����Zfz���@���mƢ��{N�/8��~�H�3��1!�b�����%dMz���+ש�*1͔2z8�@g�����B�~ҽ�Y��s�#N�_�f�Y�6xf���r?o�ȫT�K79�ټ�l(�c.`\�f	=msM�Oz0[MbD�.wa@mu�K%�ѫ{A5�L_�ѣ��ӗH_o=$�lZ�ʅ]�k+�s���N�_�#<���f'���P��|)Mg^��}/�@·C�a�<A��Uf��0��[E��~�Y�7��Q��L��po���wh}��3�:�-.H� �u���%���9�;�0W�u'NG��
��c���l}�|�6 >�'d)��?�L
�l>2sd����3���V��r�L��/i=j��z���+e����R|w���X�؉��K@'����u �/Ǹ�!Y�:�A�����'�a�l��}�#�ԙ�>�T1����3�e?���9��h�}ޟ�FW��J*�3�[��	�G������̣����ʹ$,��'�TD�x�Z�9Ƀ:d��zZkNj�d&��^����#��<�z� n�Of�'�]�]��M�D`AC��i�a�:جx�P�q�to6��y|)�B���f�Xض����q�q��G4��Ia>�P�����Hڅr��,V�K���$�vV�F+=A�m��oX	�Tn%����2a�b�K�hW�����E�� JȄ�o����!�O��=C=<=��GSJ�m<y:���##��:�dw:sOw�� G�Yq)X��Y�Y���>��5
t��mZ���Mm�y�`�JL���QJ{gδ=H/z��~��N�0��z�7K��d��:[(�*�Aq1�p�3]�D�g�|�1��?�ЬY�յ�u_��_7��H��Ɣ����
�d!��ۡK�L�{��iKA�M�غn�p{���7��Cْ�ly�;b�a�9�Ǖ�����յ�H�9�ѫ.�Υ�1���yw��@X�c��0�}k��Ņw�Kh�QK��N8��y�ǑM�0&'za�k:�e)u4�5Zo����*/"���ĉ󚫘]���h�~�F����-��;Z	�쿟��� �ˬn�˽;7;�yGH�o��JD���Rqܾ]�О  o��?Nf�����`��I��T������/���)��	ɵd`
�o'W�ˬZ�{D�N,�N��Q��r��H���Ɔz�ho��?fo!�/�=�V��ǽ��6��r���t��"�߯k��t5�f�s�p���$HX�m<��j�S�a<���.Ǣ`y`Xa�)(Y���C:�[��$�o���V�s\����{���/N�r�`���31xnP0�{�~V;�u�Sv���<�t�a��-�tMY^�鮋���e�K-���s�F�7�����x�Ʊ�jҗ�*�.���
Jj��F��0T
;�à����x�6�t�SEE�����1��ưHb����ς�t������]�2]���m�k8�[8�7��e�O�Yug��yʘi=;��bG�:d��U���+n?�'@"�e(�"�$/�q��ʧ�Δx�ୋ?-��j�g�S�<��lӊ �;�f�,qD�+���Н-oUg��*ፑ����]��ט����{�W�}�sfF�|�������$�s���!�
;83hV�*y����s��c��s|�S��sN�2���0#p�tk����W�#��tq�X_� �}���DT^�8��H/���{=��7�%���I�z{�XT��=�}�����E/6_}��k�Ԅ=N5����������&N�A�><�>��']Cj�V[LWb�
5S@n��TZ�\D�-�7�V�_�n�,[�Vb��_e���l{;<��񐃋Ke��O�-7���a���-L�qeJm�陭u"��붮.A�G?�Y�V���wY%�<�1�W?:$ZGo!������pΕ����:.�����IU���̖M�2������s�&tl�."xM0��	�*�3R'H�|�Ukd؍��mA>�(���Z����gT����F�|��3lK�O.h�
��k �\:���|j�SR�v��^���B�ԗ@��������]͡�-�4��5���ԯX��J�����4X�-ɂ~�#/���9x4Tb���
���v׸FP@"�g���6�,��G���)E��#��Md!���<;S�uY�ʨ�^���K4�5��٦�)���ڴ>�p���ʼ�F�?X��ƅ8��9P��ߣ�Ppwwϋt�C�ns4m�G�N�.�Ү�����Ė��������ܒ<ju>k�>BM���<����׋���y�{�C)hhh�.��tP�_�tiλ�h\]X��d�D�W8ߙ�<4^\R/�xp9�]B���͜�j�P��O�@-�+�Y�Kx��J�t�O��Hs���o����$1h��W�b�mo{UX���M@Vk�k=m+r>?���qO��;G{�z�LO[��봒.3��o{�.���Hr($UD7|����\(���龗G��"���b#h���wm�xv�?y�,�I���q�Pl9��~l��ִ�[�:BL��	}q�ی�R֠�/���]*�[E9W���wʹ_�8Rn]f�5rX����d�q�r��*��_�����NN%Iz��RSI�u�9��RA���21P�4�VbP4GoP)՞/�Y�]V��QF+�c2G5ʱ8�� ,R�f��*�@F�_��$�/�V�F8�n�m^7��W;�_���z/)5Z>Ɠ(����^ĸLYn�-(�Vu�o3�����jK'a��)X*��N�/�C�vm�89��Zi�ԍ~M^P�����=8d�6a�矬���:��rqю��	ЀJ�K��F@V�	
j��/�fC�5S ���	U���x��$����8��֕Í��r �}��Y�2�Z.��
��'�]z?G0#W��ۆj׭���ƊOH�7����n��6p��q^��^�ۄ���T��c�����VUE�r�z���
��N���n����G�c�W���]�1��� ��ˇ��}�ӎ\'�ãD�A�׉��a��dm_*��HŠ��3�-�8�e� ������xM�^��'n_c#~��QH�:c3�t3�M�[ZZ�%%��???e�uk�bZ�Q\��L$�D�f.e�Pe�3K��}�٭�㝈��������q��D��Z��:��^a���>��'v���|�R�o?�qG����ӭ����s���9�1��J�ُ+�ô�_���hy�sv�����x�ܓ��tL>]ʿض;����3�8���~���� -I��~���|O�z��!�\�gG�m7�����m�	�f��Q����h��qz�Yp��T��������>�9F|���4�E��B{�5�1��0�9Թ��!���s饱a�ǂ�*�W��7����'	B��f;�ʙ3gF��S�����⮑�c�Q�������ǥ���ǟ�8����pIK��.z�����נ�m0e	�J��� �~�F�O�?.s�>�T�)ڕQXyy�U�mv�]hhڜ.���D��M���-Xg��V��&]�Q�et�ː��!��u��K�(��f�ޞ1fL/_�u�����U����j}t�HQ�ESI789i ���X\�a&��,yc<-8��mn�<Qo����i?��~&��=Q�:�тi�ı#��X�C�K�b3^ߖ-�h����;M�cD����K�Pf$�C�l�����\�U�mŻ��'��}�U�;��T��|M���&�u�.>d4�dCF�?-m�d[�fY���"!��%�Vrq�`o�tC�zld �R|�m�g��>������=�_(�QE�_�u-�2ǚ��E/�p,X����U���&��"����6OF���{��،̈�1��]�����堽z��QE��Hf�t&���O*OM���'%=|�5�����Ȧ�c鐏V��$�d��� d�g����Lnh���N�5�8�Μ|ŝ�}�NM���Fh�ЋR��	�!�jê��:L1�N�E䎾�=�R���WN�(ww�����d|�����̭O�:|?�)��1����{A�X������-ۜK��[���HMc�~�d�:�4�UE��uwqj�o���<�Iʢ��_�c�Ν�[Ge^m�,i����}��Hs�Hs���J��H��2�ˁ�g���u��BI�UTԝCUC��l������A�`����1f���`*�*�[��@B�j�&r)��A�_�6Ǆ�"fjD�{���xrEJ��0O����x��~a?�{���B�^DI��j���ZG���GJB��r��>��y�I2g�{�K<3����.c�15e"�/dm�)i�EV�3�{y��;����m��4�W3dQ���:����d�`8�ٻ��6���!�����|�٫b5QE3���O�I�@�>�O����5>5[��Z�ؗ���XjET�f��Ï�2ߗ����98D�8B�/�L�v�/�.g�����5�<S	m� �)X��ɟ��x�fʹ�6�܅{l���l�/!F�t�)�3�lD3�4�q�Z�!1 Y����=�5PupH#���qحI��y}�y)��(� �C�Y��\u�t�D{�ã�~���(?��N'Wڷ���[�s��JU�F1]95�8�������27���G�U��,�(�B@wҶ�Y��?�Wh
@SPCqq���t�!3�oy���������϶2���c,r�[�bD�]�������56;l8�a��\ـ]ԳJ?V�N�W�ܕ���i��+�R0��� ׌i�h�t)�j9��#t~�D�kR~QFG��tHq����U�E�
YjI���������q$�QWo�������K�<��Svo����Z�>�aѧ(5��S�,�\��l:/-��iP�xR]�����to'�C���^K?��,�Hn�l�{���xǠ|�Xt:�e���-_I�:�2�$�gt6�������C�]�0�j�ēw��t����Zwr���m��cG~���[�j�d)�t�.����o��+~]r�1Ϊͭ6�jnL����#�k���Xkn���G9e��W6��<<ʻ,��uK���|�fG���g���&K��q	������p���"�$�&t����nRl,e.���bG^_��7K]͘�	�7��.�قNc��m餿�����L65�cI7w�I���3k�p O#<�<@o;��@dD�D�0��d����`R�F��r��.�~�W���h�x&�9{f�2��F�������O�ir�V�� ��=H>�Y;�}�"D�TGW7&T���/����t�8p�n�l�h���U7x'>4Y��%�_Љ�ED�ubQN["�Fv����k%��<M�oտ@1Ǆ_5=�s�f@"R���VY��kz!ɿ���!9%�C��,7F>��]��xA�+U�"ό�Y$��r��ּ|b�����^����@�#:±]�n��/��z�ω�Io�C�/E�
6�/����Ѫ��e�� V�c��j.�;��4�,WEe�}�-i��+�w�ܾm�b���{r���VĻS�o	��>�j=�»Tt>1<D��F���e��������;��OVUS�]�h���"1?l5 7o���/���kFɦ��_Z~x�|r���f�:+�Õ��8���t�x�	�j��15nq���K��e#+��jx4A;V�ߛ��&�G�/��O�hȒ;��x�����h�0��0��7>9�3�Nءi���IQ�$�җ37����>�H�y��Z��x0�c����B����\���sA���!	�-E�X��(�u��Q�j�0"��2�jR=p��&l�g%륿��bm�e��������
����	|��_`�P�Jd��cծC��W������|�a��_c)�v��S��i�\I[��Y֡,�s�?n&�s�Ҹq������vTk_a���k��?�aU�����e_F-�ņR0�O��.�}�h��y�q�ޚ�C:����9��f+��w�R���Gˎ}���Y�E�;��NkM����֠~� "or� �S�\�E]'P%����sZ߹��Jn�е������u+��4�5ռ�<��F����s�n�|��'��h@�D�Y.��W�.�A[Y���}�&�dh"��E���ݘq��k���c�V����*g$���yɪ��rT[�8*H���<��-�8�ɴ���3�s�Q�7M}�5���#�̖f�V�<��������D����dpWW��U7���}(�ၳ#��%~�Sj��̇����^�8A��G��+W5����;�Ga;L�F��S)C�zT�mb�%��K�.�?e}���E���NcDQ#��whђ��>�:�fu�P�l�;������H��m��d�ٕ�C�VF���.�d�e�)<xd��$~���Fi�ih�R�vx!>]�0p�p�>ki�i�X�_��rr�E�ބ���y>_:�]U7��A�q�4��o!��v���c��j�G���ud$�J��󸜊���(Rmc�N�w �(赂<^��"2Hg�4�X8��^�/���s^kK��/�A��m�?�zL����kYû(�ή�ޙ	���'`������M|wbP�"����R�����7� ���%�MB������(g�3^S*�g��>�����Z^=y��b! �����Г�*���/�8x8�Si㔬+�C
�?��~��]:� !�՛����p��9v�9��P�T�]���-*��L�}������J�#�!yQ�r>ٱt�;c|bb��h|�̾!Ԡ����z������&7��2]�J߇F�}E��ժe&[ԝ(>4�$Vr����xA]�[�#��z��w}�t,�|D����L5�0��z��X����[���7��y����k�	VRN���Z%���|'d%��mX���2��4�פ�3g(���]�h����555g$"s^�8	3�6;
�� �]xq	�%ZZ�}ߨ�D�0G����l�����#�{c9(��>@3����%&h&�����r4������wk�}�,����ic{��/����R-�X��k@/	���	�U��L��ďDwC�s��.o�i���;�6$�u�^�P9�:�\�>��\�ߎ����i9�]ψ��G�`d��B�W��O��Yڭ�yyKyF�C���x0��G���w@����d�{xHC[[j��Y���0 B���uץ-k�G����EkCw������\�� x� ����<�
~�l�bɌ�f��Ī�8�;��
	e��R&��C����׫x�S#D\2;E����L[9��پל{ת�h�In��]��n�v�J�0v�(�T��!��o���a�z�u�O�Y4q���,�W�l�h&�C��w��.���X�� ��RF~��P�	�1�ߡrq/��nWz�[-Y�b���u쇍M>qZb������Q�?�l�=��k�k�z��s��Es��d}��q�����*={k��NS�^0����v����k��aCٽ*����EƛR$��3���H�dv���6܂Qeʭf�H��35s�5���'��֤gX�+�K�(��|�&zC^˚�����W)��g�v��/�Mv^.�/��1:8"N&z��1Q��W��Q�R^H�Tia���y�*l$�5:d�����<L���O��p��b�܈��������wBϠ٪^�������Ya��'���-��}��B�k�>���� 2�u�T���`����l��X1�oN����m�����շi�$�^r
�܄;;��nGN6���$��ƻyqm�^�Y,�m19SA�����:֕9��5�3&��Y�+ �ﴎ�Õ?*�=|�{s�Ņ�Z��H��m@���<�x~��$�����T�r��Cf�k�G��.�m��X�NT.�2�!�����Ȼ��Z�|M��A-s`_����:��z���WM�ȅ��iz�rgR��ח�9�V����> |��œ�$�3�^�n�R�E+����g׿�L��P�[3e�g��j5utt���_X��cŇx�� J�O��ݒ)N��	k �I��Lr�_�#����2H#�� .�s�UŮ�3
R(}�����Ύ�~�����Ł���\y����2㢣�gv�Μ)..5��,.f���ődǅ�/:�.�	��+�Mb�j>�Ӈ�[�W��sk[Y�R�odߩ!��H�j΀�K4C��7�-
�!,��ޢ%��:	�?��<�_�$5}��;�2w�!4�����t����s@-GC|��R���斫fL���/}�����
���;���]����"���N��`t���ւ��Ί}�*Yf������BD��OR�����70��z���aÏ����~�-��|��#�w���0�ٞk�A�K�O�����z�*t�h]�-�圛��Gj��qss'�"{ӵ[J�2猌R�g�PAb7}g��Ƞ,�Mu9~���?^���У�|Y��#���R�ȩ��FMӱ�;.]+⪚k�}2��kM�k]�C͔2%�:�O�oIޣ���F�D�w!rB���z�8�[�!�8!+靏_�W��3ͥh��n�<��J�e�������� �_Dv
��ym��#��@��mq�$��";��ؠ��t�У��������E֦��O�Qۏ��&}��P�&�Aa9�+���с
�r���.�&�ޫ��tcNEj�Y���;�*�EMO�{:���l�;v���S�~�Q�%m�քowpJ�8�� �f�$:{O��N`�3���###�~����z`y�T�"�ƌb.$ޓ��T49�!	���ڵ�� 9�	Y��Cs�Ԏ��SC�7Դ>U<��IO�e�x���+R�� �>r����,	&n�[cכ\J`J�3 75��Pq���|Mgj�V�W�M�� ���f�z�^��#s��O&5�b	X���@��Cps�i����5�/�i����,���,iP�x�2�	T��4摅�T����NrH��L&��tU���_���hL��}@A��������ؒ�nҍ`)��w�F�(6s�����U�A��y�\K9?F�.d�[XI@�4�i�"]�t���G�ǍT�Yu$Iqv韔�JZ
�K��@�f���_�����{9[��$W��c�m�gt�ҿ����~���RX�QB^Az�N���P�mr��F�K�tW ��g6�)�]�;Z�����!�1�*���R'T�4�7��2A���Yf����U4�x��-EH��ڲ29�rnboa�ǅ�qii���;��H7ɣ�;M�t�q�+͸ޮl�#�v�i9����=*��AX�[:�}��a=��wX��x���rK��x�U��v��H#���L��!�Хn)x�?^ԟB�A��t�Z3x�*�����<<4�Ę��ٛ����lP!Yo�,#�7�1C�!����?���O�0
���f�6�j������
 sO0�C�p|||^I���R�b�^�W=퓑3]�"���u^v/�N6T��S0<P���e�=b~���eoAf�F��ۢ�,/�bV�V5�T�p��%J��xV���b���������ޮQ�؉���d)�k�Z�+#��O℺zw^!N�%aR��K��,�]=n�\�,�gB�]Nza۾�vє�x�2jk/ 9���}�k&��!�22�_�q>����Yc\�ɔ�(����7V��E�N"���Ve���{���\r;E�:��ijb�	����7X��5�N#��8t��&%be�ߘ����i������"�{kb��C�gY}~|��KNf�t�-���r~G�f<Osz��w/G&-�z6@�^�'��UD|	�c���I�|e�24rz�+��v[q4�u��;���/fwC`W��:#v�=)XM;
OZ�ф�Mdp�Ez�8s�v/ �^\1�11���9�μS�*�j�=��P�h�ڰqc$��|�0a1Ǿu��l�]5U��W�N	UvΑ����t[��u,�[��݆X������
W�����BP���t�g���Q���������U㓖�55��[( ��'𛗺��+@ݷ�oxvC����[i�h��W���<��$�WFrRSS���)X��
q��f+#J�MG'`ƕܽy�Ъ}û|.Rn�����s�c	mL���O{遑���"%��Z�MNr��� U� �	1��P �]<��]{�:�U����5n��w1���/��}�3�N#(�����G)��E`���u4�쌠���#g+ƻ�M�6���6�~���/ U׹[-��Xa-�n��,p���q>��H�����p���n���|�흵�#y�I5���=H`�烶i�x"Vz�{���*��5��,��^+�0^���x#���GRK< �K�H=��0}�`��M χ�T1�,pn�6�ɇ}�U0 �,�*��r�i��7��'���O;��"����:SD�#o�N���?�k�=�NEacv�I�V(��i���Կy�rL)ҮP�iP�����,�95��3�
����j�2��OH��Q���ps��ߜk����5R+.�&f�o�q1x��O�a�������uX֟�Ь9nv�9̩��`���g��>�3*����U0@���5�'�).O��V�����K��Y
=�d� lp�o6�c ���1(�yu�j�-�_`�|"���׏��ju/������P�jDh���r1L_ۨh:�v4��"��o��3����i2
����ZV���Iؓ��	������L4����!�F`���Pa�"`��@����Eaq��*���0��t�08�{T[�2����7�Y��hh����P׳��^�>��p]��O��6I���З������������ORR  <���x�6�]�/�֩M=)1l|q�AV�B�x�`GMgR�˳(��㛟��N����V�.�/|P`r�,Z�򌊒����?E
i�eVQ�� iD�R��7��U�����c޴�ǒ��_{�3_�$4�M�]Pq�藋�����'X.��l.�`�տ��=l�5!N��2���^Q7�F|��+V�z�� %��$��q�����3z�9_��%�)ť��a�7P�������������O����M�*��e�j顱�����ر�<S���4��Q$�֟�>�̖r��%��A� 5���?��r�Tc4�՘:����B�=��Ӕ�	c�C���}�(�K��a���;���m݃�1�6f�'�������sS=6�B9��Wd�+C|�!  �\n�um`���QJ0Kg�)����u�?��`Z�'զA������DK���֖��;��]����þ�7ﴚ������0m�����b9���(�jĸ�f����[>z�+�7�5w�D�r���L�
'?H��4u��*�m��-��d�d�q�oo�\\�"�Z��n.n���u��\�����%�_��md��H�zθb���^C\ؚ!`(3@����6��/�XT���ݶ�8-\��AXr����)��+]�����bϵ���3�
);�*v��n���Ou��I�T�K����'q*����)o�[h���E������h������N�{�������I"-}\�ϴ߻�x�/��ل�#�]��/�s��\~���H�ԗsw�$�.-��h3e���9�.��8���3��o}�}W�ǜ����+o����I]��HUV�c9"$9����C��+�� ����
�̢1>�Bݰ��d>��ޙ u����3����*��
B���=����r#D�T�j:��3������*��H�B��V�p����.�8�����ֲC��ˁ���*!��:�YG�(����s��J��h��K��9k0��_Ph�~h�,ޟ�:��
3�0+%�u���?�`ʶ{��I�V�<��֑$3\���j8�t���m0'�G��kY�!z_K+�G�NDa�N����4��`^�%�>V�r[i�r��7���i��yy��If�p�i@x-��ל�O�a����Ik���ϥ�<��,%y�or)]}���__c�+?t�����Z�qc�&�93V�r\�0(:�5��Wz37[e��-�N/��=2.�����Â��}7F0���-�+;�����jp����~�0?�=7�G�%��0��s9��Wp�6Y⟅��;p��n)��#�==hɭ2��ΟV��T*�5�`�� ��O�ֳ�ʔݗ�̔@�K�����ۼ4�l�s��|&�IXE���8�4X�~���ۃ�j�G���O�O��&��H�ܨH��L�kC4d�/�g��~¡�?)R
�rf���?D� w�2V��[4��R<�����2�����0{��6����f'�8R5��\	�/Oh[��rD�E!}���날0:�a��]O�W���7}���v� ʎ[�o��n��[���yW��yL�Q`��
�����s���6�8��*�y�F��
��ǡ�yx����H6ޣ��M8��J��`5�r�5j�a�.!!�ӒX8�<��DI�wI/(�s2	�ș�;r�����P��	fɌ�����{wK}m�����Hf����%�&/:��F����.�JQ�.�߶.���xm�[���U�%���G�{���b�fC�%�3cG�.J�U�m���F�8�Eݾ�c�W@��6=�5c�_��ud3���+8'�$�R��4׊�I%Nن?#ȸ�]�9Z�և��<3��k�����G��=Z�ų|��s52b�G���6K�(g5��KS&1ς\߫x|�ٽ�O[��kG]--�a���s¸t�v�oL���+�#���˭/�3�$!+4;�?�O%��ʹՑ4�@�U��߫���䴥!�P���{傣��0W�&�FE��{�+Q��<-��TӶf�	'D��vy����'ɒ��DhE	�x�r�sS8�&�p�IY��8<�E�}�.�����������^�f�h��< ��uҙTa������ 
�J�Z�ޮ����b[�JƎ�TD��_�J)3Y���.���6�~/ّ��n��B�.��߆���BKK)rM%�$N���&�:C����?���'?[\m?����0���Y��;4�6��˵6W�VŴW�{�s��r��۰�f�u�fʀ #��8�p���8v�+�ٛ�k)������~�2��?09a
X���Y�$��y�&Kʺa�V�����aB�k'�4���ҟX�&u*4��;9�z&!�$��%n�b�,��,�^�d����XN��Zxq�WeƧ���IH�7�IG�����F�K�����Z��V��F�]RsAc`�O`&F0f(���N;9x"������x���>*�e���O��{@F3�Xٍ�'�+�+��kކ�zї���r^H�3_8	<���ݥ����Y��{���)�G`U+�+y6�������uIj "3TL���=�\>*�PZ[m�\%�f��䲸@�k�?�Rµ��^�uf�����|-s&����c28���_Lr�W�������؍Z����U�Q��@�L���P��@T��;�ɺ��Nʳ�5L��h���%h�a|��D��8,P���q��0q����S2�vҌyZ�<ه�K\��_��3�I��D�o�>�`ܔ���#�S� ��R��]m
C��7�}0�ZzntS�@e�i�7šK4��.��◙w�Fy�{ͩ���/�Q\�����ℯ�Cр�A���O�
��3��dYouV%{��6�b
�ħ��=�XT�ֻsR)�[^�8i��į���P�%�W^�6�p����E���Z�m��nz=y��֋�,���P��!�UVQ���,���;<���w~,���&�n�}��[:�+	�Z��T:"���0����H�9�#'!L�g��Uy�:'^C{��*�{��dv�#2hu��ׇ}�I�Vx&���M����ށ4'��Bl�+��>�DG����"���<9�׆R�9�Y����%$vɧy��LW�Ԙ(�0ʯB��>C��rS�V�y���H�yz����m�	>sԹ�{v�@c��-� ~� !��qZ��ឬi�s��������dZW��:�ˀp���]!�o����XKG����zM��a{[�� B-�/YSAu�P.����-ﾸ}��@S�9]:;��[�Z��^�?=�[9Ғό���Yh�9��I}�/�`�)%�7CGK�Elg������8ΜtO�+�3�$=
�-LaՉ��ԍ�r
&)�C=Ce�(�g��X�Ĩ�#�JVb�1�9�G��t��

f���Z��U�Q�$�R�p���şh�.�� gk<��Q����*�:���gf�A�qVV����*����M��k�v溎���g��[�<d�wSwN��R�u=27�&��Q�؁���Ղ2�&r2
�I�q`6o"��-�#&�+S�*��&��"�������j�����|aQ�^��Ke"N�Q���WH(�.���(Ֆ\M�G}ڠ(:Yf������9��۔�wZ��˅v_�1��G���|��	�[�h)Ci�'+t����կ�N87{�����HKP�)�^�bFU%�����ɕ���d�Q$-.K��8+�#�v�6//��*��2�-ζ����ssO����L��9/(��O�P��e���T��q��(�0�,�`ʫ���A�E�ן1h��ge��I����>Y�w��^b�W�f i���ӭ/=��T٘5�e�l���)KƔ���@�m���5�z�ZD�:�җ��|�Wc?���k�L\��v��\���?zu
?��wF[�yG�֟�	�����Rº_�$lF���5�����;���Il�7}���~��m��9�o�bD�����(����7�&��F�A�����qp��'=�d��/%�Ȣ]m�F �G�wG5,oGQ�!*"�{��i�A�Z���T�H�ޥw�.-��	:�@B��z�����ywfg�gvvv���)��4���#/T?��YP?D�܇'܇�W�)���O3�;��\�j�Eji0��c�(ƽ����E�G����8�8sD��kܝ
�w�x�z�����F��{p�'K�Ҩ�㒴���
E�����q���3I�P3l�}h����R:����yVN\����ٖ]�7򧔜��:�Ѕ�������cM�Ie��5Q�k'��"j'�Is�a��煗!��nV���I�e+}˜��>/�fO?��}C�$����K���*�?
j�p���rY�I��{�Lȱ�\k��@n�f�Tm%W���ǳ�T�)�% [s�#ۋ��-BF���y�'Di��T/����m���WV�g�?p�C�]t{_�y��7K$���
��cb�t��p�ְ{�w�����))��d��g�>�o-
�g�J=�z4*o���5ո8��j�H!m9�#���&��z�).������xJ~]� <�ĬC���B��P����U�`<|��)j�we&��UI5�a�{���Σ���f�>�M��w��|��w�l8$i�
��� ʨ�A|�� ��X�[��z�?�76c����V���.J��y���ā@`_����l&��ܜj]���CU�_:)灱<�����,�;��'����''���e�����)ۀђE�)^J�4��i3.�&�Tx������p��^(�Y����[�/�
`뚷��5�6�L��I���zF+�㮍�8���aIj�$V�bb�x������m?��ST�U�ح�)hv-�b���r@$K��K�4ur�&C��F*�yvX&Y3�j�FuI�����]�{}�粙��Gռ4������߈��w���]�ﾨW!���~C�婟�'�:5��}q���r�Y�`�����ƲJ�E^����aB�>�8��܍%<5�K�H��vSf�P�rq�����q���%.y�l~N�l�$Ӄۚ\.����+ȣ�wۗ<��q������#:�uΊ`z/�y�\]ui�%[��ϱF�27�q���r�(m[?�^��k�GU�<��b�sdEݏ�2�&Ҕ�o�%��~PQ�H_R�Ux:`5��A�奘������3j�ۋ���25�cc�M}�J7��^�5�0}� _[���K.�ރ*	��0?z�l��䤞�0�K�'�{3�P���?�����0�i����]}�&�B�+�	&��5��n\�/�)�m��&RFiT��n d�F�ce�ԏ
.��[\�0��Mc�v�l�(����f#���a1����1�
W�v�ZY�F§���i�\��s �������03�M�'1��uf/����Uji�[������5���6L�¼�ST�m'/d�}�����{��wĿ|��'���@5���+�b<�J��mF���m�Q�}�	�Q3���2�d_��18��0�Al��$�z1eĉ(��R+��B�A���.�Wy:ځ6��?quƓ}w�A�e}�Y�)��]�O�İW�S�=V�'B��F�d�at^6��l�{�o+�w?�Y����y����>���cͤ�Ev:6����>�����(u�2\0�O>B���D�^
� ���6Afc=�K�폸D�y��?��;E+ʇ�=8Ӓ��R;���V:�⺴}�_,Z���6c�� D��fK�ɱ>�����{S3�6�"0̋�i�U7�wu��[��r���MDQ�_��a^6�o=͐��c�S�{k9��e���&T��e��>�J�Y������zñ�~�K[v>Znt{�s�g��^rޏ��~��:�֧�ێMv��k	]j{����G[]-��[x�K�A|(]�Կ_�c�Ks����Pţrw�#8tw;����<'�J�T6��U��~�Q-黁���D�R��hco�:���q9�_ ��]w��V����wZ�4$ �vzf!_�����7�h���Gik�t �AEW_����tY[Vd�����Dn7���pp�M`~E��n�O�,'��#{,_On0�u{`�ǈټ�󩔟�Gʵ�v���
��8��~،��:�����\�fk��j�#NU$*�|O=��b����'��J��9מTS~@�]�����:O�4�ɴ���v���M�g�mi�̛�F�Yٙ�Q��O����\�`%-Q2�pG�������ff�t�(*�ғb��	�Uĩ7,U�y�2���gI��4�K�$�{��ߒ��_x�pZ����B�D�v��a�
�V�5�~Â�&p���qj���W�;5mJ��;��.�S���>FO��d�Sֺ��r?c��գn(+ۉ��0,}��@�bZ�<^`�J��d��f�壎q�� Y 6Vx�Jᓐmi�+�&i�w��t����j#�J4�WzȊ[��zwF���R#�d�,ҧ۪�����%D^�K�� �cU^��`���@|<s%ӵ��Y*�����MU�WuXQZ���y'�S��t�z��$� S���{��Sw
��F߆J4�P�6�-HY�k �1�J�/.-��~4v��7r�K�]������1Cnh�Ä��䤈,D���r{ES\��p\]��XW������Oa�vR�`�~��C�;��>c�'HN�ʉ�G�p����O	Xa?��x��Wm��l����M9� f��n��q������c੻N��GH(��m�|-p$HQ'j%��s�R�#]~p$x�i1~F�v��J�J�u�ޣ�ʛ���b�[��'���M�Q�	���h�xz� $Q�h�`tZ���k!�O�F�c��Im=�S,�`�����;e\C����]H�'EWP�o,̜z8{=��Q<X�ص;�z����B�>_o���tI�g�6�S�/t��ɴ,m��DPB�����0�ǌ�M�T�,<be���'�C�<�Z"�]8����E��wJ9�L
���z���Y�B��e����
k�s�H���-�kዙ�o6'�U��'��J���Y�#��d�bz��j�9o�.���|���H�E�ӝ���x"���
����UڿJ��_��W7�����'��w�,Ʃ�md���� {J�V��y��o��]n�r�"I)�ߛ�`��� �ɴ��w��
[0�ri>N���k.�u~��m�]7������S�V+�29��N0ǹ]*̬}_��7*ot��]�="���J6���K�WC4�e;����s�GFlnZ�y��پ�󝡮�n�b�\���+�=MK i3:�v�����~�Ej�:a���ꐫ�x�;<���ߴ��:E=S�r�ޫ�ې�;��Ϲ8� �(���F���x.�n�א@	���ﱰo���x���:fA�iԼ��x�"Nx�gK�7�É+��A���F���V���&�V�M�����6p�US��G�2���<^L�Ok���Ѫ
�\Vr���f���0菸�2Tb#ۆuq�c,<�Ⅸx�����l�.̱12�DwU���220��Ot�9���G/H~5v�uҦC7U�_�[-����M��-��yĚ{��eD�lu�zoEj	a���Z?�k�ۨQY~sn|e�,�(U,��CL���YJ���@��=	�e4V�h��vJ�,��-�� �G�Q+�
x&��K%\��5������P�/���X���g�����W�,*0�H����-�}軑����t����M��|yI#�B�Z�����'�;���8�Z�y*�n �H�*���P%=o5�gl$��ߩy��=�%�T����L2$�zq08J�"��{�;��pmtl�z�vl|���N�B$5�����U@����b)��k�Z��
�	:-'�Ń�ӣ����ǭ��ʣ���]"g�J�6�LE�jؗ�z��P��6�S��4�'�ږ�.�8�ԢE�oE�c��A�ߣ=�!�,�E05HT>��-��-1�D��V�8��Ʋ�O�#vA�-��|��FJ,�?e}{,8���92�zAd}y�k+K��W�o�<-��.�K�U����|?�`��y�~b��jgL��A#$�Fq��^ad���5����*��������^Qc��HIDp'p7���BQ��A�[g�C�{r�^�Gc�M���2��E�nyO��LN���~����B �����20cn���k���-벗�~O���k]68��~��T���"���-I�u���,,@J�G�`���<�~�i����:̱>7�]C�t������qY@%����m��a�:�� *�?f�oC"\�=���*D�ۗn*U\�7��G�	�"�o�/����X�Cv<� yF�\�s1�[���V��Z��O�c��fȝ�B<ju?`��L�Qry���R���y[u��n������m},���<(!�� X����ܕ� �U}�}���8z3��4_F_�?��~���K���g��d�=K��U1G^�� ,S��[/�"ڻ��K �
��&��_3}��/&���v�
i��iK�����ۏ�G��G��2�B4(����t'yy���bkř/�.���D��:���z#(��h>��V\2��j�jO�� q2�L��ωg�ضPѣ���>�-�x��pz��к_Ǖ$����u�	��"r�t���~�����4\}j�q�{�����k�Δ��XKy�CyQ��6f�t�nM�&dhh�������D�W�k�~�fY�l�;�a�0��8���Ɵn&%�8�NM��'<P_}v�?s���8��J����t6h�:�YY�	�o�G&pCȶ*���=���s��J2�z�|��θ��!Y$)��	.n�Y��8 �9x�/�	,���{m��2�k..;�O���H�����S	;)�DTz/��F��b��J�N�t�RW��2�㣗-�K�,��d8��T�Ƹ	����F��S���p��IY
���X�(tw��17����wf�W�83����҄N�{P�㎉K��+ױk|��Q���߱<@J���9J������,՛cn66jRm@$ ����5�)���E�d�~�jdQ��Aȇ(X����ht:����ΟV��*u��Xw+���n�/m��*�I������S�*	�Q���A�o���a�o�^|Ϧ����M=�t�������zuD��Q�X��K������eߊ�4��_ؔ��5�4���,�=ٴW,��k��h� ���<�����/O��G�>
e��;΅�����JW��;Fy���m�(�!���p�`�X^gae�L�Jf?ft��]�<�k�UꐚyՐ{z�0�f߸��2��:�8�B�jB��y\�#�? ��	򂥂�*a5�0��1��W���(~p|9���&�Γ���ԋ�4�5r��óhC�؍��|���Y�V�^��^b�]�q�l1�d"\�d:��P��Z�tO@Vc��+̷皅rH�P��J�nw���X,G��bf7�<Fp
<߄�^��d#D��=�+Ƅ�Nd��t�`�mr�th�/|��H����@\U>'{d�BF*fy��^�MH���2�2.pB�ۨhP�	2Y]]ujrFV�&u�;�������_�!�ˠ5Xi!N�������T�C;��o�ު���?�+�t"�"�Ht7����!Ԏ�}��t�{\�������H��ў~(z*�'�#����G���µ�{��r]�-���c�L���2�%MB<����:�A�Ҹ�9U���C��Ћ�D��X�_՚`s?����4�����;�sY	�0ϩ.V�/�f�#X�Ao� O�Z&�9�jt�e.h��OD���}p��qaA�rC5��ZP���u^�*3��;9EE����������f����I�&DW�>Ey��Wz�uK��x���Q�Q "�s��Զ�4�q؇cG��L#g%�$�+I�B7Mٷ��2抴�������cS����?�#�������N�n�Z	d��/Flj%@�Jǒ>Uѭd��@S��4�����m�U^�f����Ǭ>���AN-Z'�38�)�c{����	K�'+���)���/�U�3���ӄ�߀O{F��:��[E֚ф~],,�:U:��y�a�R��ԋ��.ʧ�V�0��DK0K�%)D<n�x�I�`�T��Q�Z8K��l�d�Ȭ��i*���7EA��� �;P�qS�M�D&5��U=�W)�$��1���>/��t]��+�#���Wu�nRN�X]-������ʟ��8X���X��(��|�[��4��̪���;�񱁡��GL����s�{є9�����"]��. ���w�(�\P�%<M>���GtG�L����cR�L?]��MM��h ?˽m������t��j��/�P�B̋G�xN�n��x�
xF� �L���D{��������~�!�
�X���߶����q���>����sӕ����qF�B�J�u���O��1���9h���>����
��������1�Wl	���&�%�-�?�5k�y�8�E����YŃ���J�ҿ�H_�!���"����	S�Z�Udt�|��h[C���`���xw�����	dS��V��}���Q�=���@]@ʗ
��{��`�?G
(��`	#�ٻ����C���R�h����,���
�4� G꧞rf
�L�� �#�8�7m;�p�#x�u�f�����*���]+y�s����cI�d�<F�O=�F����ؙO3�$ć�X�׭��+,����;ի8..���M�R�����z�J�Y9H�kJ�����e[��!�����{N'��-�]R���L�/�3M�݇s�v�_��l�g�[�~ֱ�>N'��Qت�����aS˙�����<����_��9j@�\%�v�����ڍZ���O�+<�ce�n�?V�Rcd0Z�t$��z#?�Ć���	#�ء�E���1�,��XM����|�0�����1)j��ZcaqzP�������Wn��C�<v�2��+)�7)�=���Q�xk4h��SK[�AU��j�b����|t:*��-3K��Bf�c��	0����{���5�/�nA͛/�����>��Ջ�`���0�~�*ӵ")�-�X���~���}�W/��0Y��c��e
�!l�l����Rk��h}�ξ�����ĳ��1""��^Q�U���ߠ���=� ����f�<taE@%��H������B������p�8���3��F�B�bAmՙ4�SZ���ud�y����$�͌'O33�j�Zeq2����4~Tq��u�G�4c��]l��M��!�}O�a��x��+��	�d]�;��rz/M!�Z��nj1]ǺΧ��ΩqG` jkp`ղ��EUj���/%� ���\��S�us�IL�n7� ԠN�L^>f-2nzy���tR����|�:Ǵq2qK7�����#���/_���|�6;����q<V����i����{.pȨT�k�>�`�_S?��|zz��(�N]I��c{��-�0恺:Y�S��:�,���\"� ��;,?����	�2g��si���,2�_�c��lm�ݘ�W�N��٥g��X[�B۲��O���;�	A(��veNk�aDW۽����V�85�y'r����t��Q�Dۡ��㨬�����9A�r�R��]Y!���=B6�k�H�i����`~�-q��s&�@��Ε��-(ؼ5,>_I��2��x�Ѹ�1���#���g$��K�Iڈ
���sE���3��6���g��z��xa[u��[}�B�,A�v��w�_��{��S�Jk�e<�������P8p�*Oe�v*MM�95����h�Ё�m��YT�x<�'hy2=����u�y^9�Lw��I
�9E�r���;�[O��:�TU�::�u�l����[��* ܕ�I����9YO�����o�s~��C���>�5�[�r��T���2�U#�#��{��8�J����2陙�F	ɛIA�RI��C��&�t�h7n��`ƚU��{�d<��i*����=�{��wre���x�����������d�
"�5��.k���o�Y��TMڣT��3
 �����.e��������BBd,�o��H
C*՛�9^�2���-����(�#zG����Bj��n#����ÛJbm=t�9Uboj���v��r�mtn�n��h��I�x�X���\ZE1�_��W�����1L��Պ͎=������*��Rg=`����(�4(�b�/b����<�n����ߵ9�1�����J��AYV֌��m6�R�O ��n�Jh%p)��Cq�����9�<NXg.�S���%�l�� 	g�|���!t�+�G���U�ǘ������o���cP��sԖ�t�7����?1��Lͯ/���xmf�eE|K�MH����M�Eu�1�������������s�7:�y�&z+��	���&�)I �a�e3��M��N��	�G�����yh��I-���n�)_^�.��_�N�HU�2Y=>�i�a]W��&���ӚX��C{�%ƙ���	6�Jes��!#���NEU��lA�J6n�gvM�5�1��E�M��,u��ӎ�G@��S��%���_�d�TR�=��a���?���ش�0T���Z]-���(JO%+��Sbd-�3�KV��f\\��ս]�-���5�)�g�k˺Uj-�$��P�����^RD^�� �Ewd�`�ը-b���\���K4mrˏ-�҄����Ϲ%���키��3inɑ�e��9�����z��S�f�U{euX%��H���zW�1w��`���T���#���2��L�x�X�m��'�Ib����u*�{���}s��������b�Pj�5!a�5��+e�#� ��'y��"�z�i=���r���8���
>��$$2���y�T��7�I!.Oj7�="�'��!�}�[�������CA������o�;A�x�8j^	�j�@��O�����7��d~�v���U7^.�)�oԲA9�'|�k7	Ս-���IIG�p|�틙�-t5��0�,�N�ڪI;>������`�7o�����C�yས*����5?���ϡp�>y�����n�xJ��J�9L�9a���Y�q#���m�d�FsT017#ci�X5��GCR����ҵ�KX�,�/�c(ҳ�p�El�+����Uo�ya1�"�N��������XA?�Tt�M���1Ln�Ś���篨A�:�е㙄<䗛�I��,��>���x��9=}�gm��ǁ �n8��.OLZ�b�BQy�	�=yvL��>g����乹o�	��d-�>j�+��٫������S\��d�����S=��Ft��gϊ}%ΐ�Bl�&_��B��3�me��DnI��Ԗ���O&k�#3��N��L�����N���de���Q~[g)�Ȕ��NX�lZ�q��|�5��{��ߥ����X�a�4�& _�;���ݐV^���d��{~)a|��G{s���"��x2.�7"��8L���FH�AznC������C#q[2*B?���L�����tt�n�X����@�&n�#�)���g�C�e�WbB䐈B���v}���6�Q����^v�s��1�TR_L7N�U�����uzs.�����ߓ5Q>���}g�4}eKG;o���Y���;�[���2X��� _UJ�O�=�v��D���#+=Y�n�:܇�oXs�,�z�>$��/'����&�3�z�魕Z����"w�Ǿ\�'����|��C�ε&S8�kK�|<{�g�M󹘙�!F}b��֒�B6��?�.Ύ�K���Y�|��[b���z��¯���o�;dhsⓖ���.��v���;>�1A��N�ط~�6���||��z��B�ήF �uos��{�\A���U]'�!{K�g�o�����a�#em�37��������h�7��
�j�	��:
�l��#�Z\rl��3ض:�r����{���M�K��_��sRY����ϫ��� lGR9B�1-3C[�ESDY% �rG���#/���*��t.�:�&ZR��s�� �X[�쯌?o�I�J��\X-7��7�E^[G�?ܟxe�f�N"3a�1�mG�(UD_jF�Iߚk�t�}3+e�FnV����>m#^�)��g����d���O�@FJ�"����1�7f#i�A
e�Lӑ�Sb�o����:?.�ن��kt�7'�֊}�uB2u���o!FW�!2�(E]���޸��0CȮ��zX��G��Ҵ�=�Zl�N:��S��w�����M�2�"(���x��DL�%J�K3�;S�������:~g�j�Z(��%'C�[�l0Λ����	�����Ī���/��7Q�B��}�e�I���!�Nf�6Yg������wH͖k�s9>,}�F��r7jȽ9H����]VY���R~ਫ਼_�ŝ>O��5������~��Rwo��Q��U/�R��Y�H4}��5YW��ZXG����_�}���=8����Ibmy��9�}�3	m��� 5��B�4��Ņ�D�
�OV�����빆'����6�8�5)"N\{�l;�#�W����C�`!A��z+�I���=	��Ӏ�<�/���<E�����zI@��(%�qW�G9�^��G�����$�)(*f��uv�P��z��ǀ��:��T�Q���,i�Š��X]a�Jh���T���~pZ��C�|��L~�^Zl���$�J<<|O�2�y���~@�i�<o�b�����.�� b���V����g	�)��R\��R��?L����b����қ����g̍�Qe�
���z��������Ӈ�5��������cW�'��,E��H���a��x��������ꙅ���>�Bt(� b+�>��|�~�Ɗ�8L�-��� 7�7�Ρ�i�� Y[��[�%��Σ}0;�`�<?  �[i��׼%����ܱP�V�����4YL{�*t�B�:o�����
����_ދ42�����&��E����"Ջ;f3�����(}�BӔ�/��L�H�F^�ƕt�AN�!�ƨ�`���,�lu<���El�XuZ�[4�o}�I*��!�?�{-��)�B���q�Mt���&_<}A��� L;#�;r�����dB��,t��!#�#��0��yxx>���NV,�C(���Q�`�"i��UO��Yƕ56�wF�f��LҨ�[Y�1?coB;1�\��,�[�y+`�}��qV+�4ASu�K�X�j,�}P7$�.��\�97�-.O���{�i�S&*��I�Q��̈́~65��`����NT뷛+��a������f����q�Av5����W��}�}Cvq�o��xg��-����;{z���bR��l���cR��Ú���d^3��J���$ZUѱC ,N��E�������b:�i����C%��m�<�Sp���٦(Og�l����5��V:d%Њ�0z+��9����� (�����Jc��9uXE�[Pa�i�(
)?��K��h*�D���g��q�\�6hT��J.u��F��7f\ʉo-5��짣����1�&z��B���5��Rꅝ�vV
G"MB�lo��ʮ��Xq�j�����z�,10�Ǎ�u��K�R�O���fy��2����t-����?�ƛ�6��i�O�B���+Y�ף���7ڠ�[�
�'w]��������W���������|�ÈE���*=O(zꃗ=�59�(M�̼o�A_�)1���Sl�t;s�(�:�Ąg{��nBH�YԖ�.�}���KN�Ly�>�!Eܘ����Fvca����7ak��(<�-�G����P�����UȎ��;{>�]?����Ԃ���� �����WZ��Q��%�
ܭ�k%ޝr�m�!�v���\�B�갳�����VH���6G���95&�÷�n}��U�=�?J3=hse���G_HCv��^ta�/�>da.�`<�]��[g�����<'����oY�b��&��c��q{�+/[��!���"�O�O�胄�	N����1�>m��^��7���OӢ�6*�eU��FC�|�٤d�0�@&(B@.ta��~��hn,��J�y6C�Eء%�A���~Z*�����./���H�a5��^U51�<��0(���L�: ���K�BV���٣����3�a�y�װ����e��3�
�?�k�o�twrY�w���.?Uf������-jHZ�xe���TNp��z�2^\:�F�'P�4V�=4Ō7'|�e��Źr�=�k�7��PX�~*���w�*��j:Ew"\<�\�j5u�a��Ԣ ��|��r?�8�yM�r�:A/����ϣ�ˆ9՛	�x�f���f+���4?�O�دE��=�U�aQh�\���yᐰ�=���]П�~1J{���5�����2L��M���*nB�� Xު�; ��'���϶;��n�g�}E"����${�%��q��m�<�r�j��A��ŝ=B��D�m�g�}�e��)��I<�ԆD�H�TE����i��gX����.��,��%\��[�y��#�>�x�#��?�L|�N�>�|�Q���Գ{��#��p�*RV	N3 ��V���3��&���^0T���>!k(Б_�����}��Zz76�,��l��#���7\��'yP���KH�p'H[��O�:vv��7;/�;��Ls:MNӮ��=����_���D�5bM(23৪�nʖk�ۢy���x �78I��G��=�^�O� ��5�>��?�����h~{��r�|q����գ�Ї�0Y���k���iX����;���/C[R,ʟ�������'w���o��b_n�*n�\)�d�UD����ԟ%��pulB2�"�o�m�BpHp[G�܆���I]TPs���+Q��/�C(�u�	�dp�<��Vkn����~�ߦ�>���tu��s|������n����9eXU��<C}Fy]����Mb�َ��p�psY�[J,1��YW������֣�wv�z��\�'|�ȋ�Z�ev�gbbV2OE�]�$Q�O����l�+0���׻��1V��eou������\z��"-�tj��j	�������׽�1лfiX���͟Zn���c��2��K�sZ�}'z��=�Ý_i%���c}��4�.+|�06�zf�j4��]����DE��Lw����5��?��>���Q��V?�c��]d|mis.����(�)�To�X���ɓ��s���`RIos�z��,;Hk�)[�0طZ�'�i�j`�=^���㩽I��^OlPr�B�����c��4��=u��;�U��G˂�Gc2��F
2tw�2{���̗8�n��͎;��<���2n�d���ړ~
i�-�S�O^k���5�0x:�3�H�
C�ގ�?_�M��3���:0U*9%Vڦ������^Ȱ��/1v�(Ϟ��|�
MuR��������epa�Ԭ,CS?&�I���kR�}�QO��tY����&Hq�G���� �'Bt��*p�{#���(S���*l=��X���%�ֽ�7��ӈA�;�H��O=�P�4^��,2��~]$Xu��:Q���L��&F�,���Y���I����C� �#����0u�Z���ަ��-W�g)������<6��ď����~��{z<:u��5���~��"��)E6�>դ� /�,R���־Ar�C���Q�<��gj��h�P����iA$�4��(�y�S��*�V������z�?g�-'͗��P�%���+;ru�P�x͊]	���\�E��� �O��K5��_�;k��iy4�b��s�_D�ّ�~6
eK��9�9I;->�-���L���z.q,�:5��I�@ ��b�7gS�˼���vȮ��j���?�|��!Ӵ��޿�Z�3���ݫ�~��[ج�6�
H>���5ND��z�f<����N%g�FT+y����5u9{��yI��p��rS+���,7�6��1����~q�H����,?#<������|�Y���z�R�p�LI�d�BP�������D_Z���P�n�z�qv������y~v�ӑ2�y�H+Ɲ��}�V���0��u��$�ux�d�:G�֐�Ɠ~���<LNUai!�l�`p#ƫ��� �Z���p0�y	���g͗���(_3<>���cW�zJ-�I���3���4���*a}��삧�����Q���-�PJ��l�X80w����x���y��VR�x](/�"��/#�>�݊I-�o�e:K�q�xYz��#Lv��/�Y|���.��a��̍�͎�
<�0s�{� �o=���>H� �z�Z��ӕN�x����
�5Zi#`�톷Y��߉r�jo"q|Sz�����?�q�g��,��a�u�_�,�_m�/Lߛ(�����ȳr~�쾫�j�x�׍��fc�E�
!v�y:t���> $ţC���'��8t��T���c��1�{xo��<o������:���
H�3H�.�,����,O�+�/	)Ӽ�)z�n�HGo}�b������.'��Z�p8T���˨0�me�FYnT��bi|8��C09����.�(�[��g_&?��Z����k��eU�~)���Pb��* ����.�C4������g�pB�2aĜ�����T2��޴]���*/4Bc���s��`��T�X�T%�����B8�q��$'����Z,�a+���r�(m�[Sl(-�28ǉ{�L�=Տ�����u�?�������v���t ��汛�M���3�j��wb�l�uhk�����MT]��������h� �ܠ��5�|}�o�p���r��I��K���vH�,CC)2�����J�V&���~����ڡ��K �
.�N@߈B��ĕ�K��7���e�A�"�T�r?�?�M�㮃3FR(.f�mΖ���m��N�55����W����^Y_eZg���yI�]���-���P�Y��:�o�|Y��Eg&e��|9��}.�-����Q���u�	q۪L�)e�q\y��/^�%<��U7'�����E���R�*)�����2�E��u}뺁��{o@Ʀ�.RAm \(���♗���PH�=�@���S�s�A>�i�l�vF��83@�R�ߦ�ʯq���p��y�M{�ަ����^u�hԁ�9te���'3��4J�.C���405��iu�I�g���"R{orL%���xrϚ�؀�Q��׵c��k�_���ř�ea^�}l�'�QW6~9�}�ء��}��`�T���H0`�%EO���hj��=T�m��-��\B�M���ĺ넄^-+ݳZc�|=��72`D�?R$=�8�w���oް�ӊ��^(�� ����A��������4�ƣKetn��[�fQ��)�X�,�UT0�t�po�n��f;A�D�7{ۃ���me�s~��b������^I:AC)��IH9	���`#A�ag|p�����K���2�4��t��u� �{�C��@���Ѐ�4�o��E^8Y�̸{7�Al��k<��ͺ����s�l��#��>L�=Cэ��c6"�&����qmȅ������4�u�����E��!�0]d9�J��#b��
��3k����0��^`����Ή7�
XƻLK��d����#��xN��y�T���~p���G3����SvN'D�=՘6Zr��u�h�1X�iz��7��=��H!�
dca�i�u��Bc;�qO|��B�ܼRl���8��iV�v��C����b
�s~���7�{�IW�H&����Ԁ����~:��䬿W����:l�֍)D�S3���1�-�?9�d�ne�`X		璘��P\y�R�,*)�w7|���W3�0/��Np���&�S����K�$���H/�.�<�-��!����ͱn5�e�|�"�y�����+����|>�?�t���.j�P^H9k����s�eH�O9.����#��DC*��m��ނZ�,3퍱��f|@('a(c-�?�j�L(=��i٪���1��}�d�t}��5��o2-.=��j+����,�,�+��(�w���6�DԮ���4cf,VP<���|����B_EU5m\����,w��vi"Q����ԫＢAe��5$e����=�b�O�u ���^l_W�Q�mG�K R
��A~�R(~B�뻎�C��
,@�ʄ�i��-��0��~����{
D(J�ж�������a��b#O$ͧ�_OU࣭d�=&�1׼�ʘ)������{{[���W*��怷��,�b;�į��W�e�l�[Ԗ(��e�)�^����;����dl�=��q�LM='���(�^��d�qC��gO_�i���}/�l�(pD�Q��r;b\����&-��2�>���{c��IX�'u+��Wj���MtbR�����Q(������=��}C�"����Ե5��
�4�S#Xxk�Gգ�e�b��\��b��OJ�R���dzGػ����g��=���k��z����Mua:T�*�u����|ã
� U��,��Nj���� �|l7������4�x��e����VW��t�3S���2���Kd������Osz�O�Y�Ji�Blr2�͆���S����� �>z(�?�LF��5[� ״z>vt[�O7��C,�`�,	[����1�픥�ȱE]� h�>�<�7VK�6h�R��.��k%�<��&�)�ʟ�R^�Bk?�?���zU&̽;�hS%�3^���>�>_-7�c�o����>� ��M���YJ�RS'P�\�C�Y��Rq�FY)[b©H�ݿu��d�sY���J��l�f��2io�GH_y����f�>9J����oY����*Ý�����W��o�=��t�.o�G�8L�A�<$�"�R�3D���%6<ѵ�/Z�v��i�-Z�y��u�l
���)>���U�u��'�>��ʒ�Q�.{��"���|�p�լm�&�����IRɘ��X_����?����mk;�P�Q�RE�T�J	ET@@J�齆�G@zG�@h��;E�54��!�� ������d����}�^{�g=��M����?)��[��rA������a���BY��C.��٥�z���n�9|�%}���]�<�������1��"	�e��Cvvd.��*��V�A�V�j
�۬�UX5�X��A�Z��J�t8�ao�c�ĭ�ٍ}��,.�+Ysߖ������Q��J��H�}rȳ�<<|ښ���H^ �����>0��{R�,��5�̟6�n�iJ�NCW���?��y�!E�K�ͤ�M��ew�m����ţ�k�A/wTW9I�n���ez���褎���Ko!�=[7٭ln
��(��̌འ	���vM�B�	)��dd�{�<�5�	�&�Y�%;ߝݯ��pI��x3vކ`��D;�\0D>G@�{:J���[����kq9�<���o�IG�q����$��v8p{������s��C���ř�e�1e}��c0B��#\��9�C��x���6��V�����ԑvݜf�f�:`�G��	ܨ�-V�8 �!-��:=8�,�iS��,f�͟C��|?T?�Qz�����W?��k|�]E�����}�y�C�r�tX?��zN����=�,4n�0h�$�Q6�m�
����-�dŹtt�$7}�����E�K4Y����²�Q�w��I9���?�����2��s!ڙ��2�����d���8F�� ���͐����"�(��f�,#��+)�o�3��r��A�=�$3�(�D
[��Ӹ&B��%c:|3�+�N�54Iı5�F��\�aDD>�5�.�m�Z1����׽h�?��^��P �!&<z0�#��k�d]һ�pl�=�V�i���Yi�ɸ��ﶚ��u��hLM��񖍑�_�5��(�O��q�ʬ3��/�kɆy��#��ڗ��+��sp�T�SX��b�%S���jF�֜gd��}~�%g1����O��~7����m�[!�8��]r���e���~��W
���$�wonҧ�$ҽ����m�YS$�X����n{���Z���[sΡ�G}����/�g�\Y��^��j"HX�a��2ν��@�"+��$�X��s�)d�O*`�����f]=A�Â���� /ҫ�d��_\��gGt)ș�;P"�(��~�>���tYxI����ki.����*k�_n�'�H��Bf�i��*���%l�����r[�1��m���I��_/tϯ�J���.}�s��ю})�G�ܽe�4�M�����Yo0��yi%_����uV�a1���%�R�ğd��W�s�_����׳���$ٴ��w}�����.��rf���aH�Q�$���yh+�Q꥿�t������J��� ���^�"�x��?��F��5���"�G�޸�yt;nG)�\�+S��8g�÷�f�z�M ֻA��q���3/�%E�[?o�7խJ��w'd	{�>�btz�dE|Ԙ����_^4�	���ݖ|%��C�����锫���ۙ������I��-P��%,L�� _E�Ωoz�8%�.;A���G^���I��8�O��Yr~���m����QV�R���\��P�m�#�a��XP ���.�0�N�-���U�������  ί�<
�=t�F��K2�4��ˁ�!�>!�6�*��(� �k�V�8�;���߆�7��J��~ћ*w*}ǊE��i�˼�Ţ�Z�t,�]m5��8��Z�yנ�-��1Dk>���t~��8}$�Z&&������ z/����("��G��=����q�6���f��tE.D�$��K�Х��j���I��������5��"��$Ʌ���J;�Q��<����c\ύ�5�+�#-�9qRFfC���?敕�n���y.rd�wo�z�IIAy�]V<�bL,{/:��&6�����6r���2�~C�E< !2#h���r$��"Zr	b�Ks^���(���ة�u~�nx��FI��O� ��oGG��$���vr_P'��1����-kQ�#�ǲ�u����w����Z�K�����o� Jϻ+�1�3*NNk�m%�oi��2nH�_l�bİ�o/�M��X+�Pߴ;��@2��z���T�~�����NZѣ��cV�ߕ�^'�I��/S,&�G�[@��\Rd���s`_(�s4�o��|�.�Dz:�z��@{=q��.~��pn�*@�E���t/�y#[y���1nN�l�.=Zػ��Ѣi $�:���^�����z�r�AC���Ĳ���H�~O�҅iJ�j�fT�S)㥴�RHW�v>6�brz�q*Y#;X�`���]��"�$�d)��1Y�O/����j��C�tKoIlq �?��G ��eD<�n�1�Q�-՞��f�9���$h��8	��(s^s�u�ۇ�����m07�T��I��-���eXPlo��R�~9���%J�^���4�B��4w<��&���ʥ��O���&0P*��[�N�R��$�bM��t�p�vq�L4>Q��W�h#$7b�%��)�?����G���(R-�a��4AdI0�O�j�i�"8�]��������X$8h^=��Cnl(��QE�P'x#<jL5M��W�n��4Nk+L㝔N�g�ǮȾ}^����t�D8�X���K�57Y��A�y"V�1n�o���B)j=��!S�g�5�S�f���B�(Q�U|6�9Y>��W��
�HΗ�i�M�N�ITGE�F@O?v2+��t~E�� j޻�c;,Q���}�P�Oh�$ev� G�Qؿ�صI�]|lt
�4��.PƷ�:4d=�=q�����"yT�ҫ��z�LT�� �w����	q���/������{�F�n{�nմ3�dij�J���3����Q,H�^jYʠU�+��x�(T@ܕn���:���4}d��h�r���i����M�ĬD:h��2����M_0yO�!N�h
�V �צSߏ0�_��sE8 -�=c�Ԥ!ą0!Lo��xi}�n���4�m��9�G��k~�O�G�w�r3-�ɥ6�wڨ	�z�yn��L�_�T����W��u���V�0�K��xN�6	�
�+������sHFm��3�D�O���}&�9�i������ߖ6	PyL^�@J���=��N#Q�oG�O'+���x�I�A<��LB[��������'��*�������9X%^i�ihR[B�[��9E5/�z$/m�,{����6�	��p�`e$�/(В�=��&����J�ҫ����`�m�FŹ;�M���i�5�C��,Ύ���p=�����I-���9� w�"���fg♡�K�͟%��K�Op(��H�v�bHd���A����u_ӽ��������J��נ�k��,���#��W��M��z�nh�reE�0b���j����	��I��|�g�B��i��P#�x�ō!�������� AaꃄG�dWW+�������u�[a.��b�R���������EXM�4_ƭ)���p�X��3i��� ��ul�<1| �aIA��� �����"�x�4��{�C4�採�,��鎪V
����+Ŭ�F��,���z��ו��<�1��5�&7u��ARLoN��dվ�
}���Y�Z��hm_��rk[��i�kF҄���K�S��:����R����3�u��J--�-����
fb61�C����î�^#!���e�������|C����=���I�H��H�6«ղ���Q:�+�Rs�����&]��5��j�T�"�޽e���LU�}�����M��d?D^3	zf�|��fAP5i�Rg���/$
��<]��M0�f�������s7���g|���^\��!��-���F�������w3y�?�$if�7N�����K�P ]�2��~����Ʌ_R�U7��~BJ2)���ړs7>�� ͘WKal���m� �����OV�&��[Q��U�����\�6�h��7W6��	K�D�>��9�)��u��o�
[JJ���~⎾��*��e�8��+^[kS@*�����v���e齷Y�f�O�l��':���Q�S('k��n�X�n������2�v��]�rE����P��7��c���[�-���њ��Y�������GҤm�^J� ���'��I���zڽ�٬��黚9j߇����u�t< jڞ��%��C�}�Lr�#�r��H{YG8 ��J��7<�O%�ݎL{�>d���`M�q�o�GQ��g�6��T�9�Z�#���uqK�����*.�\����YU�������Q����tI>�r4�2�U�@�� /�i��|�E����V�K^K���oiJ3�IGE�=�`T�w����C���7m	�a�U����R���(�0����zV>~3�c��Hy�-�Zϋ&�o�D��#�.�RmM=�&�pP����i�n4���U���`c����Fq��������ĠL常�T1�:WH���i=O�B4��vU��8d���G�y�4YӶ�����hA���q�[�F"��D<�d�D7rҼs�?F���*a|�#�W����B�4�G��N�ɤN�ۙ3���W
ӯ����EH��le��3����ma�l������尼�����p�jAM��T���V��?cي���,��j\��a9��R������bS���>/��L��2.|�=	*�f���~���\��g�WH�/!�O��z�C3�Mw5�_U�)�����k�qz�� �w�(�2:۟�!yK���:u'�DWQrШ�m a����p�Ɋ�à8)�!m�%�}MpYɚ5|�CBH�P��4;�'s�'~�&�����M1�Ywp=I�saM��;�LBY�O,�OJY&z5�fq;�=�Y8O'����}�#mfXծ2�6L�䙛�k���;ه���C�#���r�F�W�~�R�L*&��-cu����^�ENJ���+�Vf�01��GS���sK�ŀv�5ި��Jo�OB��gz�m@��sR�R�a�o�⮉���������V�,լ�$�6o���)�3Q�U]mL~|�����E�5�W�[B��P��/�=���#������}��T<� ��g�x9` �1z�{Z/w}-�{O�GC0�g�
A8cڀ����[��P}�ej�2�r8�zt6�oD@�(��Ю1���9�����*�Ć��t�⃐�Y�-�dq6��N�"V����>]�;�ژGp��m�?��w����њQ�y^��bu���t�&Z^!�i"pP��l��F��'�(��I�=�p���=YWn;O!x2ڿ�j�Ϡ%���\H�a+xhl� ��v�Hװ`v��yekG���X���	|G�� {gXW�[`ʪPKNU�����9���"m�&����iճR�ס^��2��6m��I�e��OU���.��ZԶ->�t�,]'y�.M<t�~���	��}ż4��{��2(�[{2��to���颹��Ύ	K�_��I�ԫ~�:J>z�u�i�R��QŎqmh@"��m���J}$��q}(~��e9�{��v�Q �h��c������t��e�Nܳ�����ͤ� 1	w9.e�:�w�J�������fu?����,����֗aG�Bl\�� V痰�sF)���<�>�{��6�Tj�im�s=���C�6��X��AaATgTj$���7*m� �ֲe��9K���Ӛ	"%�jwa�B�PV{���fe Mm���+cw,%׹UvQ����R_2:�ʢ��[�t�?Q7z.�?�h�;&%�p��qّ>蹊���� �d�����Ɛ(�ٝN���K�t`��ߵ)��7���S���w謁-�8��mT�k����Ծ,AJ���{�T>�r�='������ص%�2C�<)�ʢ��5�
���=�Ho���@��Ź^��M�B)ߤ�̯��#�U��㕜z:��K˴�^��c��iO;%���T��7����r+ӌ�#�)��SE�^]�çP~��l����	�J&V#���6�� ���*+X�����Ķ��2@��=gi�s|��0暜�4ĩ�H2����a�;p�c�`m<���Y�W*�L��p6`8|��!�Ɓ7k%-��fvC_�����8��O��/�E�z�����d��jR�F�����z�[P�O�7�<�\#�N�~=;��o���0f��,i��Ke�^� \�ymO�3~p�H9�+@��9���+�%���(�i<��g4�=#��D�ē����ޡ���)?��뗾d��U3���M��]���y7���v�����-���;���ڵI"��]�i��u g;�S�����IO�f��u�m���Y����Xݽ��4�c�����O|M&�b{�	㥗V6�|Ps+n�S�𵌽$O'�8�%=���/���$6��Δ\�f��p�7�u�z-��յ�r���Ǖ��y_޺�	,*�(��B�1�n���3��o����ǓuN�{6
��vu#�i�����7���?kU�D�9��>��m��B��"�q\�`�C����GD�`�*S����y]`�ɱ�V7S�{�
����wS_��� ��?�8}x}�
޸>�#��%,wD�v�q�w=��������'w��gO�����I	��W��3�jZzz�Un*�uj����D�����%'}2��\/�w�T��]|r�����
$�%W0�%�.1��3�$�u��1�[�A�k�����x|�k�]�;Eb����z�q�`���O���|\ʆJ��-|Ka��^#`�.j���X�Ĝ2Dd���KA������>0~T�t��ֹ����Fiߍ�30P��Q��v�`έ!���[��13�������
]����Ё�&E�������zH�/dQ�7e�����J�Iz�.�r�@����b�����<i�d;c҆�s�c�_��"��\kj,�BZ����%bz��ZL�����	��V�[`6j�b:0�=8�����NȆi'K�~#�
u�o��i�$�9�G�V��p�܏�Q!#_:��4���)6�*��:!����V���>3�mq����=ta���g��u.�z�全G<	�Wo��U峇��o��&�y�G?	I\l�U?=�����2��\�]�rY=��E�O����z�߂�h9x�}8R��r�]�?�����ㅦ'����j�iv�*�ݔx��1?���L��b.��E݈i@`X��`��5�ms���ȋ��}�I�j����$�M��w{�x�k-bl,`�Mk��	���>�t�&�1఍�y.��J9;?�#ǌi^?�(%I�	����r�Dp#�إ�G8�Y�#����4$%�i�L	��?�Tm���_��H�)��SE4J�*>
�*վ��W$g ���p��C%�+����;c��j�Ean���>��ډt�{g�����-'�0��@@���c$����ё�kz�U�|�R��d�>K�	��.F6��#�XK�g�|�	a�Pn3�(�!/G���lP�ee�Ϻ;5��x�Nx��neaU��~b��u���?�� i�m�~�}�(�v{�x�$iЕY����b�x�D��B�Q0*N/��PL@l��,���7�&��7N>���q��/ߍ��`;�nOd��}56�{e�k��(�/�X��~��u�|�*t��"�ƭv@$'"�~���e1�����/�| }k�kn���+�u�fH�<�R�o���Gt䜣E*�5GZ�_�2/ޛ�D9��2�6�o�0iU��������O�9���ȣW���VC\���բ��(U�4�\�<�o:�l�� W��V?���N0�l�O:����|���?�%��?���1�:ٍ~���%�?��*�Y/|�k�~Xc�x=�� ;T�/�G_Y�|�82Vj�Mg�ߵ���[���$g[u$�Y"��.��J��7tY��Vq��xE@5� *L-1;�O��T&Z�s��9b��;0I�cw��$J�|%%!xoF��;���͕��m�ϥk4����D�."����� Zw�8�~J��!$p�,�!�����\���#/�f�|��N�r�q�\���b$UE�8����o:!<blGI���M7,eX3<��I3��f���w�W�7c�����?%*Z�^�O�Qs�I����	��)�B)|��v/X�����^m͍ȝ܍�2û~Q��q*��Y�q�����O�&��x����}O-��eyq��-��=�}��U����]���t�	�WGл�r��c:Yǁp �����^hz��봜�pY�酜�mbA������Xo1߱��Z�t�������n�����:)}����&�鱿�o�M�t��MSjc�����<�H�_KM�<�B^�Gj.��l�����;����W߇G���:_�����*A�b�S�e>ʝ8����q�Xh2�	H>�ˢ�h{>���[c�q�,����0��5SPX��=��Xj$j�Xd=55ͥ�o�h{��į���Źu�B�F�W&v۬s�uq��:ĪK���\]����,��A	�J&��p���ϒ�8�D�~���̩|GWSf�:�z��>xtc<������*zי�})�)�+/wuYu��h��!�Ꮨ0KW�.H��	s=֍K��������pg4�LR�Y�s�;�~,��z�J%����@������I�
]���y�fE��"�^�hV�t&?���4���Q�bj(�(	
�xŗY~��3�s-�vC�׿km�h�W�s�Q�d�Ӑ��#mf����oU����'¹��V��S����	���1�K�+���O�6u�UWĨ�X�6�݋��ڠ�Ca�l����U,��Ge�G� ��A�ht�X+�[��l�F�V+�HÜ��Xׇ��S%�����������f�׾�x�+L�����s��iV�����{�֨tu�?�aU�!�z��*g�]�vvܢV'�?.v^��n��x�Ē������{9C�ֶ7�H]��Y�h�蓥�1�K��J6{���^Ks���Kt�ڋ�>��?4Td'R�/-��Uk�L2ZIBJ�M0 r��������Q�����3<)�/@�%�D�'K���p�\[;f.Ͼ��*�`;�Å��2G#$���[���	Ys<��"5;Z�Y��lh �ҥ���ѻ����nJ���ZK�����\��᠍(��	��FJ��������a�7M~y�6)�S���Έ@á�h���5t���qB6�6��hF�����\{�4�H7y�P�����>nq���h.1�'��1u%Hz&�P����Ņ+�3+׿����k�I����J�eܐ`�� z�k�F�	�����:���1��8|�-x|�y�Ĥ`\�����h־�g��{Ө�}�7��n�4��w���~�ez�a$�Ӳь[HOX��f��b4��g���ٷk�e��~��u<ϵ�' ���v�B	L������ ����j��,,,4"��sNb$��q��*���{S�wl��[d��&K��o��n�Ȟ�G E��h��䉝V�$^S|:*(��l�6H������i�N�6�[Q+�����;H6���]'�G�N&���=��"l�8&U|��z���S���٣P��q�TJU.|���Ǽ,ỽw�mCTY��[�ӿUB��pd�s�U-���x� o�<���T��?�B�b�5}�_҅�n3�\~NBޝb�0�ի�,#��k[��:{�͒~K�L�Q�Q�$�Z:��~�]{$H�����ǩQ���-լ����cgP��X�HHT�ݪA�讏|E�W�;b���l��E��"}>X؏~�*��l����Iʈ�I6m�r�����g�'�߯Mp�{���@��;�����l�|�K��I����7j�K�$�!�h�cP�.��bE�w���HAx�b'�H��A�eG�,��l�G��z�ӽ�iR�//��؎�~i^����1K*�	�xh�z�A�WJ2ph�C����q��yԖ�~e�F����0ҮxE��)��~x��*:Y��6\�����(��x��q���I��&�X���N��zym�
v�5�苛�zme����*::���f���������e�hn_9B��D�ڞ��n?�8|�{���Δ'1�:�wӏO6E��q	�����Y��~���/ꪯG�����`z��`\�'��
��<�1����^�XN]t��y�գ� �~�'~�\����"�U�qpp��cf���~A�|,(.��YX M����6$����T�/����}���/��=8�tij�iIV��'N�J,���3��	F��LF�V�$��ٟ�b�͒�U10��L��ȟE؍:�z��.�����ǬNe�I�8��A'���ܣ��)�Y.	cR�Ϩ]����s�u��5f�����EAښ����]iiyh�B�pۭ�R���Ѣ���z�ڕ	3����j'��.H��l/d��1^���o�t��p0�2����~�l����(�^d����U����<eY$�Q_��G�: �
'6��,�ٴ���rT� �!����Ά�Q6��_EՎ�KY�}�W�)�R��.��Z��E���#*��#O��B�o�u	Wx�>�ܫ�6��t��^����W@���E��{���Z�}��g"L^���C�b�)%�Kv	.���z��x3yM�>��ۣ���j�F3�0�����	����I\�-p�Ut�'nj����ib�K��@T"���h��Ee�m9l.kC�]$��ی 2��9�g4:�Fp~�GK� �Q���R���)�5�&� 1����9�C%.~5���b�l`����I#M3vY>#��nlgq;�j����	�@u	��. L�",ų��U������e���9�M�hp+�G�g��1��q�$(�h�;��%��G����m�|���c��~���[>Ѫ�O��4Ԟc�WIש;}"��N���fE*�|E~���~e�q�.��}Ҹ��ko���^aq�&מМl
�cYT�I�!)��a�q�f��	�п ��
�sg[Ib�g*-|����*haa���~����G��~)J��]pfv�����-�=ȑ�z��N�?siɭ0�`����d�⻸��T�je�����8G�����^2X������+�%�|�EGH!Μ_�Z @]~-�7�%�/~���Z{zvu?��¨w�� 'C��䶒־�f�����%��4���N������W� �+S ˿.\��_�knu�)1�+bfڞ�W989&�7(��g�NK��7����@d�)�[����\��M�҂s���O?%�֦+?-�]�R?��A�)�i[���=��'��kG��d�V�����ʱ����ۆ��K/����T�Xnj��"�d���C��m �|�.n�-��P1[���@���c����;�B`�g����3�DhAzzU!����R����q ��)��:�{/��F�'����F�@��� �0��:�{C��+c��y�l]&������joѲV#U��e��(%Y��`�s?�W�i��U>�{V�mtG��R�U�O� ല��KM���:�k�)s2qN��ZO��Eh�@�����.��D �kk20��p��}3���67#�u��s ���Cq�@%�U��l�Ω�����s�j���+�~�g�#?w0��jKI@#����e�A�&h�נ&)Ό�A�u��"�X��U���
K|���f55�MW��~�h���ǧ£t��A��Y����m����rS�pX�ǒV�&�h��9�
�5�����s�; ��'�r�=���o�����	���+~��ib*|�:''����E�b����{Z����j0�~����7�=�q&06��q�-��t��}���-�W�s���U׏�g%Z�?2(d�b��N�M4�"����1ʢ�-F[������转"yȓiG����B��my .:kZ�F������&OU�G��,�?��s�X���\Ậ� �݋TB����6о������L�1y�C��kdt�x��V��:}"���@ë���P���h�CKaČ����x�l�[�L�<�� ��o:I����%�CwRLt�$q��	���@Հ�nc�*�[���/%�"Ÿȿ���/�Y��髏E;�Q����+k�F��2X&���U8W�J�-�f�-_��BAc�B���k@�@]��X�e9֋;��c�r69¸�)��T���;g>M��'��:1�a��PcD��+b�w<�&[��7-���Z��%.��(D�A9��e@'��'�a�H0�bj���k`u�Jw�S�H��9޴6w���\W��֥���.'�F���E�8�)�;���b%����R��J􎗥|��6��mD^�p��ى>�Kq'����𹼆K�}r���6��l-]����'��)�|��2��R�j�.8W��nZ�Rŝ�l�]�Q����@�H�H���q*��Ҍ�I�{��rvӝ��kI�I�&��Z�	"�q%I3��w��=��:&��,|n��k9�^1���A³2��?�q��R��*G����1~"9��7��-���H���l�QSc�ت��4<>^�'ջ���ׯ��f�Ϭ�ߓ?�6��;O��@9�������$�y7��K?1Ir��b��]�aěk�7	F.v@�����Z#�3����ߞ2;_��ģ]�ۄ���6U\]0{��77��~̓(x:�����Vv�Z���2rX�Ì��4����F�>�G��Z�p<�5$�3srv/�5k��dʱ�c�\���c�]��;��֗����VII)�`�Rg��	q�����a1��ي�u���y��wQ^���뵪��L���7������BqA�o//�r��������9������|���p�{�tW�uE�%�!_�(Ta��<�>	&�OnBMF�^�u#�RP�ŕo:�6ꢘ��w�^r�?��^oLd�9C0Õ]&�w'�l��P�=�a����r�?>�.v��s�ݻOs=G��H�x�����?Z�]�8�-5��e�&��A*:�O�O����/�.{z~Z��5���S%�3�=ay�i
���T?=�L���J&�ˊ��Y��^�=�k���1�t�o�6�Aos%�%d�˒���?�ӞI%���E���Û7聰�%?t�e�0��g)�	Y�u�+[�R���ƣ�d#á����V\lX��D�=���<9Y��O���'[��m�'*k�KZι�^0�]ӆ\ĉ��4�Xi�&���s�B}���Uj	�V��j�6Y'�wJ4~�:��bq=�wE��C��/Չ�Ҽ��6h��lo)��7;�:���h<kM���~p����Pq���a��T謧Z�/OMW�I4��&�`������O�
�3{��|���װ�:V�������81U�>5Z�؂�-��f�������WBj%���ǩ�C�X&=�c�cqc�褗!���w��}������8k���o����.J�T&��`j�|o�O|��EC��m�C��<�S�)��A�<�`&�D�L�������|$^�����O7�Ã⣺�d	��mv���"��l�V+1��Q��4ӽ���Z[��z�a��/�m��[�LrT�9��R�`�=�	�~�IEy��<j����XQY�_Wg�d�����Cg!�������.�kFLR���$���&q0�c��̾���v{�u6%B�Gz"���'�w�Jv'0�Y1����k�9`i~@�����0H:Q������1f�KC\App�AB[?�T/\i���FP�/���UZn%����uo)���^�=���o��U�?g���� ڞv^���3��� t7c2Az����bR�O�j���͑��js��Bu�򨨳����hO�~cXR��\x����[�����ބQ}�p���OC��Y݊��/�bwQ���r��"dz��c^Q���u��+�*99��n��ߛt�)& l�<��k�W�D�:B�z��Y�vu��x�%2�{C���=�+;[�q���`�^\V��`���m�����R�h�sq(�4D�1��獍�/<jn�ma��ѩm�}~��?���Aϒ�iou���ʊ�߆n��Zhr�R�F5��t;��-.2��m��>Zq<<C�������0L�F��:ZZ_K�o��"�&�@�M釥��W���<�^ڴ�.޺#"�&�ĥ�j	ؐ[����~�"�_��H���a������aG����n��-��Ĕ�^^�e"�a��/��~�YzeC��L��7��Ό^�M
�Ο��$���ϔ�*P������A�̳/"k��ʳ��pp�<�D/�i��H��;c��������O�H��@eq��ϫ�)u��@��lV��w�����0�z���U�EX��7�`p�~Y�L���r/�z���\m+W�*��W�H���� ���	``Ik�LlmL㕢5�/��D�R,���s
:H��0�?�}��O�dw�KA�X4*at�*@���5�>(���Y�S�"yx��Nl�c˞�ZA��z��W�Z���U���h��όٽװ�^��-`��>���B�Ha��wtT%Q�g�6j�N���� �w�r�}��GE���K��
t���=�2�$o�xĈkX��8<�X��[���^�u:Z�{P] u:7mˇ�{4���"�B��������i�ҝ�Ajlвl'��+����߻�x�7���8��e}1G�����bO�)��k�(�}�;t
���`�3{f�go����BJ���ƤP'�J򔽴���5+&^?�s����Mnp@ܟN��U�������Gm�J�O���ۡ�7~,�`��h�ݹc��!����Y682��쥽�2��6�F'<y�X��"�%��[~(���h&�;x���H���.������L��U��b�3~���e�rj�S���s�@6����i��V߳�#���!��"Y��h?a*��?�hz���W����{�el�������;2Z� � ��;�[�
oT/�9�	�j6�ڬ�/Tڈ$��"@��?���7�)�6�K�@:������L�i-�;���>�q5���Gl �����rq9A(J�;z��*ˬ��f|��vT���m��'��X�16��§>�"�}Tٗ�[>�eԉ�=�Y�_zK��e��3p���;���k`G�L�y�@f�O���U����AA�~���ی��-�3ӡوS�/���v�VE����`��	�
%e�'���xى�UKg����>V>4�%؂��,yH9/�]n��(('�}P���{��̶�d3
��c�TfM��8�AA��*Х^V��E�¹䒄
�(ol#�g��CԵ�M���������l�כ����bԺ?;��X�V��/kO��t։ ��'�xcy#���s��3�-19��(�Yt���c� ��W')�&��	�Q�B��jC�V���ۣA��sA%�&�P%�t�6��Â'��:D��ĉ��M˽q����->��P�#:���1�e�[�C�94��_f%��WU���;�֗0_�Dkc�_��|2�����u�9psWx����;�Blj�r�fe*�~� �x��>�J��Ŋ�=��	�ˬd\���)�֬�*�Q!x"K��_Jְ�F��~�$��J-�}�U�:_gc ~H�`�` E��:����P�0#w�͞�M���0��V�|2�ҏ���РL�З7�w��>�1qq�bno^@��x�ѥ�9S��UB[m�Z<����	��Z�(O����Z �0]˝� 3wc�6uZ�]�&�J��x觽��l�V�u��F`�[T	�/��H.e�Mu��[#�Ӱ��|��}9�:�O��^����2KUW,��Zn�\=����,d*���V�0�4FH���h)�Q�ńE־�ș)��z�����8B�a���g��~��
�E����jD}d�L3z �P��ed3q�"V@ ��M�I�P|\�bH�dۢ�&sp���
�_��(>����+�A!]fa�Y$ߛ
���]o�����C�!Qy{,�T�#��v�S
��0m�KL��c���L�ٱ&�+)��>JʂL�w��
���:�N��{��_��+�{%.���5K�8���gPn��6�SMz��xM�bO��l���ή򍙈t�>�hb[��Z�N����6�L��֘Hvo����#���A�۵�K�'[�)��_k-�����y_+���UX��0x�pYGk.��j4�X(��3ګ�0�)2�t��d�
�>n?�x^}'��I��qe�m�o�df��U���V@�Z�ʼ�(�*�]�)Z��L���]Y�X��0��J���劉�����ixy��������@8����R�ʮ��]�x��Q;t��p��F3����jnU����E
�~��kL_�gxW�{yB����'��WW�L���H��¥[e���\�c7_l���L|놌_���`S�p%2`�+�QLR�R*����a������7U�M|C�Z�+	L��le�CJ��5tL��t�Ҟ�#�g��3;?yq�t�s$	7�u������&�.���s]F����%���*�tn�X�j���<�^����|�{�7��VHm�E*��|T	�����>�1�����r�o9�d�h��5wl��o}XQ��F��MS�ה@/G�ϊ�(*D!����w4��X m��CA�Tk��|�N�`���\����VѸ�~^��f���w�� ��w��H�,��w���h�=H���N@fAg
���hp�-̕"y�+��8Dr�.]�(t�Z-����[a'�����2Rod�̡UŌ��d�hVCs?���~�gV�w�G��n}�@J*�K�M�;�H�e8C�	��\T[�����uI?i��G�u�C���C2J��R��ǡdg�]F�ٛC�E��=r�^YgSdd;��l粝q�������<<>��~�_��z����޲�.w�ͱ.?�ߦ�׶�3T����J6J0�*M�9�}+��{�����/�W&;�5)�Ѓ�3�'�#���:��j��մ~�V��e� �zh����z	4�_yO�\)Vk��r:|ڮy)�m�g��;8i�R"Ч�� �o����E,�_���\�6}��\^V���bnBq�����ڱ���u%��X5�~��8B.�+f�q]1�D/���p1ۣ/7��p/�}nñ���J�v�X��3��:\�=b�L�?�Gl<W��v�Yk��n�O�^��.p��A D�U��?��<�l�j]톷hn�۩��A����Wl��׭7Q����0-�v�v�+�%p��Gc�i����?�v���� �J��1� &�#G 2�T#�Hܦ٫#���E��6݋��' ��Wa�����;�����u@��҃+��Ư�|�9Kǉ�>i��)�,�5�V�\�����`��b��}�7򮑻���
m�\�{2>Y�	Ǧ�e��?���y+#u��⳥��?&�*��ԪS�w<�����)DBL�.)�$��_�M�)�jШ\��y?����}A_�dD�^�	}AU�i9���]L��>Ф��3����?�	���RT�����r���$ɭ�1�t*ʩض�F@~��m[`��ע���i��c��?sn%L*x�}q��X��I��ծqd��I����cg�<�`�B����̪q	4�	�5��(����9������7�>���]���Y�c?S�U�u?BI�VU�N�_Y綎ĭV�z�6�cZ�HӤ���>���?K��D�`���D�n~�y��Ѥ��DR��%�5(\0!��ɘƥ\ȋY�e9&�&`Yo'DD�+��`Pg-):��TNi:i����Ҹ��ީ�1�);z�EF(��q�c�S2'����v�~���n*�^���<��a^Q�q�>��ܫ�K��F}<�1��{���s���!یWG�[c�Q�
�	�\zTKk���9;`�ACZ�Fq-<�ҕz�R�z�y�ag/}yd&����-�f)'�U�6w��3ß-��Ǔu�C���oz���'$�F�P�΍�aݲPk_O���@�� r?8Ֆ� �Eh�42��N�w��
��4���{��1�&i9�O[���0+ݺ92�x�p��E3��2/���eL	�� '�3��lzXC�{޼����b+R��^Z������2 6^2�
�˹���^]xp����i.Ñ�f�&(���Fc{��2�꘽��hÌ��G��@QM�*����B�<�a�q��R�`��nN�,
��������c�A�êS�e�e�+�@��S���f�c���H�nr�+T�<!Q���2��{��e��$4��F�3��Jy��G޲�h�7_��u���b�}X�
1��mE2�\?����`&���?ZN�H=�|;�3/��q�����rS}q��GW[T�?����� ��I�6�B�ō�!/VW�;#T����3���,z�b ���)���8�ڗ���sw���F��Sj�%�o��//�0 F���Y*g�H=,$u��E��g��������j�Xwu���rAS�f7R'i�3>@d��k[όҸ��������r���e�|��7~ߕ�����[��:0�x7w��ϊ��b��;�y砶���!K��i�bY���n�7�.F���"�#o"���ʆ�Ў��C�ޱ��SRi+ƸC��kW x84_I���ǘ����a����������%�4�jO�5��~��<5gC>:ec�zUI�&-G�и 5�sJU�<eɕ����j�;<�����g�[#ys8���������gu����0����꺣��ҷP���4^2�<�Dg�����y$��dCbRm0��h�������S����:�5q�ϒ��b%���C��w}%�7�v��_��	���g��y�k�/��RA�����"���)�0� ����d�b0E劷J��;�Pt�����#:�΂����)(p
���
���\P2�+_+�b�4��-���Uv]uUE��5a �]��a�n�ǋLi\q�d����ڵ�B�)5��_�Z���[�ҝ��lP�J���+�]XYxz����������c�e��ɪ��9L�ZM�l�q�!���wz�	�<��I�VT�h��9<^Rx:l�(������\鮁\J
{��r�z��\�n1�*�� ���_�"H�i0�*[I�3��Z�I-�Ix�Ys*���%��D@�:!j:��k�͵B"��(a��Ѥ��[��=`/�E��m�� ,�2���H�s�N/X�S�ܦ�x�2�kM�m�'�_^e.�q��uX$�s����������S���Fb� ���wu�M7�7>�Tv�?���i���Y��sp���s�K��O���q(F(i}�m,&���Yp��4v�s�
�7=EA���--��ZL���O$Pbw���I��S�:��~���Z��{�Y�6lT7����lF>a��7�~R��Ư�4KK�WV����5��Evd��U%����Em/����P�M�뾆� ��\��~�>ҕ������ܞ�87!�:-� uHqC�R�sד��ƺ�}��j�7�B\�{^p�êwgX;\�y/u�)�Ťu7[8�΂�@��/�~j%��j�t,���k8	p��Vwww/�)���V�����C[����tQ�:�����Qlh��̍���rr�:;&}���+�Z���N�v֝��O��KI��D�����}%��@|R��y�|���6�66+��6i^c���� (�Q�Jle�]���m948�g�	Z�YT�(�ԃ�+�w*�٣��+���n�&D9͋y����Lfj%��*����%��0ҌXިs��Թ���J���8�p�ɱ�徉�jpS����1���Hzaw7�CF[��uΈ�e��0��]�ė�2߿G��5�L.�1�48n	�c1YB�02	�V�.���0���z*`y�a�?[Ɨ���דB���t���AN�{������ �	,u�|@�Ic��v�v[���&f�=t� "s@����g�R�rω�"S2>��*��`_�g�Ғ6N��d�2ӛ�ܵ�ɾ������'����6�ɖ�OV7<� U�׻�d�OM#xI؞%�e�ɂ�
�����m]'cW���������oFRcۇ�������q ��Ր4:��<V�]��Mq����D\ĸq�oM ��פ 7�t"���]vzr�Y�ٍbsJ56����~u����v���t��ٲ�݊J�n��������T2��![+]]����.i��ӰQw`/ԍ��y�+����+\�J�s���u����#���M_����@G6�륮��b�'�0؆R���+��/ǩ��`���i���^�8��'b\ξ��^a���3�U� ��W��T�O��.y�����Jq�Kɂ�k�����f�j/��ܵsr�U4��p����g�
�G�U:A��ܒP���+4grj�t	$�U�D�Z~���;O��c�\\ɪ�tnj����Ozv�§���h3!=�a�~�-��X�g�p+���x�f��p��G蹕��=^���Cz�.�����G��§l`E�^���e)�����D�zD͔���2n��dkòx��hfG�?��/�9��1�cS_�>��PǹzN��5�ׁ��Tޢ�E�X���'�(Ү�PG� �T !��q������	�g=�j���&��1�Y�2��d7��L4��� 	?/�J�{��Q;P\&��/������&b�J�-�q���f�zz3�v|�OQT~d��Sy�����hg �X��cM�pt�4�a��� ��?$MI��T:���x��OV��5�Q�/��?F���q�8��������}v�4����A�:�䍱��ÞtFo~8c5#9�E�%�D�?E���wU.�0�$�6��MP���݋�iN��hJ|�CV������h����U�s�^��H��F�ݷZ��|��w�Y ]
�������Q�e-f�B�Qq5Wk��JkKG�~TY��wR�{<����TX�h�Q9�N�����0"%�5�ʪ�My������8=]r�5�S�|��]��Jf^��;2	�?�j���y��к;�x�"������-B��f��0e���lgNNL�*-{tܛ6�_�:��b��&ӱ)�t�1!�`�5+�Ǔ��%2R��K�v�������>u�K!Ca����K�b�WI��w�����ib����o���4�lS�qq���U�Ya��Wɹ�E��:���k�Mպ���'#cK��Ι�SS�f$�h��Y�G����Pc�ڞ$wT����`�9�W��K�%͔<�Mã2{%����!�3�FΟ��ח�̒�-+ns	��Ş���@�����I{"6YC�ΩU�A�O�jrf�rrzdOw��b�9q����#OJ 3,F�59ri���М���?�����'��`C=�9�<��� ���3� �_C�e�k�_#3�G>+)��ת�_LI\@�
E��kKx��Zyڹ��&���D�J�,ڑ���H1��	G��C?	��
ZZL�M�5�:���A�H��r�y
�ic5��FX�v���f�����*a���X�=�@9��s��u���q[�2��9��b���a���Z��5A���&���+\UT{t��Ԑ��T�ܕ�����q���,���ʎ<���c��#�ڤs���F�mw�O���/��G"Q�w�Kv\�
^o_~�۷^J[�+�ze6�u	�
R�?�F8��h��U �5-�lT�jvv��}C�ق�Wh�f�Ŗ;h8���D����L����ޒ뉂��,.6�`�I����x�/}g<�(a��q[?Y'��O����
�*Lw�e�ySL��6���{�kwE��2&�v/�7Xʁ�RU/1�;�-�e����\`����fve��B& 3<��c�N��f���g��������k��`�GM�N$k�?n�_�
�X0?��d�� ;=�ϧ,q�y�:��*�K_�y�QV6A"m*"�������N<\EWhF��!(u�Rv�#�T{dE	�Q�1'��|�>�z� 越:؛w�#�[2�����B'VK=�<�	�u�
����ܯ�|�k�v�ڄ��u;�b"�җ�����@w��f��Q����eee���IM�H�e������P��S��e9�j��g�^��|t�f��]�
>���9�E��w쮫a���W���2���?:-]�R�-��y�E5{ś�ǅ��7<��%Z3Nq����a'�	�*�
�I�UK}�eu���C8W�p���C�ݷ�Gd6k������|6���Y��g�%ZU@;���Ez�29�Hh�d���Ɩ���T��i���������G��kT�k��D"-�\}CV���j�wh*#0#�~nX.b� �m�^*ڊo=�^�kv�&���G?���@
�h�k$h�o�?�\��ɃL���M7�_��c������WI}���C���&&�ʗMM}U�0�L��B2TJ����9ܩ�cN5w�$�\�F V�;8�ᮼa�m�����M�r����G���v蝽3�t� ��+�o?΃��4����"��e8;exaQ��e;7�@Oz��$�wd|��K��.#�twk��;��|��::�~�?C�����;R��<]۫�bu|�3��3=�c��*?�hvwLFĭ
T��Q�а�����������#;褺�uD܉�Fo��٭l\���Ho>j�P�Q��o���類��`����N���v�c�����bg7��Er�M��L�i��7�9�¹Ju?���3����>��G�D�1��U����oG���hg�\B�n�Oԭx��Y���.{�!��̹k��/;�������G��E�m�Hd���E2���������>up�I�)}�8|�ʥON~�n�[�h2_�l�R�VFkP%��G2 01���?�8-�+��0�J�`��ѕu8��T���H���1Fa�o�������2@��M5���j9�5�HW�G��"�vn��~0�sv�עe��K_�[�� ��Yv�5��*̤���8Kdd�p�,=#L�q��BE3	ܳ����t�;/юM�Y�Q�O8�yy���.R�������e�T^[�?4���GUuOɗ�;����;vX��
訴hl��1l�7��ß��)V�C��R�i�7�v���&7z����s���2��y��xB�E���;����^KYډ�W<W��䮘ߕ0����M��`~����x=Q�$U��s�;⨖3zuW1SF� ����NMSC"ā�� 1�C�K ����O!Q ���A�H��6t<���o��4����+x.���O��>�����w��i�� £�m��JѾ����7�T�^%oiکH� �j�l�JIn����q.(�ԍ�[#������q@���ud�]�p���w*ë7����;�;�b�#S(�2��{p���{-Xv�f�[�-���a[��.�ҥ�ub{xH!���(hå�Emu�'���-���5�|@�9/M�0H�Z���L��wzT;=j?.b�0$+Ǖ��jњOkw�
}����!�H�n��(���n��5�>#q����m̯�5H���i�V(���=;�u|�4�n߹	ݤl�e���,b�cW�laZ�F ���R�2� SO��s��3_����@ ay�i�x"��xzz�ߨ�
O�-H^c���c�>�B�����J�G�w(\Kߖ���*�{�t3�:���Br%�dx8a`���mq3�x+ڜ�A�봮�xf�X,)��+���L��[UU��M�����y��{�,^����Jr��}rjO<�z�>!;z�L[[�.�~n_	��٢�ܴ�m�s�#p�*lu������ũ,^T|HV=f�֌|��cR��Ep_q�q1\�_�U���)E'���9����������Q���b-��ט���]����t_�����]2h��7���99��V��C��b����	�F'��:�|���[s��v}���w��
�x(P���%t�O�(e =zW�1݌j�2�d�.(�_,�6���56�۷�K�rk�$o��vK���_bR	�oT�W1�����U���Ȭ�BZ�u�P�avSp�
�9F�:��:��x�K�d �"a�"}LEҽ���pV㙊x)6S�k�p��K�JJ��1�U������#㛔,0>k����h��@0U�]��L=���k���D#6E�ȸ��;�59u���|�)^�!6�U?��B�E�i������=b�]��L����L��|�Z�[�����_zg(@���{=Z��a;O�*�`��q.y`����J2��9�L%8�*j����$C�b�o�ܢ>'��74���6A���u�*s�"��bv���C�j���K�If��R׷	�8r�����j�G�+�����"�?	���v_�2��*N��"�<�u��G���ok��R'��&�����N��������Z��ۢ"mm��'�����r��*����Ӌ�eN@_8�
����8�p7���Q�E����z<u�m��c|������*��\B�v������b��IZ���LFT�Pb}����z���?�� ���Zf��x\���_A���@���Z��%k݊2�ob(^,�`hO�58nK
>�c�@��ż��`կ��!���rU$K7�R��z��O��5rm��OE�Q���y�s��ϛi%URf%����ƕ��?�o��B�c턻��Z�O��K��g�gt�/�� x �\5�^�JK�?߯��%8c�D������yTK�����k�Jis�/�Ѧ|�T��Fx?�C$�����?�������T�Qg�(��u�������o��%O�c��	�(�;$�������)�v/�,	��/s��lṦ�v���Jaa��[)5c�ԉzˢ�2S�1�N/��6х���A;��X��o�(k�1�~�8��K������ԭa�?�g|րF���_�������+�!g���99=�	lt�
:4� GGzG���[��῁��I���^z:GQ5 qLzT_��4����q�V�>����M4�ƽ^S�̮�A�p�a��4Dj7n���{���_F����x��PQ}s�ݻx� u�_3�nk�*�m�g|�Zh�xA����M׍t�?9��O��.�͕�r�ZC��N[f���t���sХM�!YJOV�ܖ��*"#:l�����i�*�y@,.���1LQ�92���86� �3O�YQ�8Ε�%���R�#����/"�#Y/�4<���%W��w�짏_��:9:t� tI�-(
8|ۺ���{��b�P�i�;]�:�6�)w.�W:�K =�'�E:Ml���T��P��4�1Ǵ;���z���^~�
E��zܳT�������X�T��t))��Ñ����:�}?�[�U�:�K����qg�pB����~L��bBl1/9@
`�=
���C�:zc](ֹ���q�CQ�hK}�C"��wO?��'/��1U���>>p-����d���iSܾ	�=Ɍ�#L�{�bzZd�U����y��ŕO�'�P����c"NX����P3�[�0����a1՘�/�$���
��2O))i~V��Mo��6-���0�����F�-K?��<=k .��:�t�8s�U�h�?,5�n8��B��aU�%�Mv�뫗�ZZ��Su�6h�+L����/����u�2I������u����t"�wx���Eh��*�u������jn�G���Ŷ����/}@c2���N|��1t��������Q��٪!�wi�y��^:B�΢�r�A���}h]740*��*����o!������u@�Q��D��s�aKc3T�a�|�9��偁�����E�6�ǀ���vW�Us�Ne!mb���g���z��(�|���]qU�I��+������dC- � ����D4"����F����L`z��1������umA���XX���{���p��,r�n�~�9Q�^��W˲��cn?��z��O��nfH7��6��� |M�maQ娎��I�n�&��hfL4I��>�r��q���f��_��A�/. V-��D�zM��᱇~|N�ખ��^~�a�f�#7�B<�i��y)��򦈕�&D�C�ZZ)�j[ ��"�/�U��|�������ݲ���gE���9xj��O�b6w�s��')����9������E��d��|鄔���%���s�'Vk	>;�z�)�0�8i��O^��Mk���I ��T+k�
uw���0�6X��Cp����މY=<٪����cJ �f��xU��~�F))W��>�ы��s�v���V��pK�����m�A�rrچ{;�Q$Rv3���콖J�O�Ύ)h�0V�V$�vl"����L\�,��nUSK���h?��Y���pI	$,G�38��o[�������j���*�7*�L�_��:�@6��6[hՔ:��4V ^a���!U�[j2��Qǭ����=#����d'S[>2D%��-Q֧��'~;��0"z�W�DbTŊe�5��	R�l�DNn�v@!���)��,7+���*pȅ��]��S�����E��Џ��@��;��)J��(�aRP�����b=�ֻ톬�\ն.&PӀ��d��_/&�ج���q�!�pT�������P�`F��C������c@�
�N�7�z������V/=K��N�I�u����͹��h�������r��N�|f'�3�e�>L6km�O4߻5 V�u���Ϥ�w�Gud����Oj+�������ߕ�*$(��!��ٮ5	�C�z� �U��v�5? ^���yd:!�x<��c�@_���Y���97�J$�����On8�0|� `��L?�-(��rÁՍ"ΞpR�<
�B����V?�}�ъ��A����\A)\V;���aDl�%p�,�e��\ D4���H��!rff�����p��^Ydʄ��F�<��w�ܹ����s&�R9U��E�Y11�| Fr@V��R�#Sy+�^��J�6�V`�&�S=��D� S�-��;5�w$�Zd�;Cv�i�9��2�Dԁ�ZFI=.Z\�{�^�g4y��KZFZ����:�6��e��j��Q��W<��w��B;�J�8�������Wu}��,R|��K��?3?�xc;��ZWn?����\6f�JM�N��f����G����d��!Ƹ�|�5A羼7��᪂�V��L�\)u��^�E�:�vڤZ���=_���PN�h�o�_�)�o�Ç��/�T�㶑u׈��ۄ��o n;t�T9�����{�^�I�(USUU�����y�}?��6��m�nGJ�~����oN��'�U���v �5N��uk��Y|��i_����b=0�y�D�{쎌#s�K�kA<.aжv�g�N� ����UBs�5�5O�� ,��>�,�Oؓ�=���#(����FM�c��H�A�=zm�m��w�Dj~^��ܢ%�6g�|:�SW�)���Ç�?�3�\� �IY0_��goyʙ$:�C� �(��ŗ�,e!���۲@#6RX��?��/S��|�`�;�Ƅ#[��5�����k��f�P�Y��s!L�I|V��UZ������E:�!9FuW�]=��^:$��?�h_�ܼ��i�=|fF�^�J6�jNlkgp],�8�yL�����I{�`�j�%ބ�q0�٨;� "���.NFQ�� �~�"tc����Cᛲ�1S_��R�ƝS�����,�R+|��y�?�;�\����ۭg(����\jn��C�X��"��Q����K���`�K�-�÷6��������."�}h����υ�5� 9�`"�9���/�D���xܒ����+3��"�Z~�o:p;�~�(�ҕ^@�QS�*A��:*h`E�\������(��.X�L��_;����Т���ܩ���P��$��_khY4K���k��6	9S�e��R���?O�8�,�����H���L�+_��A���a�,}4������$c��ݬ<��·u�pdn�8t`��}2a}Z���zPv
��H0����֘����x����>I��R8j
~�_X�|��R���FdQE72o�0pģ�+�"�<�0t&IW״9��-�tC:���T޶�5A�Sؙb\񔣿-�S41��Nmek_��OmY��Y�x+��A̒I��*ؚ��뜞5�p2�?��T�-�����τ����,=�|��4ME'�^�{���X��VS�E]��7C_d���1H?&	��)W+�|�|lh���N�s�?�9n?3���+���Ã�J.�&"���ǀ$��ȱ��c�/�Cߞ�y�VRm�آ�f�ܟ6x��z�
J5������PËo������@��)u7#��}C�r��9w�?���S��ݽ�8��q�����yT�XLH������5������#>A���/|f����8�6{{N����o�DM8�����H/k�rL���8��Z)+C�����Ѧ&�j��/tj����S߿�Z���M�A���YSF׽��
��#i�ٜ�T�)�wG�4��+�?|=�?�{Ɵ��4C�i��o/�4��-4��0V7�:(��B� �lQ�kR���}��my�t� �E���UW��x�C��\Z�h����ߊl+<;�b��ů�M�%�?Zm�h�]^�q��YM�/��������a-��G�ώ*�@'�]Gto{#�AQWσ-�����ίͷ.9���� (Ψ�pr�����J�ާ�c���!�cl���??)���Q�=��-�Z:3�l�Z�1F7�O�`�T�_L��m��%�.�Qoiu% ����k�_N����ݑѰq�.���,��;a0.�w>/��@�C#w���^R��ԣ�OCq�b�����xg��%� +�@�:#��<�[�(ePyq���Qjֿ�;-M�:N�"P�������ќ�+��T���y��+R��3��:u/iQޟ"g�z�����w;|)K$x�Il����9C��O�-�HK=ه�Z���;V�""���j��������k{���#�%���2%:�{� )lex}�Z��Vq��c@�$�.�/�h�mhP94
=� $yՙY�h"_��s���[�V���<�z�+c� ��֩(w���}�����]�ٙuLG�Ni���~]���(�E�m~0�[�B�p�0E��!�FS�_��>�V 7!~�5b�����{O�A�bgg��+s�Ƞ�NI���
��n9\9AO�I4��TX�7~(^k
3�r����.�F�y��lӇb.��H�mE�U�z��~ooR���o��e����3e+�ދ�I��G�oT����\}^<��, ��~�A����@Q6'2��2���O��W�9$_�wά��/4"���`��8��l���(�b�m�ɪ���d7�)Ӫy�"(�x�"7�.�~�v��ݽ���:�I1H���ۆ*dM�����Pj>���F�vك9r*�����=+�����2���g��n�����JA*aruρ�GJ "lV$�YXD�ۻ�]\�$k/}�ﯥ��w���ɭӹ���(5�(>:8W#4��4�b�J��p�ݒ2�++�*WaVE��6=b�+�yc
}�r8�ub�f��n~廹�zNf�i�j$��Р���AU��&��IC��͂�{j��iM��u@���v+��Z�D�<�k,KoX>�+� � �h�1�hv��/��9�<�H#���`���y�('�Zn��S�?3�gi���gdtǐ������D%%�T5�*'�[�0��$����~�j�>E�ü�nF'�������س�wf���}�IM�]0���O���@U;�@�K��q�D�\���{����k��������ٝ@!��ڼ�F��_���U"SB�4[19��������l�����Ѹ�r(O����NN��}���ylv���ܲw�C�(�}ۛ0L26"J��q�F r���o�K��.5��=N��g-s������qh�߈���.�w҆����EUugמN�>ޟ��඘�vPP�����$��Ar^.�|ە��cX�FM"���'hUw����߇�e�`_�o��O[m�Ry�md_d>'���{I��I��ĺqVɱVQ������7]7�/�x}��ﭪ�!���ʙ6����ؠ����u���)�Y۴�i��$�?��	I��5� R��}dj'���Ĉ���Xo��_��z�b�[��j�ģ���D[GH�`���.�d��C�,�F7�mc�s��,p�L�-#\|�H�TO�7�sT�	��+�3��򩣲w4�� �6�	���"��~�h������C�ҙ�_-JeeK��6�>�@���2IU���2����{��G��m���k"��F�O[�"Rll���+nY�%�UB��fW�<̱zA�p���	���ߧ&��h�J�U���x�>5����mX�Q�Ao��W^�bZ#�fݳ�JZ/��m*ӏQ�%�l|
�B:�����]���s���OMM�ަ���^�gP���׬{��,�dE�~�,|�)}r��<��E[WՆT�^�t��o�A5�yp�`�)vf�^���r\�%n��8����[�k�-"���R���w#�6��9��*��n�I����N{::��v��RW"��ޥ~i]Jr�6fZ��c��ɧ*�����1�?\�$JaR�s�d�8*]�!�ԣ�
���.� �
QHH��u.=��r[Ve��X�<��V��������N;�C�Pk`Q݊J���J��Vrٌ|�'8x�>��5�mE��L�t����c�&�v���R�'R�� '�IN'/��Lh���r壗��b�8H�+�*e3v�(� ;�����*$�[a�\�@��:����Ӏ���J��?��R3w���`��TV����hƿ��9��>jY�Keh6�۰Aʪ6���i�&��[ϼ�G�l�'N%v_)��^H6��s'�ҟ�#!��֯�}�vR!d>���ދQ�ɧ�p���句����a+�?������?���5��ܼh'܍��������XT*�{�����&��R�$STaЀWFTA�af	P��"�N؛G��/߭?�� �t,~���im\g�ϟΒ؞̖�����R	���/�sE�j�q�]�9�Z/3I����
��~QMjj�c�����e���7Aj��N@ $�aXELYU�Ȣa=�d�	���/�c
p����i"�Ӯ^3g���fUCv(i��zf!��!x�y����hwhqG������xNi����8��
>��n��Ğ�*.�9ۡ��uS͘��+OPح��1T�5������wԞ�^~����w����l�O�����o�<Ғz�Z��n�ֳ)��ΌlW��D?c�-�������X30՝NDDJ�!W��9���Q��L���F&:�����ζn��A$�'�r��6e�~W�2���fߴ��� ��;JUT�1���t�,l �jqp�&.��3��qM9{�c0�9nȇ�F��G!�X���;�+"|����z%�(�I�P������O���i�ݞ_Q�H����t��2D4E_��v0l<���~���.���F1����4(�;�.�am�{�IY�2LR��]����ܕ�	@j? �C� �k����4���,5O�,�%�I�O�h�`9�`�tS�n��ouﾅLVp���姽�1/Q_�����*����َ�_��;/��k�u�]��= ��L�y
���m��v@���*�RTN�����jB����@�ԋ�W�դͳhiS�,l�����
�+��C,��0Z������J,�����e@�����|y2������u�U5D�(M��z=#���ck�ìp&�na�ɵ���@�n��f�eA�%ڻc�����n�Mj^��둘+�˒���F���R�~��-��N���X3��/C��MS�e�k)��J���4#��gB?v&Od���2�h�޵e3;8�=�po��Ta������/.��q����N����ߚ�X��7>��Lŏ���p}[�ǉs~�d��g9�¨�@Қ���:��ج��`��d-�W����oV�=��B俞{�5#hPmV��a��~��y���G�rb�������s��&p8|�,�c�"�Lϫ�8z#�Iɋ�ΐu8`1�[�tb$����r��~�
t�|ax��*�V���_�Y53K}���~%(��~`�w����.��_P[J���d��VĂug�qa1Mqw���."�r�7Q�2n�����p.�n=M͎��߱tư�+IU��qg����n��>�Vgb=j�֡v �?�i���YG+�]8��;�LδW�ח�>t�]bD���(h �]b :C)�1�4P_��r/'���tܞ�	�Zρf�d>^D5���q���Z����_����P�T�m��i���vn�=`��Q�c��v�pGc�"���*ۈ�9H������jS2��q�(���4�A�'+P[������F�S%Pͅ���.`�i8I@ʙ{��EVk;?C���J�lZ��X��<��d97sRO Uv��<t��O��	���BvW�w߾���8C�Na����H|�}��/5��>��f�4�ϫi�)��cWbM�cf!-��C]s��w'�yN��#�mJ%S�� :`�L�߈���f5�h`S>��Z6P���-���|�qT�{� ��ҏ�-�2�z�z�M�sf�O@{n��r���C�o=A�-��Q��`���l��\�>�s\�s�9/�%��8äG:o?��mC���[#�?�yp�&(H֊��mz�Dsj�[�#��MOj`#:�m^�l��K������Rd�0:U9�x��H�q%2��.' %=�g�̱��7'Z��uH���Oν�֦�N<<*~<��:9�`���S��n�\Z��1�s4
�슫� ��>�)���o����9����n���34��M�u�#��^#fc��H��6� ����L]�{����(���M���ΰdy4I?��v��Ee}��m��7g�w�c�ˋ�_�����V��b���>:6 ��T��Sf�93�,:#(��\���mdd+ȹZ���:�)O��ڙ�M��&4;�H����5���*L�A��#m��N��� �1��B��q�;��t'��J�w�����͵M�ϟ�$��[�z3)���Um�hzd�5��0� 2���If��7~x"�Dx�Fa}T��V��f�<��"qo��tVpK�p�fP�ao�x�!j�S��`�0���)͵�ī
w�兆7��tT�{l��-����Yr�և_3�'f��p\�W��:�-��b��C"�lP�3�CD�x� ZЧ�˽��⪫��m;v������fa�&W	Q�	���?�����7��<�Cb�	G}�%�v�@�t;�F�W��6���]_5µ�K!) P�8���YM.F�7�e�M�p賿���4᭞İH�N!�b��]qc�	�����J����5Z��AV�����&&iV�C�k�,F:"�i�)Cѳ�	��B�:(�]�T���6�]�}mz�����������~�����������e��l�p��&Wɦ���3�W�?�4�M���h���^�)�?Cs�^�%o��45����\B!�S4�s��&B��EfF͹s�#�Em�����R�ޟnx�gi��RAm�3xƨE:4�-|��־���mIV��Ѱ��tײ���ӥ����N����,g���Sb���cO>��.�۬C��KyГY7m:����jzyގr��
*E@D�.H/��t��Ez	E:!��� U���;�=(H�D:H'������������	[fgg�gvv��99`��)�d��1���u�ίG�9r��	 ��ɩز&e��������خ}���G�w�Tr1�(����%>����x!������.(�E�$r��l]�G>��w�^�0'[�nU��ĖV����E�J�-��P'� ��]g��1�c����L6ED4=���
��~�ݥg"�F� B6ڀss�'ǪX�������&
Joy�?o��Vb��������۠��i��k
�%�&i���k,:��Muƹ�#���=�.�Sں!���������$�fd�8e�1FKǁ��eU~׮
�d���Y7P�� ��1�ך�O��,(���R6��ߔ5/<M���&�I|����|,#z��s�����l�Tqi����Êa�Ac������gϿ��q��F�*���^�%�j�kx�򱠉���~���������^mx��k����d2�b�LC��Vіzoh�*���"GMQA�������B��YI<m !�弫e$�4���w!�� :���#��(m/�>UG�Sl���[:jnpA�]*����.���6_���z
�.���
�w�=ozZ��ы��9u|�Bz�?q�z���4��*��<��)�|fns.����������b�9s���L2�;�l� 5<E𪨬\��d${#A��`��Z^b�����u�lS�OA�F�*�-���z��KWF��w� {�����\ �J!H)�x}9��HE�.�����pT�*�c��3;w��CTd����1؟f()��Z��I�[j���mհ�z.T�o��Q~�&gVr�PQ�� x����F���
͜c�U�����]�Bs�����,A�t	ʶ6�P�;�Z�Ż<+ި[�T��_>�R�\[���2vI7�]�R5M�������8ɉ��r�f|�5����z���&�*9���B����_���3`D����4b��#���Y��dmwK���A�,�Ế:���O��-��d*��Xz�  /K
���?DՔS�W9�;맊Ô�:W���Eeʶ%r�wb:{C:���u��(1y��B�V��^��\�p��J�,[�h&�4y ���h��~�F��w�\�p� {��W���f����]�(a������v�<+ſyϾ)(*!����OKW,�~Wf�z�t^Չ���(��Uk������<ԟ���G�͹��`a�� �5\P��P4��OwS�T���|\��Xx�E.�:�=K�������y�c�1
Y�$c�ο9�Xq�_X�kn���ԣE�/�9؛��%�@-_��^�D+�lG�m�[�d��P��uF��&����
�H�r�DrG]/�f�﨤�`#�$�j����}�<���.�ֽ��p��58���=l11
����T]��,�
���prM~��m����d`y&>��O��^zwM"?�;�z*��"%gmG�ݘٯ�ו�v������RV�TZUY� �������� ���6X�iQ�a��E+�oY$4ߥ�ٽ�����t�wT	s���ʙ~���ZE_�v���¼�Mʨ<����:SY�3K��BSlnM�U��|l��ͺ�Iǀ.c	`�I��r�&f�.�R" [�.y\\���/�K���Vʥ8����I��I�}��=g9W
v��\g�i� J*����ܹC~�W�n��e��}9&���̀�)ǅ(�`/�˳�+�9����n����O�zn���k\h�8\�~9��w�+6����NA�r.dA������Y����o����Hv���-h�4�[ccG��Y|�1]�ZT��T���v?�o��3��mc�f�J�N�)2��r�9�<b@`�|#)1�$��.d�w���  1LKG��I�KA����W������ւ�S�ѫ��h���?���3�{	Ybì�ʞe(�8�o(�L*-H�~��?u|Ė,C�C�t���J��dL#t'CMץ�T;5�?�og�:���C��M�)k��m�|��	�1vťY4�⭔TQ�C�{�fc]�n����L�li��f���hh#�^K�X�0	Ȗ�gd��-6]F'W����j��F/)�r���'�p̮ ��c�oh?�pĲ��8F7���iI�䯫H�xh����jF ؅�u����)d���:����� ۹̔�D$o�۟�6�ŕlPo�Lۘ^��Ե�m=&����^��i%�u�z��g(Y����e�R%d��]<�g����o�*U$�#�xq��7(c����Ot�0���Sٲ��	"�C39I]�o]�ƹn��$����˞�y���DH�>ǹ���PZ)���\(�5��TN�a�q���i�#�͌��#�Bu���n:J�p�AN��#a�@{:a#��CP}+tnP-&����H���2UY�/���ِc��|y�X	�L6"��2�����B����BS}��\��s���8_�����\A�̼j���ȡ��'T��&[?����"�j���Qmz�6{r�ԁ�Y� W��J2�ǔ60PS�fc��Y�꿕���
.`�k�J��rf3H;�Z'2��/�����o2�|�3�������L��0�MҺ���^y���'����W�)RB������N�ͻ�:x�3������5����g�KyJ����o�M�W��=T�d��2�֓0Q�m��M��Ys�H���P�v�eL-�W�?���!�X1A`d(�$�G�-]���92\`��zYz�>�fe��-x��D^ԃys�mؿ�����*�^������f�����T���[[=^B��e�,늯i{x����IaNy�Ҽ���8Ed���2����M��(�%ɼǮ{(���$h[z���<����J��E�{%􉦤���S�r#�>���Qr��D��*�e+�T���L6�<�w���udw�x�oz�<Jc�U��9�����O��Fn�a_�,'|t�n�Ep6 �}�Lz�N�᱑Xt���p{�%�{��߶������P�&���H�w������(8�����a�0��h��f�`�N��@��`H���L�<&)%�� @�$|_L��o�L7��?�7�9�X�߮�f�Z�z��|9$���?�FqOФ<���!1���
�,S,c~el��n}�Z�HP&�s~ Q�K��#���@��3� '�XrcJ�~TT���^�N��;�mB�J��Y��\L0a��LW4����8��B�K)4��[eH���ʽ1_j����w��Mn�{S%�WOʛ��S�S�����W��쭪��0ۮ�id-�M^rۦ��x�GMs��mݢ�j�׼��If�0if�����KU
����k1��SC���U��z+�-	$��h�mG=��F�l��͑Sʵ�>�q���U@�&^f���?�m��u����r�����Y:ۥ�c����3ߘ!�d��퇦�`�X�j�d�	t$:���7��7&������8����4�Y��=m�P�v�\�;~x����#�Hx.x+�UiG�:Of��p���gL�״���D 
��<&g0�a/]c�O�_@ d�ڜ���7D���[K6�I!���3��Ec��;��nH'�,o֎}2	|9 cα��	�����+Y�]��Y�2u��\'U24s�H�����hU��{����y�v��X��mL�4��lfy�m�&�}n����jO-�B�a�][ t�l_PL��W�L�E���WYh��U���*����z��<�3{s���m߉�f��xJ�0T��e��86.m5����@"��DGh���$���@l��{�0?�:��Qn�Ur�'�e"�=a�il(�j����m�y��{�?zBk`�%�fd�fc�:I���t�#N�;�:Jut�y���9%4S���j�����i����a�*�eՊ"�_�9���З
�$t�H�Ϭ�����(��Lf`	��NU#��t'�����F�*�25��~��0
	I� �+��'�����4>M�C]�8���<�����x��,�*�($��a\����Uz�е�� 6�ֽL(���哊�����U��o��*��L]��b�)N ������E��}[�T>N���j���޽�H(-�է*����,�3���v�[:�:�}������.�04Ҳ_���F�#���!YJ��=�x�L�c�q���x�3B-�\���se:�n��w��\�E4R�/c���o>j��/��4��e�E�܍��/���u�z��s9`�=.�-�kVSL_R^��Q:����lj�WԆ�U��o:AV��/7i��2�ʘЪ�/|CVjůs�b���f�%��EVR�6.%ӧK���` ���2m(֙r�m>O�"��.���O�mh�^Zh���,��g��ܩΰ=f�'�v�sO:C����2?���Ͳ���a-q�Y~w��;�ȁo?_�݄����8Z�-"����eT?0ٯ5��W�aw.��W��sK�WHa�.Z���ާ��_k���l��f��`��";;�@�W^���>b��~xl��/��o���ͭ�e��.q�O���sMH�9��z���ø��4b8T�O`D�ϩ���b�߅�dn��4��\n�ڧ?I�_�f��Z#����&�4\�(���I�B�%�q�n����l�/�;�$h4A�y��K�(��O���/��G�>�Z{��7�g.�`]���$a9㕡p����,������[X��x1�*��%K�SRg&�3H�M�u�a�ʔ��z�[2��vM�T�g߷�z�@@�{�ȀC�=�gx.�����SXV�V����ٷ?�z/�F�Q�}"�X(�p}]:ps
2Z��t�����$�h��<Ɍ �8�aQ;VB�����n�'�O�����s�}F �'m)�&�E&u$���up�6V�V0��̂����L*����O�H<Oh+ltN;��v��	��r����& 99$�{��b.�{ �|����#]��$>���p�)�?�(����}ߐ�n.fv��i��x�a0���/�.�?�`�[!nԕ'd��}o������w7�N���5j ���pmـs �Pjş1P�$,e���t˛{�5h��/�̹.�nݤK�E0:��]@� ��8ϭ{$t���R���F���#P���YM�ȣ4G��g�eH��=������V������֫��=�.[�܂�N Y�X�p0�Ȣ�ŝ}702��h��T[�95q���H}��[���>�&��_�����q=�C�óp�qɗ�r4�
��!���4���~.�W�[�)R��U[�L^�/����6���a��
�ݾb�A,v�*^*nd��#l��H��S�}͔��Lz}ݤS��_�:#Y�s����#i�rJ,v�Jȯ�j��.6�b�	�	Ѯ���ˑ��!��O(8����J#���RP������aՃ�cqu��M9{a�n7%�pZ���	!qӴhO+�4��x$<��}5�{��/73�R8�h{x_NX�5�������&g�"`��eB��1c[������O ��6X[	�.�9}Cur/:��n�ǒV�5+���"&��3��FQ���UoL�Ps���#ϼ4�$ڕ�Mb�f�l�a	1>C{[��^�۸���~�0����4b%�U��u��J����Z�$r�s^���x���r�oU��ߌK4G~���%�choO��1/���1��y(�Mp��6�ޏ��#�ۻ��
譲��ee���w>>������a��u����怢G2}=�HC��}9�,�*�;n����<�`�G��Ė��j�8��ӥR�¦��&Hݖ�y�G���t���a&^oY���c���0�X::^�/��;������p�)���v�#�1`Dڌ����I�a�2:��Cɾ�CQ7�9GSf��}�4�a��!�����g����Y��1�[�+f�����72�i��;�<��|�\%5�R�/&b$ac�3��J���=�vyEwi��ђ!�Try60=č!3ޙ�R�(�c�=9H_���V1v �X��ى�ڏs���z?+hL7re]�rݧ^I:g��Q��>�m0P���Z������;&;ͷ���2�O��(�g�0
��[�X����`���
��˭�0���	;2�E^�{��m*��v�b%i�%�H��0P��oP�=��Uv/�Zl]�)����S Z��$��|�u��=�%�v�j�J����e�m?%x~���Zn`�|�n��q�ʸ�>�����b���^�U��PG��X�����o���=%���g��!�I��0����Y�ق��)��pٶ*N�;�
�� ��O8$�	�t_�R�!�9��pA���S����Sz�O�Ռ�v�藉�򷅏�S���2��0j"�ơƵ 5Y���]�a����A[[�d���k}���S{���0�VI6�5�����$�ڡJ�1�X1s�ή�9��8�������٩7��|�'��|y��E���ۖYg�t��f����c���U��#�72^�����3[� �2�����%��\�R�i���v�Ok�����U��*0~�E*�|�xf9�Wq+fP�n�5'�#t$P>������0%w�j����E�IWٳUTn����+)ǂ�u�ڲ3�0U�t�d?����-��t!�ȡ�������߷��V�eh~���y�*m^�KD;�����s�!w�]���w7#}�� ������x{[W���Ͱx����;<�σ��]�y�����������ʑAŉ�}'���\R���������׉J<���*��qH�~��`z�������g9{�Z9���%<�ʈ�U&~��7g/ۦ��}�'��#���ac>Ȭ+H�V�O:j�$fa����1�:��"��_�����'��)�U��[�h����H����AH�^��!�KZ:��j��P�/�&el�I�N���[*��E��>&�-�Ǐ�&z;��ڕR�ُ�^y,#y��[�}zvL�¼�yV�NG���L ���k`�V�B��FZ��	���b���`��|�6i�F\ʕ�vd�����?c�,�MW����UD|�R�zs�Y4�찶#f�1��@�]�%H�!�E���F�Ww&k���	kl���2�|캢�Ĥ�Y�(�������+{�{����~	B��
zíiM��g��gⵏ�������M�,j}��T��O��:Mcˇ��Ѩa��}=f�����Ҩ#�����q�A -���Y*�wm�r����0�#|V�a�1�������Ѱ��z�3�_W�Mv~�|g�=n��z׆X������;g�@��i�	����\]����)�י��R����w����xd���a~3��ui���:����5�#@�oB�����X�-E��f`�:D\�"�L�.�R����s�,���U�^�"���z+Ō�ҿnN?������/�0�M��ݐ�)p�:�1��cw |�]G�`�T+"����Έ�W۲���Mm~�n'>׬].ϕ�/��]뵧�*�svE��2"-�f`��7��=eʂ������)�O��.Ҿ:ė	�P�Q���������X6���L�YB��+�n�?{��K�ڭ�s �M�����~�\+�d����0~Ѫ)�� ��?�r�\���{�4=��N�x4���F@mw�X��$ڶV��d����8��A�ځe�t���x�ӂ����#�;I)�L\�N�6|�B�^2�E�/��	>�l�E��4�Fb�L�p�)|�Ȧ�x�jf�m�6w�+�\u��#!��U�Iiq�"%�9�S-}��z�?���]��w��0R��ׅ�WI�	�zb9噏d�9���%�EN�e�B����=\?y@ �V^�-�1]��<��
�Ue�tY�x��_�;���.�#D������4��9,�9���Ve@�|HN�3�[场!{�ũ��&��%zM���m�0����['�c-=�(�5Q8��_�Pva�wϾB�&���^��ʣ�x�; ��� !j�Ah��~�m�S	G�9
�o��o0��YZ���1�����O!L�!��>Tq��H/Ĩ/����������j��N����~���/�m�
�����%o��!jj`��F(O^˯,h��R��+M�ʄ�[��=�p�#���qI�@���P�sh���x�dO�Qmz`v��>�u�[IIܱ��;��/����	*�*�m ��D�E�ڋ��|�_�n&��S?m1�S�?�8�!��Uf�����L�	n݅<.{+�#��m���C3�����*��(�zQ����LAZ|�<��ſ"Ǵ7`�k����A��;#�|>�DxAB�Q#^	���o�� 6��tI+���RF�;�u�}c���c���T�In��c�3��kG���$7������.'<Е�"~9�_����d�oY��=^y}i#��|��S��h����
��ݏ;�$ĸƺ��=8��:�lٝ[��m��b��3ԧAg����R�㕼iw3�6�t�3�ص7a�Į�����̦�!=e9i�j�����Ih8����5a���M�fW�7��?0U2�ȇg��v��;[�G���<@ ���/��S0�<{VTn ��"�]1����	��bƯn�/�P�J�S�Ն�Gh&xC�H"��$�UAi~�j����	�2�ڞc�~��+�'���]I~ݱX�YE��a���]д�">r6y��I9�16��Ӈ��C���ﵮ��U!ya_�z��,�%��|�Aʂ�v�T���r�Q(�^u��X�����u�R����{_����x&������3�;�ј�������� �YF<�i�s����������u���&K��;w��Oy��M#���(���p簐��z�!�l_�P�Z����#��=��������w�~�=���Lr�9��wkr�mϱ�:��g�,�5v�kPͬ�}zx��ɩ�P��x  ҡ>6N;ж(gf��H�W���J���0�!�ow`�E���{Kxε�rz�kk5���\7]�{T��n<� ���eD�Wu�X���`�
����"��M��69����g� ��s仳&�RT;u���1^�]7Js������iN�ijڥz\�mi\���s�Mh��[7�x��y�!G4+k �g�>&z���i�����e%NJ�$�Խ�ci�ԝ�<5݇'1����l�0$���K]�p�L��U�����ߣ\\z�2�QS�->�LCؗ-?e*yȹ��@��QBE��w+Q�Ŏ3#�2��Y⣘tW�yU3�&�ȹu
D��w��d�Ha���&����4t�}^%y��P���� �N�׃5���ť��]�2�5�)�d���� -������L�>[X��b����N��:�
�]z]��4�����p��Ywy�ݍ�f����:��A%k�2��Y���0-����@6�]�x�ϩr�f?_A���a��2�l�t@ N�눎-t�Qr52�o��s�.c#B�|\�	��7ih��1⩽ �	Ϻn}�����qWl��˶���ļ�~����U6
�����<aL��K�ͮR���O2>�(��B�k�۟�YkT�G���,�X���;6��?���G��0j�hi�M.�b�-���oW��]�⠿���Cv._Y+�.8�5	�V[��R1v�l5�P��	u�{�ˉ�_QY�Cv��#I�Inu���R���o,SjI����㺧lC�0FME��%UV��֮Le<�e������Y'���d�i���w�	�]Hkg;�d��L���
C�M-9U.�
�q�d�:�_�c%�N��]))��־������,w95�ՓP;�e#����M�0@���6~�Ձ�i�0C���+�.�~����+͑�U��.+Xd�b��,"��$��y)�.GT������Xu� 3���(���S�/Go�h�Ŗ�o���/HN�������t��-����t:.��J�4{م��퉻aG�V��"���fvN��>�M輖rr���!a����6p����u�6�N�w`!p��#>��wo���2����?t4�-V�ru��ߛڎ�@M_��L0�8� jo�W-�},H��'�N���R�v�VM��r4%����4�}�H��
8��.�eBBUXw����o�g�YpU�49-1�4T~�Tˌ-�����i��*�z��p���נ#:-��@�'.�a]�K�눮�]E�T��}��24������u'�}�m�w�>��<;E�۩.^��-����2�^���AX��SS�$-��1��oc݌m�kl0���u+K��0�-����qGU�*=���=��+<-ߺ��4&��û�������W�
�c�
I�|l'����, �vͺ��i��cM��[���$9���_���^�,9Zk�Y��rsQ�u?q�^�ϛ��{'5�5ȱ�iI?��n�~X��`A׋�r��=d>v�����-��n�Wy�9�e�E�N��Sx9��ס ���CW��1�O�v2��{��}�N#�*�x �W�+�7�N��n=�Q6Y�	�%�-��b:ص|�^;l�EH��W�|�JҢ��Y���%����d�Lޔ p��b��Ӳ�O	�l��K.m���F�)3L����V����͈�;���u-��1d����Z��%��(ǧ�V�[��$2O�˒�F-~%:�^�ul���9𑷎@�2���~^(P�U���]S$ ���i�D�R���6{�"��8'�qx/�Ώ"�x(�9�,��K�/+�N�=�>�|��Xt���3�r���_�0l�y�Zg�5��G�z7.骺r�W���XiV�d��41�:��N����|���x��B5O��LO����6�SA.�}�u�@O7���5;ո�tm�-�s���?��/R�����s���Ɵ�8����F��?Է���R��<{I���<��[�̺A��8(S�b$����Ѣ'�`Ց��"���J6�cp@����}�@ֱK&��ۡ`BXk���U��g��~���6��{WC�^K�z,x����[���S;�_1
�>L����\��ŵ���a#��d����;PN�C�t���`�����?A=
����[ӌքӠ��i˛llnS��m��>�o]~W����Rו/&�����Bt�g#	�.�X��X	��*�Դ��*M-�+UE�n�:���2Rƀ��K1$5cJ����l���m���ߟ�֤e��vv?�3� �X��@�ؤ�흗֢���P��[�B�PՂ������ kM>�m�.�S��a�����SQ�}�p�1��sۏ��\a�r��_VcM�������Ԓ=d�ܡX7����@��M��q���� ��N���2۫�"֌�W�أ��v�Q��]<֣�E������Ҳ&N�)T��,�"e�h�Y�=��M���3��
9�����tK}ar��]q|�8���ff��1Tl�{��UU���Ř�T��#_�S<����0O��Ͽ�����zL��{ON-�<�F�D�r����+�)�pu�.���q�AW�	C�^���]�!)�����e���If�<K3���<\$���K��*W�٬�3��8��8�K��P���m�2��.�8�����۽�ox�N���l�9� r�}�~���cL/qtf�Ϩ��(j�K�$�)W�II��,W�kj����AW4��+�Qh@�o�kR{���T���uǍ]U�c_��c�[M<8n���4�]�ښ�/���DNO��eco}D�x��%md���ٷ�b5Z��-���sL����c��fh�ڧ��,�=)W�,���~�&�aQ�75Ot_��o975Fw�@L��e�j���g�U�!�QO�k$�F¦ΈJf��&	�ӡE���@�S��^V%}�iQ]�ː���F�;��G��C����Ko
�I@�o�nl��q�k��/֯��[R�"��	��051=	�`���'��/p���]�����gV�|�bY��5睾]F�}UW�R�.��D��R�
-�tg���l�q�g�.@OL`oB_�6x��c��>���� P���;���k�TAo�į�>U��!�'��x5����@���?r�}&6M�kk��C�h��mW��l�?�.��%EY�T��!y�x��漘�|+2���Z�|"�œ��J�< ��w���<}����ՓL}ƹ���P�?�������*&D�Fa��4��׫���ɧA|�$�&��b��p�O�	�jЕ(Ǳ�9)*b(Uz��|�P)�U�c}��<�pt����կ{����~�"�¯y��=
����Lme�r��Ǖ��Ё����Yh/m�&,�UGN�����`VYx�누~1b�z]�&�kc�*����)ۦZ%X��߿�%�	����?�[ܟd�����`�|�+�;���4Z�$�u������$�6l� �B���39��J�B!���9`.*>EM����L��@)k$��*�բ2�n�Ƴ�an�(�2Tz�C7倫�<������7�gh�W���-����?q/7U.�o��43&�Y[n�	
z*�����^oK��sQ$�h�V��N��yV#�v\��k}�2ď"��.� -GF�p�6�����|ܞ�h�ڀ����'xыy��=���ǣR�����0f�^��bE���3τ_w���[5Yp��l0�v�>�	�V��p%e	3�7GEwϏqN�8<�+�y�<(���0ߌT�3����F��gC6�v�?�ڙ"�CW�+\� gL\��ɤ������Tk��e>�}
4#S�~8-�+k���*�nyU� ��0)�-��2}\@)u1E�y���l��G��N��R�-�0��Q&��`����q���܎d�% r��gı�'�.4�X��ʟ[����Bi��r�b�w�3��1y,�!	p�Unw��+��^��3�@�5o�<[)���i��+�2��U;�6"��,���
�i�:��x�[�Dw����( ���A�U�h�>Q�#;� �S�y֚�����	�X�V�z�r�'яlν�7FWyلS�둖wC�<�=/�S�;�yו��a0�RN�Y�׵[�aI�|�nd���R ��~$?\��̖lk��b��QJh��FQCn�B�1֯�� t���5���+���������Yg�K�<Tp�����^�9��e(8=Rء���[X-��,�O�t&�3�g�<�/���j��|��s�v8�h����A��	��|���u��Iw�T� 
��ߋ&����[�\:�����h����2Y�l3�^��uS���(>��H��犥���������擷u�������B��J���-�"�Hk��!oc����nu=\b	�7^��6t)���TV��C��[4����|.��hd=�l�AO�`��>����1���{�~�m�
+[��ɱ���oC�j7��t� 4�c�<,�2�����^FqByO3��)�h�\cC�lɣ�J�xk�nd�x�BO�}p��V�K��w|��	0�/s�i���驅�\c�u���wf��hJ�ȓ+�g�hgy�^�bP��a^a;9�I}<��ly�sS�s rp{詺Œq>�iVE��/ �O!9z��',I����G>S��m�п�P��ҭ��c�]T�$���k'e��٠n�Y:�ٹX���}^�������8�<���]2�7����Rl*-���B��!��mD�"S┘�{ ��f�2�t#dj�gr���zR�F�Kǆ6n�ٷ=_[d���.>�+bG���X�Ш�;�(}<��4��h��h�:j�5��J@�\�����pSdV�����m˜F�9� ��=�Q�N<ϗ�	;�t�K�R���fI�E��A��J���Yy�C�;Kz��I͙ F#��mEo�v"�TR�0l��mlA��E�)�1Va_�|Km/���+hC�Oj)_�F+��� ny(Z�$��F4Y�'�{ms8C8C
]�VI6���R�R���:A
�$�5�llՒ�'V)��W�(@��<Wr$2*6���OL�>t������Sb��h��t�*ͼK㉠~��GP���(��֝�d���S4V�򥓵NF�1�0�*}/����q4��ZW
�:z�I\@N�;�H0����3�:��-?��g����S��N¸�/wd^�0;޹y���W�Y���<���g缼�5�&WЩ<�}����ޗ/�Q�|@A���C{G�xLw���L|k��_��l����s�g����S|$P����|�E�N������5�=��L����E��sĆR�K@�?1y���[
�>V=W����νĻ��������D��������j���r��t���I1�{}uoN��kOH�]:Y�ct$��T��o�@���B�,�c2~&6��┩��b�+D�,֍�>�D'����XA��o�^a��fk0,��z�;KA�cE���u���~���x��Fq�*��P���Ơ���x�s4S__�O�[m�?�Ĝ�­�����G��^�[��tgl�[[�[c��j�MK?-[R]�ʣ��~o0�������K���15nV\lMK-�tl�@�b��:��7hy8#BO�l���g�(�33~��O��Qz�B���K��'cg����f��b迟J7D=����,1�9TX�0ձ܌����ԬZxm�����Р?�j
��brN��ko�VZ������m������߃"/co��E�����w��� �^�#+%�{�T4�h�<�[W)��[����Q�Jܧ2�_>�;e����p�=U?i|�ǁ�:(����Vu�?RU�j�sv����/��_{<"�~��J����%���q}�������-t|çc'WBRwJܺb_q�P�#s��<Q%�D��T-�l�t�q�����l�r*��vj�������SSh�]ש]Z����d��V6�y�"ҘIue���N�u;S2�������H��8^x�=^�����ӾӜ�����/n����'f��wݰ���`6۟o+��&fW"��)i��#v(��d�LGu���u�j!��OA�F!�Ϗ��e���<F������_i:[�iK��I���E�˺Z
F���MW���oy($��1kV��Y�g������]�c�C�T݈0�mX]yw�����Qq�������9tmg1��p�?Xl,E��,��N5vw��l���ngD�4c(Ɋ������RFJ�@��Ul��٤h�z�y��T}�5-�4D�[�[��l(�i��u�ː�ُ�[�f�V���S���FY�n�0������}�q�%��oU�-㤷��U+����o�O���ӗ��y6�$�/�`F)�|٠)��3���<qy�8���'�wY���g����� _��w�+�Dݹ���ir�"��H��x?`�7��n]����qj��\������m��k4��s��\�?n9GD�I�����p�\�*��:Yr#�y2>"��C�H�N��f��:;���VZI�b��n��15P�C�*"�T�~�\��_$�� �7~��Z����sV�29|��**��}�ߎ��!>/��ӉVҌ�v��3�0��	�¿�?���b�ġ�u1h\�J@��En� �u]������m�Z�=�I<NÊf�%���?��Ǡ�fs�Xؕ��Y��������33.i��-F�
KJ6L��ڮq�I�J3��J��hV�7<v��dx��+��5֎�wr0�8|%��2L���6�㡗s]AN\�X9���6��qe�a�6+�t�������UC�E���_�{�\����|�V��{Zr�)�����%d�s��"���Qa����"z�Ȫ�>����OK��S����n?p��.'��u��cۓW���E�o�fJ�j~�#��7����F��qz��q4�� 3%k��Y׭g���u�����{ߺ�14G��"�����kǍ�'xm����Cw��\�j�  �[	\��ɡ���/י2Dؖ<W"g��m��?XlLOx�LC%��p�|���4�iM�"���Up�P�}N�5`ZF�|����;�!&>Z���U/pH�������g��^ѩؘ���AY���+��t �;ў�{�'�U}<q]��=�� ؐ/ �""�5��S࠰\���Cj��G����?�K;2F#��ݚ��P�dR
v����Y(���o�a�T��5����GT��wu���ॣs|+-{d&b?�����^���f�+ѩv'�wДrS�{'��
�b��\îT�iz1��p0HU�'EI�$'������m񴡹�U�>\؞ ����	��x�d��J����Ri�ѩ��Oc�O���E%��-�M3Y�b^+�$2Lk�?~̌� ]�V��b�meC"�k�2�KN�q�Cx�랛�qN����QmKA������Ӄ��ڭ˲r�&��U(���,0�,rL�����mװ
1�z!�x]��V2x���Ȅ������ޓ���z����H�rJ�a;t��n�vl�\�ro��BH
��q�+��^Shr�\��Ƭ���Ʉ%��DxTĠ����.��Y����<Y���L��l�)�l;I��r�����ˠ��<7���ʺ�M2w����T�bh'����s��:�!	�z�F3���J�%����5%_�^�$l�&�t[�2F��g+���;Y�/���(P۾Yp����T��Et˫	�rb�DOZ��S ��7���^~��^�;�izK����utio��]����X!;(��a�e%8�րփ��2�C$;��)���!�'�7o����Z����@݉G]�כ�ȶ��V[��_[Y���V�A�<��k�7=�|�֪mQC�x�౲��K�T}�:|�οǨ�CWW��q����+e(���F�x��m���b�Ƚ�Gy�
u�!kl��w� ����T���;K�v�d}��)
��7��>{B¼�����)��O3��K��1���\k��g(i��rr~�ؽc��+G�I�j�[��nB�ֺG�y�����Y����D� *�siқ�*�tAzG��Ф(*R�Ҥ�t��B	��R�	=��z�����sfwg�yfgv�eG�`<O����-��j4��nJ�Ns�����*��T�j}�������9L�_�#l�� *��Қ�y���+i���o^�J�m&<�����u�*K�}'lYR�hD���/9�W0��ĕ���;���3ʨ=�7Or|4��ݔ�"}V� �:��U�o��oH;��>��𫴠.�?UAfǚ���WM�C�)��� ��Ld��c�P������80,� �P d���t/�N>t�ғ*U����},����O�����;%+�5���2����j�#S�/֨j�4���[b1�#�n#Jf'��r��>B΍�k?��X?����f�>'D�=����g�&�wk�u���)�Wϒ��qT@M�|#�PR}[:��y)Oq����R��������$��H�*�f�Dd��ùyav��@��Ã���石���=�(��D��a���#E'��ς��H��Y+�-��*ׯߘ/Pl~�QKh�]]��P��<�C�����V�S�y?d\y�͗.w><����d�]_AG;�p�I93sY�z�����s��Ʒ2�iR�j�VpBf�i�5a���5���숷6|��o��F:��a#�M|ذ�F6<:4��f�����({���ѱE����a���K��c�!g��~p޼׹UYi�|��.J"ۗ�W������G+�cR�����@h���{�Qe��+�^�#5K7�-=��Y�w��h0���}rٍ>�Wq�H����X	�``��ηL�Z&E���bX�hi��/�������hb�4<x�<m������}z1�a٪�����ui��e�[��w-g�NR�*�m�E+�H5I��,�T�byA%��t<�������%Ӕ�?��7Y��Z�ĳU?s3���$D��%�{���5�~ �3;{��׫��V�Za_�$����_��L�f�O���oNg@���Ѵ��2�Q�R��5����Ρɣ+��2�`]�����
���G�O�l�D�7�z��ƥ��~�U,����E�*�:�o�_�L��t?G�n�?U�+r�l������z��4/%vY�����s4]o�[��l�NÅ���Q,ᒕ�kC�T�2�kmk{۲j�����]��?���d??xb�ݴ;�N!�,>�z��=%E�]7���_S�Ôb۶��	�2IK]�u�G��긒�����z:���7�Դ�S�4;����H�Ȟ��}$�U�6��<��֧:��GX�ۧ�d��؂v聨���TI�w~���K���[�xW�^�����@`�hHkr��[�Q�%�,�)p	.�v��[�0ƥ=�pH�����#6J�ŝ�w��v]�V�{ɻ-�����b<E]aӓ�L|��(q��m^
��&�RqU���y[ĭb�ڭk���g:����Yi���\Ӟ���z���7��K�?�PrEyziD!i�KH���*�[�$��́�R�8F'�z��}m�S�Xk}��#'3+*�Dt��ܷ���)b\v��7	 z�@�l�n������rqss�g�`;B�u'n���T)v�W�Zz���Э�/� ѢT��S��Ҧ+��kSv�xF��J�8ϖO:{N_5:�η�
�>��y�靾���_z��bpe��.��� ����z݉��ҦVL��ұx����!b��>�z��v�.�(t���B�L����Mn��ó��o�	�42�T�B�m�As���<j�%.�T<ؗR.�!�um31~��>jFEl*V�KqF% /��NoQP���2��
�nB%�z���.;Nq��F���~݅�����n�'��h�+ :�,:a�٦����1`íg<$ưj���=�7�p�;l�\T�p>��Pq}\��[¤?kY��*�@��,�o b憭Fb���ɓ�	��;cKx0�3���n��u,k�VvU�$!鰠'~>6,Q�����ס:���j���{�y��U UT��#�&�-�|�AyE5~BP�Uvm�N��x�r�tH��i^�L�D��5��{a��q׮�}�bK%m����Kx7����m�0F�͎�}&5Φ�!g���V\9R~K��T@�9�i�{��e:�&��3�U�){>8�cX�g�huY�9����B��z���Y�9��������5Ȱ(!y�_6��մ���n��V���K�X�>N�樛;��R͙�͉B_�#��c^�^�Go�k�A�;HB(?�q��1�=�l,���ߗU��ouY}iL�?��9yRt"�2��D���g���E�����vu��ss{���^�_���ւ@�RD�B� =)�Vy���vNq�����9����TY�@�X�7��SU��鍑�O�X�Տ��������aʭ��1��h43�,�Q����c���No��7?���c?�T����M9F�4�#!�;,���Y62X�,x��.�>�ʟM���s��T���Im�YVْe~j(5�O��>����A��'�d\�c�բ\d�|����l�'��EY�\�hU�C��1bgS�Mw���Iw"��k؆��:`�&�����P�i��R&=ۊ��?��jv|ѭ)b� 8/���|�l2�JB2�RW���ȩ��>�J�����0�����x�Ƒ���[_�G���eZ�p[ƌՋ��ݖM3��Α�Cݏ�I"c(s!����{�ɨm�>�$�9��E���>����;>Z 7`'�1l.��.˗ݜÛ9ۛ�%ҁ�9��l�>i����w�
>�5Q1O����혲���PLy�yk�y�`vTO�H��Sx���O��0�����~W�PW��R��zBᓒ|�,�prh���r�A=�K8����h�!e<Q�C�c.ĂApd(b�5���seK5�!��J��S�r�uN�vr��"`��ڦCvF�W�D�hS�M>ԧ=�a{�`Sݍ-�.��"����v�1u2����a�����O�L疎C8!�l���k��P��YKk�e�x{�pꪢYٮ��Li����O)*�}���N�_��˲�r�fP��n}����o?
X���t��q|r���}�����1�^���w�)���>�᳔�yQ�R��RT�ҿ�SK���:��KY@ �n�͊����M���=�����n-��U��v]w|Ѿ�׾硾�X��u������݊q|}����Ψ
�x��\���-��zOL�K�;����5�Jfk��.���^"(k��*��꒶���]^>Na�E�-[c�on��sky�*u��P.�jse����St�ѥ��m��u�%�����N�U��ELwV2�M�YYU����p�� *�����EG�����-��9g��[`]{��B'q@�DS�Q�<��lڜ+�u��=�a� }IL�������'�=��^�����2o���lU������!�G `e��4��sO�k<8Y� ��]����/��2��in�Y~7�kr�N,��W�{���Yo���doz>�`[,�9z�.���eO
�$�����tVj�VU]m��k��Z�N+@a�k�V���;��O|�_���/?���l�qL�~x�B�Qh�+ptV��р�P2G�f\�W�2w7R!"+�3��<|�]^t���6~������.��NG��F�Ǚ�>� ��u����s�-^�(�(W�~<�n�k��i���3���(J�.�;�rrr�,>β24����(�	�嬮��y�bTB��j���0����������3�>�z�(�Զ];�'ث���4����h>|�l�Ԏ-��5�j~1Ea��'E��9��~�{>l�ܿ����*��!F\�yx���k�T�}r!�aAa�ʭo�t8Ek�ԉW��^;-�/�{ZY5���f}�$Թ�ˎ�zk�<$���Ѿ@*�`̤�57{�~t�kr���V5�YmN��j�l��M��w�A���5��ٻ��\ۻJ�I��<1
�$o�A�'�6	�%��˹/�9��N���H航�EB���-r�����/W�5!ZxrO�"4'��wO����	sc��Ө��fZ����e�1���5���:ӻ�M��C'H(��~.��LԨ,BU}�M"I9�1׫C����G̗�*A�f)��0�+Þm�w�\��YJ��( 姞��+U֫dޣ���p������Z�c�� �O ���$���lp��Sྜྷ���R'db��7�ˊ�S��yO���� <H{�h�sf7�Y����]���>X
F���#���o��R��~�l����� � ���*��V��N��hi� ��i1�{'a��RQ2�Q��X��
M���Vmt���W$�q�	33��䥥F�Uwd�.����y������w��b=#�B<�*_窄�=$c����,�y�{�B'n��J����$I�����%љ���.��d�ƠÕ�e?����FP�qy�vq�)oA�j����fm�����!夊C�� ��='� ��2�w���`��0E�c�U2�º�"Z!.�-�E�R�f��6����� ���Q�"[�ں���מ�iz��J�8�\i��Vl�y~������1����s��f�y����ϱ2-|���)T�L��P9�s���&��<���%Ĕ��%��Be�0�,�m4�� �u��S'�iv�y���r��׶X*��1���v���z4֙ARg�p��%/���S���.k���?\��
����ٳfjߴΨܡ^��Z��pX�*�1x���fU��v�K1>	<c�mKqԈ-m��E����@�>�	�pp�\Gf$�{��f�U��ʇ\ZBn���h��j�W:�O��z4jMc��a9�9���'� �� 0�tMה%|��s '�9�鴜c��#��F��Ƕ%�����J|�B{6i���NK|v����������V i8��*���[j��7-����s�/=U��mVO �l~���T�6д��[��P�U2�I9G1ʩ'AǏ���S,�����*���}��Ad�=��Z��.f^�B�檲\$�z)Y�[�fh��v7���^f����o�ӯ��Mwǳ�F������.��K�Lgx�n�M!���p��Ś��*x�'�,�zVB�AQ�oIC��R��K��pM;���t�>��Q8�u���C�s%��CԴ�$i'v-b8W�R~�tMs`�񂝔�z*��(�jl<
)�����JK�\�qt��s��g����E�pr�8>�P����.�7�?�~��/����^%��?�{iy�YK����p�F�H�4��r<���Ղ�ssl�S�ƽ���va��i�2������r�}��֪1�x�s�5��:��MJ�Sy����
�0l�\d���	�����ܡ�][A��V������ A��>�Y�\�u��;���|l�k����4iʐ�d>.|�]	��c����\Q�2|W�!z�c!��N�����;g?椖4b�B#LpBWߴR���ͤ�F"����j{���N`d �9l��憻Cc��b�LG�l 
6�v4�\��$��45�S�АRŴ�y�D*��9?���~��ڍ��9�T��ܖ�CkhȒ���}��K���{�q���<���Ӳ��Mj�h�����[3��>���]i7�{l���Y�������謞���~�)ķG��g�����7�x�:�޾�\��+�?~ejz�E���;�>��-V� �]����,'�|��7�0le�01��ͫ!�(�9O�n��I�z�j3��첲]��SC�O[�|R�&�����9��I���G��vV�!*o�V|SȺ��tù�⮪�mn]�~R���g���:Ɉ���\$�依�.����;���f�õ���d�G��/��7�>6��!0���B�w}޴�X<�V����*G?�{/�tY���U�2kNqUp�
�3R�Af [�����?�ꖲ��l;i���n�sE^�^$�=,z�8TV���r�Ǵ�&�\�J�R4)�lV�h+�n��ģ���	8)�RXB��9�9^-b��6�VP�Q.S��-!޺��Rg��흉��,��%��v�����kb��4<� ںS[j����?��<'���%��O-��2�9�<ļR��h���
oib5Ϗ��AY�]lT���Mp�p�$�M��>�ʉj*]քjЄn�T[hu�pxD{�Dg���l�)I�����5`j�j�a�Ok|�u[ ��*���a����Y\��I\w��s���Q!�,��:Z��������)Ǫ�]�wo����'��j~V븁Zk��FM"���T<^@X$��h���� ���_���%t�s]�]m��C�`����n�S'J�ةj��0Q��Y/�,?9�Qag��NzfI�?T"Q)�p��=�v�iDYѓY��mfn�}��T3��Sz@��յ���k��ʯ/�J<�r|XP��R�X�ϛ�I�x�M�aa�u�wy��_�<�ܚpF9q#�f5�%�bH���Jq��W��u�/ܿ�0f�͜Q��r>&:��{�4����X�՝X����F�P�ڮPR���oz_M��Rr���p>�T��_Կͭ�{�E}i���e0�Å4������3�c����������|X��+C�D�Q����딿�S�M�����߱ۺ�_Z\D'(F�-�c1�z�?f�L$/sO,[��v�:�E6V�h����F��_GgȐ�p��x����2hL|�f	&)T�u&�zퟺ �74�Ң��Uq�S&���92275�c۟��7�f'��IJհ�o=f�Z�oY��ϽKo�����Y���3=<��C���f��s��MWgX����AϜ�Ծ����]���F�Yr���b�
IhM�v�8��A֜��8��>�c���O���|䪝Ɋ��覱����l�*aR�U¤II"}Q�,W` OIy�,�֪B�j�`�FKʉ� �Uδ��}��M��1iF�~���pa�Q
sw��"��Qh���KX�"���i�ԹF�f�3�nQ3�6�x�d�c|�SÃP�6C+�����=���6�c�#w�/�B"���JWe��Z��K��
"���JRx)�e����7!��nN��֏jw�K����4ȗ*�Εk�V��W�#�ϸ����ڒt��"���b��z��W���?[y�=���3ؼ݇���)M� ��ҏ�/,���o&����OA[Х�S�ک�z#k��a��Ψ�`�|bХJ�Ԭ<s��o��J�jX�(r������ Ί�o=A�(ppD�<Y}Mԓ|Y�"ohK��^&�JK����TŹf;����l�Q��O��d���m��^8����,x�?��"#��hv5�\���Y����#n5�h/��X\U�-n���Uy&��I྾�T}"����#�Q��&���[��
%�C�Dai5#`�a�n8����^�e0��b�cf�~6�6�W�Kֳ�ݟ
�A�]��� ْ��!*���9���E�n�}d�} #��pĲJ�$���pvl���`NR�
���䁒�3)�n��S�j �p�9�����b�)&�v���4c�n�q�m|�����b8;�i���A�4㖉��d��������kۜ+3��>��=n�:�DӺ�A���������C3�
r�2�E���������j��`����������7Eu�d>А�(\�E�����e#�$�IhH1fv����ؐð�cͽ��<���K�N2#W�kNDre�!v��aTB"EM�Rw�Ϫ��a�F�HO��ʆ��#Gg=:�	5 �s������&...���/���˹����r��m�5&>&��J��ǬW;=ˌy=y������\�2=Ǵ��ʄ�{�.���*9�.)��X�P�q�~K"R���L٩��.�����iT��j���2�Fiu��g.7�����U�\˯��q��I_��xz
y�R��ARS��z�\j���q�u�ӃJ�(�W�G��&}퇾~�e0��L�My8�{�ҊUoX���;�購s�D%`��E��V�S�nk�r
@>��˪�~tK�=:�MM����뻥 �s�7��E���X0L��V���^�|��@̩��Xi	����8\d}	5iM{/#��p3}�5^!�c����\O�����a��?J�sa�M�/6J���[�qL���[���4��|wt�q.%e/&��O*u���1����jI$�q������<�;(;/� �2%e3_ |M���C:Iyi��7�3��С�Y�{�%pL~�4�7��0�w���6��L���,y��W��޹���xB��i�/(��$��i�a�n��NT	J�ZfS�k�$rX�ߐ|��cb��h>��~�Q Iy��^�����|�c�0��ӝoZ�q!CE �r��Z����GT��D�N��X��]��g��l0�t���$�df��vQ�\tr$��|Va+��x
\�}�+j�;-@��2Rh:�!�Y� �O��YT��]嚝��� �Å|����?K��~FC=���f����32��`����n�~��<C���le�H_O�@�S�7�~�Z����1��f���u6�zKa�4�笽fN����	@��������Z���fF83�n��!���!e��ɮ����;���o~��z?Pp�-��%�R-"yFr�ΚhZU��tg��Ә7��5n!1H�uXk?4L�B�hi���0u��
qy�!�^b�4��P�F���3&�r��{S%���B�ڰÝM�3�١�a��^���{��J�^n
�;T��9��R�w����u�������Q}�)�"n���J���/
]@3���w�m��<���U����L�y�^�?��y]{��H)�~0iw�ҪR�k�����ۯi��L�,ў6�"�g��2^���]��q��n�c?��4�
���p��Ui�G&r[	��w@�x�P �H���	���ů`5�v��YK` 2���ų�ſ���b�����7/[
���s�o�L!%�d��Q�S��#��!�w�/�ϓNRW�%L�mw��+'S��8u+�>Rݓ[P'ڶ�-_�浂�DiO�}yG�T��ˎ^?�{�@;��ƶ|s翉k�]b�|�y�ͼP�X��S��]���e��� \%���n�J�=��nTV��MQ��rJM=Բ*�B7deRQ�V�-���_���R�� ��9\/X���U�i�"������e�u�g�A# Ws��[�nX�D�/�`���1`�����ü� �d xN7-��n� ��|����I~ ����P��%#�*{�)d�G"^S�Qx�_��SK3�R4����!���Ct�֣K���Q���G��8���߷��-t��N/�6n�d��L>����L�=K{���u��=�L6m��A�E�����������<����FTI�ګ�������w�m{�����焑�7���@N C���355S7��i8w !�~�v
>�KL뗪���~Q���PTI�ٳ�{�>K�T#���N�.?N�l�h����d�� ��~�"b�e�Ƅ٤�DY��^�|��E���ZF�1=��UqP��YK�N�������O�����Ю�n��x����m�~�k�B�r{e\_;�Qf8�n�O14�2H�'�Win�$#f-����Ҝl����w(j�mml�����Fl��m�3Y:L|�&-}��(�X�#��=kR~�u�Sܗ�t&>��F�߾���>b7���%�K��M��\��s�w�N���a嬞�M9�^�|ز���K-�qz����o(pwc"i5�B����kLhGD���u:ڀ�"̐P�_��#v�oG}���ϮUP��r236��-q��}�NJ��u5z{{��o&>��]~~}��ݽe]��<� �YX��74 z�պ)�%�a$Ǉ�t\k�-��*�$���hj+�O�Ty�����xi��,(h1�͛7�����b�0���l��]�8#�F3�=F�K�S-���30�:X�En@����NP8�B	�?�oĈD�E�7��T"F��~&މ��X�c�\v���V�ͼ�`L҈�J�y�g+R�PC@=V궝!��e�M��A0q��syu�`nn�1���2�@U�B��ᨴ�u���e���V�V|�V?��P�-~�/����2Ѳ�x���-k����`�1<=;�ɱ8nP��'z`��ѽ�~x���I�=�jYI��Yj�n�55z�_L��iab�Y��r�/�sUۃguM�����-OzO� w˓�V4^����x��\1
9q0����8�OǮ5	�iɚ�G�����W4��ġ���?�5��������o�2��!1�*#
=��M�	ֺˢ��1[*�{2!0L9n�%)R�C��t|��ma'��hή���m��Aһ��"��Z�}((I_���zf|莘pFB���XڊyE�5}`a�E��r���M���Kx��""6�%ޕ�x�B���b�ҮV����Az(f�%~ �h��<�PAn5���k���*�N���\2
\����x��̐.������ґ��Y撈8�m��+�5B�'�,��)�~V�7О�3�b��~���i�h֐�i�C���$�{���=6�pة�_����ͱ���+��'���>J.|p�3��}����^r?�A�!�t�Ŀ ͑h����2�Q���'���e���`��o��mF��x}�k�������	^.#����Jt�^S��ؤO��O�;x�2.رtFJ��؂�.G@��q*/;�F�"x�%Ρ�����Gǵ>��b�����nt5h���Jܒ�,��xAU̜~$��JLb"�,����|U�X-w�5BhtܨÙ p�d��]$~g\ Ɉ���)	�C�ʾ�\B����H~��󾽭�{�c!�
`�{`^�,���]K���siNui�Rg���A}$;��a˛��΍'�����2$��5_%��i�A���#NyGt���Tњ�)%��I{�k����P��5Γ�� �p�L�+5Өp�^ml�i�-�;�t�s��E_l���ZqY�\S��Y��hcs�/UF�n���z7���\|��!E3�>����kC�m�(��>ND�6n.��П�M����Z�Sꀵ��r��<��O���Cd�=	�;�c��K�a��H���r`�iOѡ���[�<�/s���/�+|K�r14}[+��1�|0�g�v�7b��Y�=�v�����ȅ��s��e��b\k��u.��C��Y1����Z髹��l"�^싍;���V��g��)Y!�:�.��d|��S���wˠ��`��`�-�ϧ��W̆�_�8h�ͮ�� ���Nss#t[��xqГ�&�B��T��03L�]�Q�J���Єrw�}(�'�<��;1��˂�(<9Ҥ�c�/��9�B_Y�0��r*�ɭ��*��ݗ��!:��s2����둠���Y�-ғ�(�g+��Y��~'���ۮ�$�J���ذ06���2��%]Km�U/�G��o����Q`a����V�_�>PQ\kX��u�zd�������zD�}�������ԧ���K�=]�H@E2��~�^:�3�#Ӕ-��2�2�Rq'��NصR�Jאb:>
ǯ��VmD��Eٞz�/����@��u�T}�2Z��<�9�I�!uY�k�"�����q^��]�ao��O�B��Rz��)yH)�K���wy�r�_��8dj��=D>hf��N^ÔD�U�����>�~	L2%���s����:���;]%�'�jd�֖��t��x�Ζ~<�&Y�9%z<�J�M�Τ��!$���d�o�ʴ��b��^�KW�0ĩ�ax�n��=��f�lx�%���j�w��bV��_��.Sz��!�BS���<5�F�5���pRKwZ��S�Ub7��v��6������@�w2���@�c6�TJ�����lT�5S�&93DMl�l�|��GK��b	!6U1���
���ZZ��W¯W�����*�.���� �!�x����u�(��H�/CWZ�(W\
���CI��u���ᥧ���\.�̀�w��Mk`�0Os��~���z	c��rL�eS����R�4�f��;6���Bm��Ho>Ar�j�|ᯰlxߥN�M~O)����| 敇T��ț'!�\p�oci������%�t*�RB�w� �`�����%�Mڎ�t�%�bF: ����U�j3�{�y󕳾e�d��
��gN�(S����>���v�2Ȅ��G �u����t�Tڧ�Ŧ���.ױ���9e���g�ݾ�<�?�3_\)ͳ5(��"� 1F��V�(��6�cE���.�(d������磋�-�os�[��>�F7mG�ӎ�\��xE
ڹ�������M�&]-jŊ8����c(���z�^�j��w�K�`�o����K�-+1�R|����"ي���BQ�f��>�ޏ���F�w)I��`Bٖ�'���sp?���:�{��������۠�̌���L��mxOD��y����w�홻ܾg'��� 7o�QF.�/4U��m�8�ke��+��*(�Sb�����PB�'�����'�����`����@iH2��X(��6y�$�+��\=ՔP��e����g��:�d�!��ә����iҍ!����Y;-��3�����Z©�2��+^�ؿ�i��䢖 ����W�n	�3%�a�j�].������dg��n�N�gδ�4Six�6�>5�#���x����s�;��2��^�p�_���6���ڙ���Y�}$nD<��_H�.�حu7�k���$�s�.T;�ԣ5�%��\ �uh�� �,��o.�2�'���+_+]/r�X�6�&��ڧ��i�����I�׵�D}��R�bHy^-|����	Q��X�Xڭ�~B����X&�q����o\^����RD{�G�uȏ]���5�dƅk�1�լ9�}�SY�Ӻ��u����ag�
�����=��/�L�Ǔ�}�9a���WA��5Ͳ7|մ;�T�><q<��$��XO�ц�[��"��O��$+�-e
��G�-U�["V�,.��ޤPP!Y��5�V�1~o5Qegqَ�1���<� l�_#����H�W�%`�A�z�Y���_o��ƺ�<g�a�&�ي�.���3_���RI�8A-��!��Dq|Tƻ�Y�`)=��}faI�ߙ�v P���vB�����s }]�	hZ��ʹY��f�j2��`�B'�ʵ=WL���
T�gnr����ߠ%�U
�e_Vb���?�-�+ɣ�����LYu4Z̿�%��(���us���V�+!>�3x�]�;��K�=A)�LƤ�]�zlG*w<�u{r���<s�)��_5�+=�֞'6�e$�#���=���?y���֋�8� |k�~O�wT��o�4��ٱ.m�"�)U���(����ӗ����o�H�x�(,=Z���)~]��䦫���Q�4���b�Dbym���y)�9]D@�hג��%����F�ۍ�B[C'*r[	�S!Rq����c�OW�??s����`��B㘼c��µQM�YQL���ѳ,���~>i�D��K��A}t���oW�Qk�l	[R͋Wב���U�q�7���>4�蘮��}�M�w�V�KPFt���U���B�%��lFO��OcO��8�Z�?� �R����0�1�	d4I&<	����ݳ����7�$�('�d��@0�Z%!��
԰�L?�=��d��}�+�MYkz5�dGt8�C3OR��[�T���"�
M��:y⾇7L���:��E�oڤ��W�Z�����>����W�F�|���-�zH���O��!k�c��%�=I�<���7����y�����6;��SX�*���#�G=�~P��1��$n���^q�&$�`� �[�Vڰ�=�z��z�QCb�2��]�if�
����ů�%YT�ǜ,R�r�3��C/��ܖ&��OOY�0*x���RO��Ӗ�/m긴�����������x�L߼��sHu�v!�*�W
�7btO��Ti�F���$�-�AFk��G��xG�/����&�T�9v.:YBbQ>d�{j���i��[&�'��_ ;��{��z��]��&�{�Z0p&a���H��!�"���v.�<���hB����s�#]�9;��T'%��t�'����$�Jj  ���F�GL-K>�i51�2��6Sȃ�k3x������B�>��v�	����� ���rn/[�����L��\)qR$7�䓩�D�h��0���7��m)��k��T����6��vG���$�ѷ�6Jȓ�h�����~|�X�9�:���G��[�g��"�M92Rԃ;�6t�}����C%jūwI J��{���}��ߡZ���s�����){��D��V�V��a¹�|��b� E9�Y��]�ƥŮ�Ƿ��M��߉,���yTn�kP�h���iBV�!{�>��Q���+wEVY�8��O4�n�U��e�0ԑޥ�ea�@��J�ӂ����_m'>�)�J��1ɑ���A��p��WO�8�-ʻ5�AK�A�R5�u0���1�5r�0Dymz�W��4z$f��]RP���u��d�q`�JY�l� (z�\����PqE��)�\�����G��=`ex{R���/�����>�n�Zfj*)2�<� YN��</��S2N�ͱ���W:Ը@Ɩh�p?�4�a�z�ljE�sk�38��.l�FE7F�`�Ɍ�w����$wPP��KO{\	Xb�;m�MQ &3�a�2wyfҾ������qO�-����K?���+,..~vws��Ц�5�[t3|K+D���<�S\F�'��کVx�ފ���y3෧�
�L���� z�㋔?�^1�!�J��V#
�1�"��#���6�������G1�콃���V��WC3���f�N��=�O��1����[��\��'�d��W�ƻ,�XV��?� �]#�복�A�Q�Ϛ*̷ӽ�7f��|��^�pb��?�@��G��%���{�G�'�-�.�,d�K�)�nn������:�fƭ��Vj���4�'�ԏ4�A�O֤5j$��en���2r#>%W�}���؇N�, ����*��B���w<�^P�@=4m��'�NKL�����/�aT�z�`�>apsI��y/s�*<�j����.�O��`��+�C�^��7<����u"Иˠ��L s��G��3���!MZ�ɯh�J���,�<�*�X��� ��r�?�Ey!��كV����=�	뭿F�X�g�G�?�/w�1Ag�o�l�Z�=M���ڢ�k�Ι��Co��HЩ�&�-����C_H�ǳ�9i���#�-p��%��H���|E�(����[�Q=7�<q�U����Qӗ
T-���N�X<�����s�APT
��1����N��.[#΃d#�F���g٬y�*�ލ�@$�x�K�\^���@㫂��}��J������mB�yUٱ�n�v 8&9����ž��A]��CG���$)"A��ˠſ�+�KB�"s��߻�����z��+d�Q?yQ��//fB3�Nd����̸O�$�W��`s���E~�V_�!B�O
��h����W�����n��R������7I=��H���<~���c'a����ϑ����K������v�.��P4e)qhoC?V��W�Y���S0��sbڊ����74�Ɏݗ���f;d4�"Ϋ��"�T�d�h	�+��%+KP��N)��c�+�w1�N�K��d+�V������jħ�S��f�]�z��������]�����,����p�z�-2��v��9`$Z��z4�V��Y�l�XG�c�J78�n5���˧Rξ��H�4Ѭ�c�uQ����A�b�`'���(�ju�����b*O����%����v�L��7]=�Ѵ�&`��\&(+�Elz?6x���p+z�U:��D�����;�z�)hc�ʶ��	q`FэL4����緻������ЁM{G�N631��#����0:>F��D���?�Ԉ�Fª��%��LݡJ-$�)��L���t7XY\���\�ď�jYBg�lЅL(�NT��r�@1�<�6��O�"�b
�=Q��Ή�5L���Z՚S�s�������M�k�N�X�^	l_�/NP�@Ǻ�;J �H���f�d0����ŕ���p��G8�w�b� ��)8K��D ̀V�((-�|����aVZᎪ�W=�Ƌ�⒫^��S)W� ��r�7������-pJ��"I����mb�خ:�V�}���jR���[�^?? L$�c���WG�u2�|�=/Lv�'�=�n������%k�$��%|k'���G$��IY�S5q��S��Q���b�{�D!/
(����xv+�.�I	h��%�f���~��
ı�����z��$%%S�C.F��N�2�����]�5�=Q��8�ZLm\ɷ��4�,s!�2�o�k	�YГ��(yt܈�[�WxV2�?0�'?��2�*��"5�@Ww������g�7��$%��{	�^9�����-69T����{�M۸��=ѩ������2א,�6AӇ��#EA��"��@|䍗2˳����=�}����F�傖���-���������A�o�����@(KZ����$���#<��4p�5��S�>jbgi����ظ@��э�oPA������팼�2�2��׮�YJ��-t&"rl�44^���⩽�'�8	����{�X.n
S��gWؐl׳��S�_s�ϟA
��O�E�wJ|͖����\J<��FɈB���l��71��n�`�u�W=�kN��^�,v�2kGF�M`zw�m�Q�e����s���Ez�"�2���V8�|�clơ�͐e$�i�={��ܚ�N��2��U<NE�m�t���3���q����J�iF�}n�Z�$ە��������#����\�GSƯq���Ur�(�.n~4q����r�3^��@%��\�l��`�7�j��߻P���ε�%)2�K�/������l�ԪCx���\��	{����D��������I���/���<����x�{Pw�epg��[�V>Ʒ݂B�!'��3s�T_k�y�Eׄ�bV�Y@���( 9A���d�%.�("y���d�9��9�%Ò֕�d�����u�Wu�n���N����	�}�~�O�$�=r�����x�Ҕ��ft��*�k�"�eW\�G�̩`�f4�J1�7tw�a���Ǆx��Α���G0�����R��@P��}���;<�X�~$z�1�&"!��L��S7xJxm({],��տ�ӛi0�M�.6��⡉Mװ �*�[d�w�+�BbS�Ӓ�gn��;��a떝x��E�spE6��{mY�.evt+��"�7Q>�IOz.�y�	Z��,��j����� ��7�.ގ���~D#`�	��'��l�g��M߿k�s�s�.����\i����pS5�	6M���6���n����ޓ��PZ� e�F���F���a�<��*���J1�4E�)�4=�GR5��� ��e^�;�z0^���sm!� "�(ȟS������:��¯I�¥�鄧�>Q��pU&�>�'���WO��V��\�:~(.ؙ���:�b#�{��-��9�Q)�S���{)�){3]���Y���=�r�G/u�U��R[��2=F�+[���g�j�}9�[���;��.�X/�f���1�}��qSƯ*[_�@Mt ���,�Ԩ�#����"�C�L�|Z*d����Jjt~��X?e3���Щ[`0�.W�Y�+�U�*6k��+�S3����Jo�+����>�3
�sJ(j�F2���x�2�c�#��X�Ձ/���H;��M�~n��Y��JY�}���is9N�3p3/�,�(��*�[�ٰ�<�z�Lg�kw���j^ax��5���H�?��P0#+,l���*�NM�:pu>��`��?-O�=o2�6q�7��G�!�\슆*Q�z �x4���'\�0Sc�'���
U�,^�Dc���VO`w���P2 &z��R~� _-DS�!B�'A"�W��	+b1�_j�է��?��ٛ�q���Т�ZVqX��S��6'���2��M�ccn�?i�ۧ��AM�j��ħ�v�"�Tܣ����vHv�0�݊�k0��wvx_r�WK!�W[�����Mp�*�˫��Ɠ�I���Q�������6���I���l��°t����	H7Q�u_ �8���w���|�]�$���8�r�oZ�g�ۀ��N����o�̺���%�!��u�a}P�!�糒t��026[�)����� �MK�/@F4 V�~�<Q���Q!�V�9*_E���������X������D�Q�ԉc�"�r|�h�06\C�������U�{\>�'�4<?��e�e��y-.�t��vɼ�����cw�v�q�Ӽ���8v��(̱L�>d�����!a��['��	�GZ(�m�� �i�S\dN�_w���zab#Ya�u8�P����9��7t���򲗷��ϯ&"�vw�����ѣ�5���7�M+jY��;�,2��m��*k,.�@^�rz�~���
N���8�?���ΫwT��H'0�o\�R��R��v���0zM�>������$�/����~{�/����h"!~�"�(�WSH�*t���%�#�3�h�
Fg^��F%�RP���d
7��}�?|G](,0�|�0U�BS��C��sJdT��2_u4R[��f+O�L�}rh�A9 ́��Ő�8�_d#��48�7�և4�8ع�����7���"o��w�|�.�ݛ�ƚ������"���t��0X�0a��:���J\�Ũ����a|��iy� �I����G`���m�RCo��v�j��E~$��8{��r���-k�� rA^+���i��>>�I��(CC7�1vc�N�]��.�*���M�w>~u&��+�'Z��/��;i���&0tMS#�n~�����ȡ�
��E�A���sۑ������7.�C\�I7`���k�+��3,>~��iW����>k�-q�ڞ���|���tT������]�*�d�kb����R[�OG��ۍ�}��1�ؚ�,�,'-`��ǅ���"�4���s}��󷎀�lҎ?]<��2�d���E�	������=�۫uFU���
sիBS� K%э���SS2xxGZ����S��"Q�f寢<����h�����:�]px#�=�H�9�"��ý8 �c"UX���I���26���4�ֽY�	�P�������s��.e�BL~r�>�h�� �i����6�E��EIir���&�Ws��R�st�\q0z�N*�A�{���B�
^&s����k�����ˡޑS�ԙ;�{5�t7��J�ILzXw(Ԥ�Cq�
a0�����4)��j{0�X~=�1�,�$j��7����tv�T#��xC*WLHK��;t�5&��s��;�y��Z��FP'�4o�m���
J���K�\�E����Nc��;=�{�:����dV�_��Vqm�C�i�BF�Zr��2ׅ�P0���?LOۯ����l'�$�Rt��x�����63�#�J�\ʝ�a�
�e�^l�n	��JZ5v:_X�Ha�aTecg����[�RYZZ�x{�~¦�a�_x�X�3Q����D*?�����?����睕Ŭk�ϊW���?bZb��P[�jAex�r4�nzKe���DڳC3�ti�<�4���q�
��)[�C���:�J�IE?RTT���5�/]OU��i����g�;�oJ��n�|#'�$��" 7RCu�]�v��B���:�ұ��>V��ͯ�����g�/̽#Q�'�\���^lU2���G_�G}Ԛ%��ZV�LY�?�NVڏ��g���N]��f�XP�e۸����O���5��=5���pS��=Kt~Z2�"��*�	�ި���ƶmIxp��H�,ahX:CC>��J�I�ǂt��m���ɬYB�EKK�@���+ ����fV1�*��1i�1�$�S��E���{��t�n�m6�J}_;��k�+��2�I�-�@�}!�Y�^�h�:�[�1��l���q��V�i�Ga;���y�w`Մ�'9�b1��O�����|խ�5����S3��h���/��s/���	5.,��xی[K]�iR���(��	�
���q�vl��;�i&Q�Cg�pO��6\x�Zp5'}�O��y0��J.`����V�I���v�^a���?��m����^��VOs)�60��6W�����V��wkG�0E�\^��2%	�+
·U�'�h�ђ����j�G$�h'�z��Ɔ|�\����"}�$��V���y�C<�����$����ES�'��<~�ћˉ�*���^�%��ޠ3C,p�'�ٔR����Bo�د��!�����u��?>_��eP�7�9#��T>W�'v��!�vUJ��1�o��?6ے!�&����񊊊���Id#�.����C�w�V�C�Aܵl݂���Z�R�����^Vc$���
{���d͇%�v%�봉	���{�%|a
;��*��mhb�Y⟟�FL���lm�$�"���tF������ݢ�I��g�<0-a*uo;+�>���:����"���Jg6�����Z�$����9��)�]F��-�������^��9L�~̮c��e1�5�<��ƀŶ}���DB<Z^6"�?�`�b[�JQ�&˚�����������mC\9�!�I��A)��i��9����s�������ih��u
�L�FN�{;E0:�ִN��NcHm�����R�/0W�-ˡ,;ѓ����%�=�����QF���_�����ؔ� �'�illf��7j&Ō������'Хk���l��F��֓!�{����]��[ڸ�M������<��AZ�:G�F��5����o�::1�v�J������ڒ&q��w�[��� S?%@��Z��Kd�M�B8L� J	�����Hb�������b?�\F*�Z�<=lxm����m�����KZ9��|������f/L�\vH�:R�7�X�
��Ѿ[�1�..�!;�x����e.e��H!:�"���e�im�Q\c[=�^]�D���*�o��,̗Ŕ#LCf�(��bOh��u޴e0�a�����o_��a'�ǔ�zޣw[�Hߦ�1�l��ʔoMUJ���T�����-����,p'�D��N0r*,({	br���A� ��%KY��焓�����s�!K�|ç�\�.v|���n�F�i7�~�A" �����r|ٯ>*��p��\���<F��u�|\T[�4�,���q�U6h�X�	cr����^p��FR#�nJX@C�˹d�-{4����c`����f�ذ�o�.��s����e ����l�6���Ad?n��"E$Jj��NH|�/�=(�`7��*�i���o��!q�l���T���oE���#��|�ǹ�c�����a���ߏ��:d�u5����������J����%{v�-_IdX!S���q��j.�j�Tvs�Qo�#�?T�%�Z����Yh@^Z`+�Eo�l-��6�ڎU�B���p��	��a9�HP��)n��H���]V.�.g����9텭�N�2L��Π�����-��}���c숙v,),��u�;��n��0��꟞��m?hTa���$�8�m�#�����b`�(��ȨQܨ��T?�@��۹yN&�{�2-���]��:'q�#�q:��?�=�tU��?�|X��Ӽ�l�X�q4��!�>��3>��׫�@QjC����f;�%b����_8�j�^�̬�e��/���.G���g?�(���?|��<
?�q{���z?&�÷Z���F �5�,��)pL�����x���{t���2ҹ\�LW[1C�ȋ�;?����' i���;��d[S���%�~��c��M���X����xkiO�qu�����S�)q��Ŗ���{ƍ"��s�{_)?@Hk�~�1o��x+٪.�n�Vh,�Փ~Ч��#j�7����L:/5� R�+��OIt���A+���$�rlQ055u�E��Tc��}�( ��_';�Y���}�~FZc?�&��C�J5��(K�2��GDQ�d������QCy:�!Ӕ)G����'kD�]�G�h�T���)������%m�������۩l2(����\������"�}� cV{	�,���5wQ���|#�����7�U�)�d��e2>b��\Ú���5wQ�z#ƨ�Sz�q�K#q�?ck�	.�Z{r��^Q��k��8-���r5�Y�|������������VE����gpp|�n[s�ɀkrڨ���R _NS���/�%���I�1�ľ/�/j|I�,1�\�H[�����f��h9�' Cv���qE��2�������ҿ��S���)"�&)��A��/V�61$:���m��"N-ʂ�}m��ā����7c4�/&U�m9��G�#� 7n��Z�?����Vz����xZ W}��ɐ�o��ɏޝuUZ�0p��|���Ǔ Jxh��O����Q}�����ܿ��R/)���^��^�?�\	Xr�*�*�B:�c���y`q�+C��{�<�p��;@w�́�8=x8���E_�<fr�N��� ?Vr��[�6p2���<�N�8zs��#7���0T2��(�����~�$-�	.�-��Zs��i���i�M�	�_�0������� PlI}��@�\��[�Ec2Tk�O���eT/����¹ԝ� �xVh���G��;��k����镾t�'ڪ_<�cK�1� o�h��덎`B� .4m�g̭�?.jq���6�EzS�	���_��M�L���q齀�x��~�@�\j���@��o(�>@.⵿��0�34N��<~]]�Z�6Y��'-�=���L�3*kW���)V<95�Mf�) <�w$�����?]k�5�!�ބ�<tӗ m�к�K��|sY�@�6��×/�Ӱ׸?��Ou����Ī=:���V�7#��A}������o�����sU�W�޼|�/��� ���/���_=���~#��� j����+eT1D@h���u#�.��1�0nbdj�ym7n��|ݛfF�c�&0���z�F��l9Q��Pe�2.�eD�<���<�f�>���w{�̓䬬��, Ȩ�.R���#�ςՆ��Bt�U^	 �pLQ:Z����H4���{y�eja�������_��wY�	��	J��0c�v�C~6������R:g��H'9u�Q����d��K��퐅�=���I�Ӳt1��~��Ν~<PY�����Q�M8�.z�~̐갴�nA�F�{r�~�b`��!;��Կi�lLXv�����b9�d����զ�Eng(�>
�(���2���ڿ�K+����)��Z�N�G~��h���I��O9�x�U��Nw�t���������7��Vݫ���sqY���n��k�R|�,[�N���������� w�}S���	�e?���g~N��j�Z�����-����7	�UH��JC�m�xU�á�5��#�[�X�J����m"d��̜�*ಈ�%l�<T��CLM��^-X�x�[^R셱7���
ڰ�d�x��[�س�<��\��g>n����L[�N��3�ul�.2���T6"]�`���F�L[3�ZQHN��{hX���K�k��R��2�T�|_��aAV'�N)��[��z����B�[� e��rr�[@�p@���s|,�M�l�[�����}�
�_$F)e\�W� ȩl9Ri]�r�� ��4��;r�R��k���5[��U�, ]o	��pv]ɓ��{h<l���xs�
���k��ﭭ�"�ׄh���J��V�����72;�^�.7.�2a��p���*�!���3��c%�
��;�G����������Q-{EO��Gl8.h%3�Ķ4�]���V�Y�!!���r�f�͍��~9ݷ��u�1M ��Ӹ�w}xm�ˁ��pU��w�oŜ%d�Vlo4Q��¹O)��crԢ�1��m��z@�'��a���,:vںe�^���IF��l�13w`�s�HG�l��lJ���f$��A�Ս�rާ!�:��j�qqa�k���dh.�&��p(urྡྷ��m��z��&��×�r��v���39��&$�*���o��SDJܢuP�3]���oT��j�Q��;�rr�`�K,&�^�-.!���LC�I8o�|����-���4��T��,��n͐�<8����~ź�3�y_��`��Q��bئe���Y��+6~;k�!��|����4o��	���L-�p8�~���T��R_x\�)��>.��������է��A=�����5���� ����āҀ����d�u�{QVtV�x�Wj^�i_�">Db� �,z���-?���`G���x�*�>�b$�V����[�tI̀�[���ߵo?�	�6��{��M�ϻ�{�u�g0%�LLr����ڊvS�~S5�����;�l��ֵC'ר1�أ��⑩���v�#s�ɛ#�s$�������,L�K�Y����<ƚ�a�MBF���W���"��O�۩��c�xj�<�ڙƑr�:��� Ԩ��r�I�ML?�%��Pf� ���@��B(AL�vM@tF�; ���o����(��7��:<n8�)lMĚ�ƅ۽\�J�А��z���<g.0�����Y�Q�㝼�{Alz�N !�@�[�ɐ>���T�MU�E���DG�&��M:{�"N����x D�>�ˤ�.�dV�oe���׭h\{:]g�m�\�\����(��#�ʈ��6�z�̜�y�7{���=��XY�F�+�ָe�k����\w���\M�Z+@��ե�Z`��r�z��)W���8.9�fk��P�?w�uX<�fXBi������c�rU���}�i8$��l�9 �[���ߣ�r'%Ŕ=�j��=s�H�8�����%x�x\�^2�\�03�@Ţ�mw���pi��̡��q��);䃻
*�_�<���m�V�Gƀ!C(G�i�yK%CPK#�C��f����H���i�ӑ���>�8H󢀋tZ�h[�x����Jm�.���V���|�_C����b�� %��D�-���InKq����;��f?���`�EvR4$�k���UU�)Ǔ��YX����2!��'f���-D�t5?6-��R��mR����;���2�h�DeZ�gw :Ů#Њ\��pE����x�9��[���d\�H��)�Z���p���)Ba�8Y����j#dZ�p�^kw��Z��`��4E�{�(;�VB�]yK�M?z�'��Q���~lh�b4?B<�P���C(�?t�iU��x0\��d�y:f?���/��D��Q웒��03��|�MH!�'���1I+Ї^S�(����B�5rU�C(���-� w����Y���3�mv?��~e ������P�pKʷ�������r����r�7�����o���5T\��Jr�]��I�O�����m��>�� ܽ/g��T�j
8�^��-/iy��j0Gݾ�=��,�00��f��k$,w�|�2f??3[��_F����� >����?{�1���Qf�w��k�/aT&��5�Snb��c*fN��A��J�Yb�NFJ�&[���|�ѪɎX��K
��r��Bh=-W�~i�δ��M!���਌e
;6�/�e�1�N�?JCb"�'K�`�Į8����V&�ݙ�j=�?E��>WZ�!���SLb�<��7¨:����(�V�Z���Ab��T��-q��RJ��6~����-�1�M���OBYᲦ�� H�t����L?�_�o	�gYt搪�
��`@���،y\��x� +&D2A��T�U���r)�u�1y��qO��ϳR:cM�8��C
,��b:�jnt��W�~���� �is%��>5O��ܨ}t&�?(!�"FVm���m~�cUJ�J�2���	
�L����7g67V��N8y��9b��"P��o���V�f{�Ӧ���k�,�.]��':5��J�c�v6k�����g�x+GN23i���d�ƴ%�5��d��L����{��� *h���{�@?�)���<��B?h%k���or�����o��:n2������ ��k���)��H�r0g!�	��t��n�z$p&��GL\�L$�mح>�xD*L��Q��{���j��g"T��X�8�Rۼٟ��������|�H\�IU�zy}�E ��?����M	ߛ?�M2��.~�`��<�ޑZ���a&g�pc�'��I��~�Y�V�Ч��"˕��q�𸌘%�\��W=W״��JgHUn�@�M@s==�s��%�sM�� `:��9�Kp�@?a
�<9e�)� 7*���(X̏�����t^0}d���葶a����� q�ޝ�k	��
g�k�7kFk���A�Y%�t%��OKm�A�Q�-�����/����,�����Гـ�K'��O�l � �aV��cI|u+koh~�/t��h�k�ޛ��k������'�<��+����������L�yr BZr��(u���+5��k��T�N$�_�0>q9XI�'՗�
����-daӃc�Z"g<� ު(��9�N}%0�V 9#73ZH��Ҍ��1�^nJ�� @�~��n��P�O����A1�ǂ�@ ��&3��
�y����A�����-�KG6�@�N������9�~�ge?�sFGz�?�x��c�Rӌ��v�zy��n��}-��j<Н�'�4��~��Ta�7� �/����P��G�cEu��;W�	���~�v����9�ZȈ7j.�zd��b��QO�.��NZ;���9��L��N�ʷ�����ȉ����y�^Y0q��e:�����V��$`	�-~�@�K˷���#�g�g��i���0ݦ�R��t�>I�?�f��X�)Vp��a\��"��h�`A�Eʟ������zd/f�4�j�N�R�Y+��\l{���m��cK/��	]��`���I��A<���<��H�~u���Rs�`���t��˥s�9���b�=�����g��p�@��n���c�e�'�/�2��q�� �����;C:�t�q#��Ee������%�2#Ζ�@�"ښq)l㓟1���XT)]��.�u�Fyٴ+��b�&���.�i�e����ڷҹ4G�k��O=���MS��7LQS�Ou�_ɮ��P����IP�U�r�$ܙ�+y ��Ps,�+��zx-@&��<��%n�^Ex��W�o�>�.KG���G��#E�A��W�	�2�c8�7b�(�59�^Z4�K��<K�>�@�_��P/��;1�����|�A�4v�q����X�L	x� J��	��r
���GM)_����E���À��B�&�܅����:x�hOw�ݍ��+���t_+���D���K٢8�rM[�!yE�`B�JjFz�������
u}�C�ߵL���m/�"P���1ꊑ���� ܮ�4��2f�BWfޣ�x�����]V�r���d�{�|+J{̺r���ߗ�_42��-�2{�Eѓ����pu�iܥ��(q 㱦�\ZZ�`�)�r���n����G����m�*&&�0�Jd�B8���:��IeR�$�o���M��e��h��a��`c��!X�\	�m��dΖZ�f��6j�a#M+�����U�{x�)C �6?s�N����/%��MJ��Ӧ8�Y���?F}9�xȉt���"���D7��Gi�;�V3���k=)r�b|��u`��ڙ�rǖ-Y��'9��*NV{!�t��޳�dڦ�����׹�O�zN�q�\?�=�K��7�B˺��8p���L��^N���}I��*�p;I�a�s*��߿�`v� ��_�#YNt�;�J��&	��(K9�G~O����s�1ÿ� �=��ca
���x!+����p�M �Q?����S�%��KC�j}x?�qn߄!^Ta����Ҩ���"��x�hڵ[Ĵ��m���v9ۤ���n�w�E���xk�,UY�BR���6ǆ�R���8~�ژ�
�bq\Z��.Xr�%}�t5�:}��Z�E�.���M�Ai5%9
�)E�G��>���P�?@S��#���h�1�='�`��Mӈ�I���).o<A����nP��!��:|����M:�����z�8���V8[��B2uK*я�CTem^ΟF�d*	�P�`t�WMx�]�&�YL�1E��������X� iզ���g���h�P�8n�%��uד�M�*���0)����z��qz+��ȹEm}/k*q:c����J�T<z�XJ5r��%��0ҍ�8[�t��l�_�0c�׫;����-y��7a��Ap-�܊��x�!&��.2f��p����jҊ4y�5�0�$,D�{�5`- 󨜚��3��p��c;�!dk��K I�����8Ep�c�p�Zi~�Բ��Ҵ��� �܅��ɾHq]m�r��;�|H���|/�f�Z���駠qn��i����%rW�}l�Hi��O���k�۰�F���Z���-wO�S��VC���i	���ԡ���·kC��cP=n�l��=51/S��(l'�	�|�ʬ�:h� r��u]�!樐y�=
#�Wk���~�&K
9�%�bF>a���.��\���Κ��y<�aUh�븣�a���[9�l� ��d�Ŝ_(ߠզk1#��`�Π��v.�%�U�
���":+?x.�tc¥��vy���h!;MZ��E��+vW1`x11���X���ǡ�����0!�v������Ǖ������T^�W)�B��EINRy˺�>ek�
4�5y�1sv�S]�d�psSW'�3(�YM+x�sz�4:��ڽC�5��Z���|�'(_A�_�E�Һh����9�	�`����p����?�1���S��?z��������(`��]�]ۆ��S���)���)����@��i�9QFC\f�W؆�Q+�11��ǉ��}���eY���ތ�=���*F��2��c7��s� �]3�G~v)"Q^�X����+C}7Υ��mхY=��d6����<�&ҭEQ·�JF��Pd�8Mب�M;�߳�v�K�H{�I#��1����mi"�%�^������������LL?�ҵ���V�z�����":LL�5�)�+�3ߚn��9A�j���O�<��\�nN���2%j�#��tS������}%���U��=��o�-�镽T�LX�J���)F ��@^>�Ǧ��/��(_?�m��'����B'f�����Hv����E�!�/t��v�44F�P�dٞ�ᯌ����i���������WK��/�������8p�4�X�c%����[�Zց[�Fv��)�v�-�=y�,T�8>�XY8h���Ȼ@M2:�Xa{0%��P��g\�@_�3�u$��$�y�+��Z٥t9�<t��F���d�2�=�e�{�s8"������8n��<�Ȥٿzem��(�����X��Q���wg����$�n�{�݌��x|f�Y���g�]
Nw��تjJ�W�Hp��]�
J�=���9]}�5ٻ���ɡ�P{��ǡj����� @�����#�^���`���+����N%�©�����J�̹Q�/?��&Y	��OE�b��g�D�[�N�X]8���<Ef5�8.㩆<P>s� ����qvjg_�He�oSCb�����N��rv�U����-��=�wm)�~܋�'g��^[�ȹ������3]ݢJq/RITȱ����Z���cgu��d��7wzܴ�S����<�1T���<��7��UO~���<�H�ٖV���z�^z�1q��f������ΰT��a*���{��Y#q������)ߎ�NNÝ	��ߟ�t�ݎ�.��?����1�M�Ԉ���U���bh]�?v�x�\ �߀@�֠ W�Y��O�[���&��n/Sa ,H��`�'�:��5�CC���k#E�!%}�3s�.��0�� �������y?7`��U��,�?ۈ���ٳ8��n �������	�nV��օ�Su�AyPX��������ԛ�s�6G��)lE�;1�*QBʋ�nf%���C>R�����RÒOXE��a��:�W�k��V/Y^��.q޼>ې��ľ�L�3m�Q:4���P*J��߅o6�G�nbS��b��i��[F��V+5-�ui����L��07r�c�Klv��9��m��,�aw�Ku}����^ލ��)�ָ�;�V<��p�תg��{��}�S3�g�Y=�a�'��gɶ�����E�e/:�F����VJ���Hk�"�\���"���� ��=������3������#���u�p�`vZ��W��kׂs����F����{�\Z���:��p���yx�F%��K]�0��d�/��Q2bm;ܤa�	���>��F�%ס���
�΁�� ��آM�4y�A�:VSS��Q����T��ؽյպ
Ov\�Փ"������1�й��f>������[[œ�X6�6٢�<)� 6"�3�ٴ?�����V�f�89�Au�����F��zY�XXۋ94�B˗w�P��ce%�4l�xF���iJ�<h��to9^#��<����ہ�W94�e��>"�Ct�3>�B�J�I��H/�}	$�DJv�������L��=vsw�K��][d������s[bW���N���ﵽ�#������7%%%�#�3Vlll3
�����F��*۱�UvH��*i�GX���y����YI��dQ�bKi
�$�*l/����>�	�$%'g�����v��PPP��nmn�(
�y[P�UZVf��I����b2��u��l�vs��c��D�do?�b��>4��~r�@�=�m��`Ŵ0Xȵ��:���+�g��t��Hi����ZI��_U(�ͫΠ�I{l`MkT��f&�K��R]SW�P4�]]M�c,s;5">�k��:VCŉ-HM���ͭ����������˹/�_r��.���ׁa\\\t=�c��<�q��H*G3�p���]�I`p���@$�n�R�6�mm�|�a��`�ޞ�o��a�f�	���a�u��h}{{P����/_>h�no��	*$�����y�A���n
B�wn}��͢��6*2��I��kT�]�%U�f�ʫ͹�.��r����m��X�}��oii��֖T:~�ߧ�>�JHN^�Rd�ET0��n*+g�u���,SNE���V��k�\{��0]�T66>V�έ\�Bn���j�5�B����F[��ttĤ��j�
xk��TR����]�������Ru���Z-�M���G�ٙ�v�����������.��T�OI�X��䑍��d��==9"����~V�����7x'I�/SS���j�6��	���ώ5�NN�}����d�;z�/22rfbP�z���"�血�lh��s�5+��Rpcƹ��"����P��0�e����;E
��݂�|��W���E�_KJ��\�����Q�����(+)��1��}29&&H�=���p�m?��ji=��OW���>_�#����,[%Y��s���;��������`�P�9i3�r+�lst��Y���iQ�����۞{$��yk~��jc�:��\�H?(((,9��b���{�ވ�4��:�MGw��k��B&Ǆ��~�l}��MW�(4�#�g^R)����rH�js�7��C�;�a�U��[��wChiҤ��KJo���yQ�P��s��ːk���`�/�\UWd�%K#��%�d�7�r*���e
������b�|���3��+�1���s-ѳ_�$	���6�:׻�(��;:M�̰ !%%���OHD/қ�ceeU�y���68�9�&r@.��(`7�f�St-qm��P��C$}�`-DAQ�Ǐ緺��҇������_���<m����Ž���A��=rf6AJ`�z�"�0@qy��5��~,���{���*�(�`�JTG>S�yb�jd(9f�uq99y��X!`����k�d��Pݾ��vUUUյ|gF	�? h�����4�*����Oc�dVj��2��T]��㕍�_f���J+���'=ۚQ��oZX��>���ʲ�#�����kn�^��k��4������bb��6�Th���׋Dmpqq�R�ӧ��8Ptp�E�E�1 �r��p:��TM���Ƽ�����Ҡ�rd[G׷tY�j�c��
��K��z��˫�v�"c���0��I��r�)j��j+�M}�w٪)L����5{��f���Sb>!�W/��5EtM���YRb$�{wc���lw���.yP��5����؛�Ò�*Q=�a 0�����:��w�[ӚN�n�	��ح��?@p$�R
j	"/�����>����q7k��b(��ĢW�.G�S�a95�����(�~Ǽ`1��ᑰ�;�����5��`�4DMf>|ٕl�i�-4�a|r�R�LY��yX�����mÀ���,J��\---��۔'�u1}<
�,Wt��:xȆ��6D���"u����W$�t괣�d��tx��D7�om�k_ƐjbK�����w�^�����$'%�)�b����"䧯$㰍��]OOG� 2�I�7�^]"�쩋$�!N������Q�z/�#BG��?&�f�ڞ�ђk���	g�8��������]���Ha�p�Bg�0�F�xكB%�oCy: P�3Y����ï&P<1#\~˗72c���i3��I�(�q����
G
��
KD����*�A��)��SJy�b,OibXz�ށ[��ì5Jk33�b�����8ͧ�'�+'�����!	��^��9J���%�#�C04���h}�L��0��I��!�E�Ѵ++�ʤF��^�~=���L#0����1�V�mަz(�4
@[�C+���p�Jܧ��E�߿_��9/��B8\�4�J���`ꗮSs_�)2nu��d6X٠�L��p�1WIyr����G�7R�F���#��k#��ce
rwn)���y����Qo��c4�a��8��m����&����v�����6 ��T��Ag�G���w�0��^�x�m���&%������ʹ�ϵwI�#�^��][�,�Z|� �` D V/�}����@�k����K<�v��j�ni��W�z"K;f�?^�<Ν�n��
C���'''��-����]�>�}{�z��if^��حَ蟥�
�{7�̻^���I�R�2��,�/�T\Q�R����U�	��Tii�}��2*x����4��m�j,� �6X	�C��tT�S�qZ�n�峊�,)/oFt%<�l)9����A��-|���yxx��߂^��5k��}�I�w��/"��f��H���L��B������,ʱ9�["$!v�	�߹�ZL���0-u'�C��[o(�=��4�����_���S��[�3:=M��=�_Uh�pO4`���1?:z�n��5��Z����Vo/\?i�S'����NG���)�p�?ڞWwws{�^��X���뻷��BL�����7��*�L���Co��7�D1��!�'eK�-�ifk	��DWٙ��$�l��D�D����y��8�6 I�J���W���;�CR���y�� [�M�ȔC�J��)y]�_�S�����B��~�`�_@�7'�Jx�v����-�r��5f���֣j������~�f��t�ƍ�����G����I�:�}�A�m�^ ���o
ر����4�˄�gb����xw�*e��ѡQ�|�<��}r���l3�I����T'AR�srr�6vs�¬'�^B��c8�F����mmא���و��T+�'�3k���@7V�� 6��&�T]���"��17�ů���y���0�r�y�:\����tr�A����,���x�V��{�Vxd)�!����3�tK<:RVEEE������r�Y&,���ǘƓ��7���=WL�~�%R��'7�[f�HGb� n�����L1��eIDKP��Fv��"$$��|����%M���3������K�Z�_D����k���>;A 6��Ll��2�|+�|<Ip�p���<�^��9�h�%��_\�eTM.H���N�w��$���[p!8��������]��{�7k��:	�i���#U�ϖ?�;��|m���fW���D~�~�***j�FL�g`��rw5;@ŷly���-�Y�a8ג8\�����HX��n��\7��K��78�H���H�W/�ￗ�Rq 0O&&:	z�#��GV±w\2�=���W �ޓhg���;�o?�@���>^��g�t>�nܲ�E:�'�J���V�Բ̓ɚG�_T��J���3ƭJ�����S��IBB(�]�׃~�R���<���X [�XIf��I���`�ciU_=a����+%��ABBڑBJ���\?O���������Fe�e�'�4�|���}W`hq��fKӕ�*�R� ��Q�EPů�_P2��=t����B��>Pw4qwk:��'Q�ݻ�^�\�b��W�ԯ��5��7ǥY���p!4:��U��.@��8YSb�MU��D�r'�{�uL|�T��ؿV����n��'w��Q���6|S�/��xピ�+������M@7;Z��%qZb�K�e��sˡ*����h>�����%�	ei�"r�ͥ�]m��|�=5�|�V*�p:��\V
��x�ʧ/�ru?)98�9����Mr� [z�5zp�������h���,x����[{j8&�w��� ���tz�L��/Q����X�2�l6�0�C�?�QDDFV	
��>�."a ��`�����2Pm8u�ll���kX4�k-���;6�pA0�C���(�Q��K�KK#�h�nе����!�_�k�bA��� ��O�[���b�=p��G��fm6�G8��9����	�~�	Ѿ�k�G�м�^_wg��ys�t:^r��kr� 	�¶�i��ϯt�%-��R�~]�MV��xuON�a	*,�T���|�ϲ�^gAF�t"���y�_�Oy�L����X�Pl�+k�����~W�ԟv��*D������uM���P��K�75�)B����:���.����^�Xkv�ŭ�
�v�hs9_�s$���F��پ�\�)��K*�g݇�o���.�na�"xz� B�=C޿��iƥ��)������C.�h��d�X��x��J^����aN� ��E&V���Ɍ5��Ӿ'/��	�}X��?���,G�m�����:�� �O�T6���_�j�2R���FXJF�D ,:E����A	K�e�n�"G�.Z(�Z�k �Ob�W����K��IW�Wu%@QY��I���)BMP�B��qu//����O��s����G^Y�&i��U���0!��g����5�&ʀP�H�c��_U;E���+�M���'����W;\/+t�tX����� ��y���vQF���B��n�/�;���Sz�&�Ro��jR����Q]��v�xv%�s�H���d�D���*��Ko�k��P�$��EdI	�~��^����*���aI/��ƚ�Bur���#W#�[���w�8���T-~"����������:Ý�����x�T��G���{1>x�s�p[[RR��(�U��N�;��I|{C���'�%��ѓ�)�����kɧ->�=
C��`:ŋ�hDçx�,l�nL��'�fNo�!V�L�l���[�������O�j;d'ҕ^��a`a�1�S�[�㲘���_pLv(0�����)���ƫ�$2�eetu6���h�Q|����MMZ�+���z:>A4��TMn
JbK_}��V�(��$�N�R��P�rf�SG7����F�EP0z�s��\���LI�R����)]#W�T~Ǝj���ϭաyH%�+Է) �����}
u;������/��V$OV�ܫ�	���1W�p�)��D�2I�l,,��٤I7k� (�g�ʬ�!�2���w�:=�\&���VQY�N�ub�FQG'
��Һ��Gzr�RS�|U��4)9�+��g.F�h��5z�wl��5~>����u{�1��&�ybNYE���}:bb���L�jk���'MMM�����KK��}M@	���+})��j�^����1����U��]=���T�dBU	����?�⇒b���|u%��(yt(����x���6��z�Ma���+C���r��)(��=cZ))�Z�a܌���m��uC�)�k�������^AYYYb�0�lj�:��E��u[�����b���Ay�޳���u�wnÌoA@��Щ��'z����NSKK�k�z靪�Z��@t�y������2O�AΌ���,�ro/�c��:�C���R�p�>k�+�֟KKK��ҳje����) ��,��~!n�rH컳��\O��19)b��&���f�,������1~D>2>Kr^i��r/i{k+kڼkvC�k�T=^�k�1��Υ�N$ӯA���Xɼ_��Y�ba��j=sNk�4$�'U4U55��������&���P�F����n77�	�!~� �~�GU0�����{z�M�qS8i� O'�c�Wy��n������ݷw86���'5V����.?�^��#�¯������k�
�-a�������c#���X�d��s8��[d����!���u ���O[�
�7�����a|����<I�|zV��ֻ�!f$��:G<�Hwbvf��9�����?� �dÿuu��cM�A�ؘAm>�Y�i�����nb�qѮ$��H�\�٤6�Q�55U6g\�b�������OO����������x/Ӭ��6���ĠW�8~�x�2\q�=�s����s�X҄m��/�l��\ꉓWR
L:�9}�c�;{|F���7�h�
���1�n��W�n�l
>��S�;`Q`U9����E��6��v3|䴴FcE��Y+C����{�GH�}R��/R
��R�4|A����g�?[�3dԌ������X\���U��=P�n7�9����.;{��칐V000����GGg�(�7�RZ�yט�;��������7r�1��ιX����]������l������ٱ��~�&���!�z����4��q����
[�<���~�b�z��+n#+���8��v�$��ա'ޑ���(�T�A��A��9bU��bb��筺�����[��\�4�$e�s� ��˳¶Xٶ�;uX��0ɴ�v��]O����|R��ìu�G!���x$�z������Z\΍�l�4c�_ǡ����4=�ɜooJ��W-�?[�ݵiƟx|�v�<�^{ 9�������O��w��o�����%1��}�>���k���kJ�knoX��)l�a�2�(K���#�N�f2��;l:�����~��_�0�+�A3j�W�+i�D^��h��r�b$̰S&2��K��'v"9�fE�ٿ=;��4I�j�L��e�H�R���x����.��᮰"��<�ߧ�^��p^���Y�j1:"b��㔓�3�ɺ�_,��}��5TT�i��zVV�ӛ�\S��mO�a}���������B����ݫK�r

��c�Z��V����e��A[���GȊ*��~�LL<RAG������:f��@�T9��-�+l�)�PWǝ/�G<Y(Q�E��C �Mn\417pkp �E �!��/ԕ�V9�I�-tDGF"����	Y~����.�
;�K����{��M�D�(��y��XUD��������(�j(N�nҊ��ve$�"���D�o�8�;��D�T�孭�W��@��mI�`������Q .��������H.;5V�/�t���e����꺌��������������n�=�K5T{��V�}������E,�;m�=:^dP�6v
t�=o�\��+��}F�� ij���wZ
�V�h8�^�~Yv6)�ns�T���/��&+�y2�%$P����F\=u���Zl���)i2+�xh�-��w�i��a�|{���+Qg+�5)�k==�B�^�i�v

h�ڕr4nP��P�\�
6FV��y���Tь��J�F��i��z�Y`�mU���7�
z��a0&

蝁��Gw�C4@��{i��`u�|�
Wg������r�o��U{I߰�~�/�U�s��V�['�8)���Y��dS�#h^%�Z����%�)Z��V�*����;wX�o��( �<Q�*u���Ѭ���;�o�l�vv����W�#�+����ڥ�*�|go$Qr`����e'���N���H4�y��z,�$vHNMm�LKt#c��eg�|z�\S�)���@������.��lzJ��Êxqy:**�؝�,a�C��Z���-���T��1���C��P+�,��£��q��j�гB���������⪜�M6`_�'�v�Ԅ!:���A����+�3��q�-X:�[�ǧ]I�Y��=�@Zw �79��!���۫�l�x8�* ���s���h�&,^�l|=�ջ�#�����3}HߦdN�奭�,�)<^72znSn��żg]~o/u��d  �J�1���I�������[NC�ة�/�i^�QX٤S�wP�g6�5!*v��1X0F�a��<�����@HZm��[.����V*~bƧ4%&�]���4����iV�'�Lw�<@�E����i�Ra���9;��$�v�w�V�S�_�GJ��ګ��Z�<Y�|�F�7!�93�PsL�u[i�o��/̤Bd�2ҌF�z��F�Ύ��{��Ġ�#�Cǡ�n�&���MC,R�l)���2ˑ���8���qj�z~�T���kp9b����AB$P�x��R�$6u��|��R��i�����>���)��oV�֨8�lHj�N����4�2���2����B����V�Ro�6HF)�==>�dll��Ʒ{[�x8ׂ-�d����P�<V��u��]t�BO��������5���q`}���N��z&�~qeeg��/ZQK��FFFFp,y����Aj�GR������9���{����h`�rs��x��� ^��&���ΦT���-(/T�Z� hl�4m,))�#`T�0������ͦ�~� �XDС� ���L?����$�FAAA�ɉ������Mt�h��V���c�o}}o�V"��O�q��瘘XU6�}��*���&бs1�����X�i``�Ob[>���R���x�i�t�>K0�-���ި
��#��bL�7aa��G�eD��>��Vf۽��'\.��-U+�_9�P6��\m���R�O.zf�DP� P#s��Z��5i���,�m(��u��Ƶ�M+��;�:+����� ���n�#�FXR��`v�ѻ��R{o�8������k#,liC��89�Ҕ|�T�ݸܛ��9,���+_nc��'e��TW?�䛹�R ,$�gQ����T�b��j<ssݿڈ��㽳ϖ��FW(t͟ǚD~�Dj�~,[v�{m����ے���?[��ƠdY��rYU2/�#ϪL�3Ì�&�`Ʃ�w�!�깕�ؘo�.ZYC�#���A�ӳU�k��`g2K�Uஉ��kq�����r���bV�0����j���q�Rᷯ�0�LBFxX�<�rZ��=3g�)�/��$ ��YX ��mK	�t#���lV�":H��"KJ ;�ZZFfk&����h�g��92})7���o���|8UC�~{��1N3��[�jI��z���<�%�t�YnkI� H�s�S�(�]zG�!���	�����x��5��L�f̜��B9�4�3�%+�v�x�D`�~5����LAs��oUIRq��y8̲dc�0\��Ɛ�I�o��h� ��,�)/��7��SY)WR	�����hݫ�� ?>��������.d�7�'02��~��̿�O>��bO�6�����Ұn(S���|1h�f�c��������9��Q
"q8��p�ɹXk)P��KdН�:��*��'PHD9���iQ����l��%�Flpx�ǐ.�9��	IH@����}p8���� Q��l���7t���'��_�����V�bR�)1��n�����9��;��F����L<���`/�߅�|�)G����==��~��bQ2��"�1��)�y~p��UD�,��}5;�Q����ڍ����-��ے�4�P
m=G�x��%�����x���Ƿ�x�&ZMAhG�ZJJ�R��`�2R}�e���ښb��\��;��5�{QQQI����o:�ߌ�bj�������)9�C5����͠����;Z��� ��>�&�<K�G̕X�v��0~��� �������[*c�^HpAW��46�Z5Z135���������u�)_]:*��⮜�3;;���y��ަ;7�lwQ"��i��ʬ����O7�5�,��Yt����Ӿ��?<~�\D�vAt����U����1�.q`�,X��/��v5�T�t�P.�I6��Z��h�N}U9�4ٷOb̦��,���ӟ0���q������uS!e���zm�K�7�PF�}�2Rz�Ł��U��:��x�����Ԡ�:r9u��B��^��V\��n쌧qvƐ�W�͘D��b�}��ڿ���=����%X��digV�IX�d�v��ヴ! X�,>xx	ñ鄶�^@��?��������}��_�>Kn���P�PB�S���b��A�j��a�n�q-,�Н0u��Ê�ɱ���}��Įg�F�⢚��Ѧ�+�(�?q�t��'��=�e0D((�$v[��� �e��ǻ?x|�	\�WW��bs���D���b�����x���� ���p�wFy�{(@��- eg=&��%���%�[�����!C�1���sI͋��'@�S�$�WQ��7���}
�p&���8��y]���N���N!�[K1�����|�P�s��`O�NT#i#�;TLi���G��@�4��e��QgS&��j�!���7�������B~��i��J(�U#ft���"=Y(S,��eqAHa�̗�P���;U�a2�e_�Y!�KL�$#����F��`�+Á?5"C�fw�m/�S'��1FG_Q��赛s/S��d���2�1Aʫ�	�?�
�EP3ddR������Ŋ��B���t�rgMa!(em��X�P��L�(�	L�Pl[A�tx��|g~{��Jp=^ŭ����х�l�AE���:��%C�p�q��e�
��%��|��
J�4撄H���F��*�4��?�<±��O����gzv��\	6ϊ�5-�_T�����ef�����.W �H�����V��bab�O��O�ɡ��$q����ѱ�w�_�>9ju��)������������abBmq=�v�=\�+�����n[��ļ���4��;�l��x	��� @���Ȁ�t��g�"�Ҿu�uw�I��,M�PS���:���$�N�������p�͙�`�P�P/��P˅��'����uҷ޾���+�yqRy
|N�hscc�ϨYO� s��Yz#!��M�� �ٿ��Ijk�����)�t��܀�C��d�u��M�%�\� i��͞O08��g@���^���v=p������sFV�9?��XX��;�Ȱss�qѴ�Y� !H���6��lV���6�Q�O7����!�L0M�Sv2��01�4)#��~0f��X���,�2��Fs$oǛ��j��h2w�/�����3t���mC��{��|W��A�~�"��e�ԟ�D�"�kI\�xVf��0���Ԛ>W3����G|RUUMϛ�oWBi{Ӛ�426���3�ȸ�_m����*z�1;8��/p�?�����7R�E��29,Н�VU1q=?��Å�`�C����䶱��	�f�W�`Q���?�:m��)(����Έi�������%�^~(�CO͋��xJF�K��������� x�W��p��H����A';n\s��E��a�$Bʽ����6x�����2|f Cp鵳�mg~�^8A/;�p�WVUMg�3�����E�W�C[*�0���{k�s�ӷ~upP��B�L��׻%��LfZE�?n�a)I�ˇ��/��-��WdǸ�+.�S  �3}g�}��� �ˠ�ڹ<gi6�.#-��N�tR��(dZ��T��: mS'����]8U��-���ƉDđ	jA
x�̸�>9h�#��O��V:@!E���K�%6����?(J�I�4i(B�v%|���R���ǁ�����su�����l�����~w����)�����
����ƻ��\�4�/���,�^�ߍ�/)�à��67�PX�B3:��wZ �bg����ҵ����~�%���D�k-�S��%�֥eeS�c����z�W�f�`�����!�ɮ޽�ڥe"��HG�O�#��%�b�Xo�:9_k���	_6}1�NIK	�; ��z~�hNx6iE9[�wWɓ-��m� �b�5{���I��+>yr��j/�����v!���lPKf�ϗ�r��F�qߙ�'�v^�nq��d\���[2�� +��E�c����V�}�]O��c��;)��+`%��dZ4X�b�����w�M����F�OJ�l���fc���������VH\\�֡Ȭ?�0�"��<@�%�1���`�#��񝿨�	R~�K¸�����!�#ot�U�t�P��P�J�<9C��= ��~�d���p����H��۰���Y��<�%==��������;�x��@�iE��2�S�4�'����w�&hf����&�u�@���J�V��7T���#2֒p�7��bP��X��t���L����˟�8Mv�U���h �}�C��V6�t��m����%�h=���T�|�f
�����z����-��`BT4�޹Q���CL�nB�>B�����6��з�`�﷋�>��ӥT��N��u�DbG'�?���TF�rm���/�@�A���.0���_2�$;�S0`־����m,�M(���Z�n�~�ll��\P�m�TF�N��$?��=(*H�嫪|�[�aN�c�l�����5F����Ia�3�(Ϊ�&���֖�l��ù�p���}��iBm��i�訨��[��I�K[��B���D���A	6�6{�ߜ�c����!;�_Vv���$N��Q�_.r0L�(n^n���=1�{ѥD��P��Eāzv��9%J:��Y\||��\�s�Yr0���D7�Xt:�  X�V��i������X��7��^%�ט������|��k@U�jU�3'G(�ZYE L'��b]6P��z����RHy�?�6x�%i���)��03���x�q�~�����;�"Y���2�("|�ڨw5�������o̒R����CZ2rH���`�u$H��a��⓲÷V�����vp��2�?���4�Rr���E���+��F���7ce�1�*7���L�g1rx6-�L�̸=�Ȩ=Mf�W�s�� �����U�lˊ!�W���Ka�YZ4V��n��#uHy�=�
)��Q����}V��[{�C�!�-�h�h�(�g���6��J��^����[������Gbk7;�K�ث�_P(��E�h��m	���+,H�e<����S�4�$��`N��7��-)�_��**�-0�n/I����X��ÉV�щJ�z�;��)���y������/�ܼ��3�-�����z]x}y�����z��m�$�G�����װ�+�~���b�	��`��?±�333%�qg`hHe�_�T5:��~�ŗ�e.qqqP�k�}1�@4q�3�1�{vhV	�Dv%e��<���JK7���,��D6{�vj�v�auǰ4TVPRʕ[*���>\` |�:�{���cwu�5-b�����amC�xx��TA\�?k��5��ǣL�}�>_;��Ƴ��O�~Z��er����d|��4[�;�_�b�v����NKM��(F�·;'�|������ocUV�, `�{D���u/,�:�=���������D�lll�f�ڲ�mu�eA���|#�����I��IU *$p,�a*#s�		Id���?���Ԅ�F�5M��Jm�����B��F�o�U�4y�q�i��-�M)RJ��iL�h��>2�&��bP����W��I���+C�<�ZUGxGZ�v�(Bqr3+x��-�NL,h��7�H�,��Q���"4$$7R}��f=��3��Hm�WmV܄n%X��3��?(ir�U��MLȫ��q�e'��c���=;WVWg�Fg0QQQ�z=D�p �w!X__����4�o��Iw�g�i윎'( ��[��Hy%���HI�I�
 ��y�S:�t��	``���e�c� �_|?3�Ɔ��ff�A����m����%[*�t㻌���k0#F�"�S�!!�ʞA��;�s%�C�^+.ߝ�enVZd�W;2$�$3�� O%�!�hO+׷#7ϰ���A��7:�p7� ��_���O����P��4*���ibf��zO��|h|�P��6k�{h��#���]��i�rxA{Px�m�[奐�Mppq������}�N�E�� vZ�s�J�m�{�V+�f2V��{��v~\�t��7���������6��>��_��|�����_�t2��i��5���bc�~I�:�MH�xDK���SWE�����B_��O����*lmM���D�='H�9>�D�O�Wdn�<�h���`�!�o1��N��S���������b����o���I�J2�h5��ޡ�8�?^wǘQ�����V���&&�k(��<rB�֠�6�ҳ_`�c�suA���h^^.���� �D��ee�'�����D��#�o<��Z�dD���rs�z���4&��Zq93���1ع��׾|7=���ņ��J�a<`�/ooAkbZY�>q'��c~�AW�j��-���~~����Z'g��(@���5(Q�������J分�^�8��dUX���N�C�
O������E�Ґ�k��$C"����7��Ȼ$�q|I��JFZ`������G�Yud7����ż=�Y�z���3����F:W����^P,��cR��O�!5�"`(^�<b�S��O/�+�P�ʿ��$���Ml��l�5Rt�0�6V�q��G��Pҩ<?����ë�ϸ��7W���A�붔OVn
I#�����Y(�e__]�Q�P2����B��Y.�o���]�94���v"u�=!��v����2F�>�Z�D��ϳ�x@&���`�[��� �����#�[j���_�w��S9wÍkMM,��m��ҫ͢�_Ӏ���2����pku�X�-`N0�w��j-.t���둸�X�\���s޽��;x�} Za�S&p?�x�/O/]��!
�;��AE�;�L&�8��Ulm���#�N��V(� ��ହ����`V6��(����g���|�%8ʛp��B�HVZ��t�Z��En-`;��H��ϥ���z{�ϝ���B�c��}�9`M���C�D(�kjlԛ�ոk0��逸���	��X����q�ݰ�p-C�������OU���ip�x���3�C��[�+>!&��MP`���ծgo�Y���P���������'���I������%�i��@�"E������*�*M�F�xu0�\�P��Å�N@�PRJ���������oT2�l���Z�+��cM	�q������~���s�
QoV����sv�{tOĢ�����O��z^��E�.��mvZz��YD�������5�����Ճ��&� �FN�w������U���&e�! �$�3'�b���G�x�?ӷ2�������Z��
ҝ���4N'�i�Ѧ��'�s%*[�A8�KK$�׮>�~A��Ԙ���+�M�VG���~���$,����_/)�E~7 j���X(��	�FV�D�s놡=3n�B7c�WH���� a�i�t�l�s��]���5%��f
���P`&�đ^=�ϕ,q��˸�2՚M��c�
#�\�Ent�(�rj@�
�	#��i���ONP�I�::1qt 4��_�,��4H�4ם8}���{��ug��b���Hd�F��ch��Ya�씫^�OB������`�JL,;�&�{*�������R����⻦�y:ML����N����yC<�^����Uzk���K������v���C�oA]$����i���\anS�4&�@��9�L�(�����4�H��Fu��4��f&����.�D��.-/���ΐ��N�v��i��v.��?�$K�6X�o E&��^�=+��5����(wڔd�
R̛��Zw���>L�wO��
-A&���0iؿ��k��*��������K����'5����S�<"+qD����P6Z�V�E��i���w=ގ1U�u����D�6Q�X
& T���sЊ��!*��XR�9]�7�c����xo�v�'Me�-��ߡ�)`eE�4����k��hvoRקkb#�#٠
�*"�GJ���־Z{�p���������l��H8����,X�v@�� ��L��vg�_|s���$�(at�2y����<K��i~|\\���!�\��0�|\	���G�Ʃx����Ϗ���|]����K9������y&�y��a�_��%)!���/[�o���}�X5en�!�?��d�.��+}x#A��a������-`��p>��~z2{�=_Ӵ�p���eV�z�����'�4��cϚ��&G�9�ҿ�W�+��&uDX�X*Ŋaoo��}R��L�!&%E2�cmumk�5�O�4RUA�x̚�`�N��,@(�Ll#�}���¨����t��}��q�0��k(J��M����*��(�J��ST$~��z���"#���/���� �:.�_g���]�۳�G�_�#ō�����V��v�37�V[\u���R|I��x�7G� �zy������J`P�(�q�{(�v������ *&"����㌸
������y�9̷j���F'<�g����󥅥e��M�^SSS�j�o�)p��,RB�Z4	����9	������ZY�ى�|o������$�0a;\��~_��*
<<|Н��1hR���e�`��LO��R� �)��2����$�
~�Q�7בpr��ۮIj�Z[G&���̀���m	��n�27��Q�ئh�U���D� �����zT'�d7�����������u�؂��^�^$44����%^xxx��oϥ�?�~p��������tߣVy���t�$BA���7h{�j#a���b����(�ǯ2�)�JR�\m�"c��D6������X���II
5騵���F7��VaJ���Ϡmt�Sя�.b�D�b��^��m�%c��c7�W�T�a���#����	���=و�޹L�VHS�$� ��n�5�~���bO������'U���ǏU�q�~�|^/�$1�0��i$v��9L��P�� ���by�R[X��I(a�P�D}0���b�=�\��ک�-�,Q�S�c��+����YL(�:� �n	�;d��I+�x_�Db����ޖ�5����%�e�&�-�������(A���~���E(R*V�X2r�b� G���f�]_�"Ɛ4�Y�`�i�{� ���Ytfj$>eD���dV��j��?�����8�,�s��@x�&/�K	`/_� ��g�����	m#�l�C\�����i���pNy&��;�u�qddd�O/�脦?3s�ǂM=d^SS��ȅL�@�Q�	��E��;Z���vOz?4!�8nnn��L��-���c����lzЮR�Ե�:P�چ���ׯ_7'�|�5"\���6^�:Hz�S{�խ�@e�#�����i���
����k���$B��?,�������绫�L����L��O�8��*e��x�6�O���5J v���)ԏ������� ��tP�Y��˽�]�r)�A!���;�����6굍�	��:�"	�FV���2���
8�a�oyL*�O�e4/��X�:;�r��X:��� &Á�uN�o�B_Ѷfd�R��y=~#���̫���ݯr����H�y
��K�>o���8�C�����"R��V7F��N%���0����kڡ��*����@��9?f�͖k��^�\h�k���_�\�r�]k􆀾�P=I9��~�KUa�H�đ���6<q�6 ��.��#T��E�K�$�&1���h*��~�Z�j�sJzz�_�h��1�K5v�16FF�.g�Y�鏷5ů'�e�


f5�����o�.Ï-{i�B7ЃnYo�����t"�9���F�a9	��E�m	W���]�P3��^p());�@���8�-�\	j�b����Ҡ��[�ƍ=��eVK���O�'�9jR���̐����nz�qq�Z}��O�:Vˍ���l�o� (((T^x<�iTV?���:6� g**<���y�𽷷wi�v+x�:�,2��oO��_]�_�x���r,�#��ׅ����q��;"E�Ņ�d,)�D��X��!�H
�-`�8�thB�E���^1��w*|H<p<U�H4�о�du#��p2_��dff
��8�M�����[�Bց 9�0	i��S��?���Oj�k7�c���_&�	��ii T�b:.7�ıP�D��Ѣv���u/����x)����233����9�-V���VK �	Ē���4��6YǾ�<+����{�Vy)E��u	��`�SVSU�u��b��⊱�w��"�+�M��|`Y��\���G,b9�,L�������!!0�w�`uF�O���6K��*�^�k����[d�1�߷G��O���H����I���� t�k-��7�99ճ��EDŶ@K���\�ǁ���jLZ���k��<� ����׿�TS@ɠ�& Fͳ5=3cwv�*ޒ[�g�����g�2J7��N�qӳ_�o���s��=nk+��kKKK�ښ���SPP��mv**uӉ��¥'������b��a�����W�=��:=�M��~W1�LM�Ġ��r��b�d�e�)g���l��g���ޫ�å�=����C�[�@�Md@QQQ�sHXD����lO��׷ʳD]5YU99��>�J�;j JY	��OR��dC�?_� ���{������t�ڽ������'.�7!���Û���5�qpG������^*C35]��u��Q�{��4e���S)�U�{8(�܇h����nk��A�q����Ƞ����282b�V����8PArC6�y
� ������t_�'�gfN��p����5�#��%�b
	�Q�9�7�w�@ض����abam��yD,|��G��5Em�����D�����L�Z.��~:�n�;n�ͅ�ut��xKikx��'���%y�S��������΀^���z���h"2u��|��I�i����9�����y��~��(%���=��ޅU��\@F�"��uԛI���e/	`d�.���
,W���cRE�U!�!A}Q<R9|��*}|z�j^�����Z���i�f� �G.=��j�DEECBI�X�_Ԩ�2���H~t���uhBhjr#�KqZO�s��JĚu����<��V��:�ߣ��p��)��^a@`��&f_R9��Ǵ�PPP�n���M!�{� ������bc�e3���M���F�ߧmO�I�越(��iZ.�N숏����ĔH�M�7~�%���vA�`e�9���A��Z���N�A���;��w�Y�:�y4��r C�5u�ir�Z(s�?���Xf�-k/P�H�!`��B����o����F$��6 �«��A�P:�i��^���I��c��^z ��
�:�2dK����=���1�����u��z�T�.lWyw��+a �*M��Fu3*�ML~OV��!�1�p]�.�|]���.�p$ί_�6��f5��oG�H~SW��+�����d*���z�Ua�lS�>�Air\s��J�)[���u�\)��t�����K,�T&���}}}���c�k��acc�o]��^����feQ�6�8j��+\��-�C\[������-�w&P2�++��{�ޯ[Б�s�yɎ,�^B::D&���kh�!M �#���5=0)�m����k�#ז���/��3��W�軃1p�+�m/��Z/`�y�2)
���T��J�6�{��ҿRT��2��T����~Mq4`Mɗ7��E
���GT*�-�N�r-��lZ1����dlⲟ��v�����V��N�N?'s'��gkΫ<��,r��'#�MH��S(�	,�d/�h�X���_mv���*r,HX��%&�v��
��CM_O�~6��8¼�S���2��N�:>�ݕ~<���)$��tJ��⺊�@e%%��h��C�mF̸��W\�55'"�����rv6��@�h	��./d��g�ePqp
�mn��yCoo�F�M�q�p)T-}�&���w�S"#�"�ԸE��04̭���B�p�s�jr����},Kݞ��U���i�+V��JC�:칀��V�қ� "R9�3�KxȠdcS,=���̯CgDDD�(�Y����/��*6D�P_n�x�2��=)5���h���ӈ� x߫O��5?.��l=�L,<�U�K�@d:�C:VYd�b����N4:�r�l�I��+�5��p	��>����v��;m;;F�=�X�����=ӭ#thD"�����%�^��׀��z&5m�kp�(@���������\Yo}�0�þREW����?�L̥E��3dgCz0~����ЂY�O%EHH8g2V�Ֆ�j�x|ȉ��Q�x}��u)�H�����1~vǗ����:�?-f�����IϪ_���
��R��mp���˷f6}�WU�؉�R��{�,�خK69������[�utm�X(� ---� ���tww}��.锔�����3���������s�o��{f�Z뺮=3k4�Ԑ�����L����[�ۖ
/��%K�p���E�r?)�bgՁg�}���a@E��%s|��&:�pjMM��[<8���9O�6K�W:7G�c��CC�n�-��7�G���Y�Y�}�W�Rm3/��Y�6��'�G��1�Ijp�p?�N9��M��3c�=����h]���_�>���l�wMUe��&�D�/�X��X�Q9F=Z��q�ϥ���ñ=Y<�0���'�V��vcR��kh�#��@���Q����N�"&�Р�A�2.)�������k���;������e^��D�AɎ`�QQ��Ml�Jѯ:Ǎ�(Ĝ���O�-<�/�e�B�-������1�k{�S
�]o�q�<M�ԉfM��A�RUPppA0�����#�����F~$qQQQ��t��vn�����q�~��c�Ñ���U4�OG䲦�z�����D�xrr���3�˝1��1Ƥ����L"��z��k�@�h�`�#����y����ovn���ک;*���=e-����௶�MY�q<��^��5>�E���ps���t�� Z�L�����V�ŧ��_1��3	����Ku��#˫��0�q�:�`�_��6G�j�N�*�ግ�3)N�%%J��D`�s.�s��������l&�����tn�L*��(��o�fi���9p��8��+l_��
�P�s��q*��N���@X"��9�b$4�`���&0������E^느�Y���?`b��T��<+�#�7%!SuT0��^�5�R��k�\���j b1���Ƣ�;�9�YWEss3�4�CDX�B~��Qn����P������O3�;I�rL�F$��P[t��Di:T�V�ؠρ�>�FK���S�0�qyMMMd|^%�`���t;]�t��&G���Yb����Z� #���F�M7������m7�h� l�n3j�(cZ���
���m������\����2�B�������ne��ʦ�(ӫ"� �@��ۧ)����+A  %_i����r��ű��e�tߗ�13�@"��Ӄ���>o����wr�M�-66�͖ԦzkqWO� s�C⻼�	�E�t2��p�5�-�Eg�CX���Qt�s�Uz�Ś5v��e�p�4�kpY��fg�p��H1�JMM��d���HZ�~ё� �놬����ET��Q{�'+)*���C�γb��f�dyqy�`)x;Ϋw^���AǜAB?�3BB�ƻ~���s�<0�kt$�{��R9m�{�"��ND%�!�K檱S.,�yޞdշ=&!�������^i�_�z�L���@��/ND/\�X3�G+e�WWW��p8,EB�BQ�V�u�mq��S|�
�o,I���ӭ�Z��i[[[���3��U��h�3����ѵ�=&�Z�
h�􊪨�M;���T��ex)�]��	-
���|*�����M��|�μ�9��(�I��A�c�<c��Q���R[+^
�xdơ�w��S������9T��x��?\T-B%�ë�&|�ؕ0h]܂Ι0""M�GEӪ�Aa;H��4�i7{��1�(i�/o�ed��?�/<�>j�i�ݺ.�z�=��]�����APqtD�=��LIIyc��,����A���w?�Wq�ϣ��'�m�/Jf�{8�~�#'�(X`c!�XV��J�;��Ou�9�Ǿl%��ݦ�?=}8ZBn���V�:p�%~�+���LM* B,���E��(��0g�����fd����B�A}��A]�'�R�aMⰄ����Z�(�nO1E�Γ��,^f�c���ҚL2�!�պ���i�b�^�����&'	(�(A��*�ֳ�p�0 sQAA���pDd8�Y#��[��Zv3���z�d�������XX^���P��������"岃[em����/B���L�B:M���qx�b�R?y9'FI*@W[b�ҜI���+���Q�D�PF�xR���K��qݧa�Q;��C��c9Hi�Ǎ����%zkm�A�`W�T����&�./��G�8��0���
��ٔ�EAo�7�����+֑�&;���붹v^�G��t�1��%	IQ����F��v��sa)0����2y��y��+<��J��u�;H10:��U��&+��1o��R!��־D@@x�Ȩ�ijj�ŖkImcI?몮R"�7�a����Ѓ�L��p�\��D�ϛp���� "�:��.(2`��������ɉHЋv1ܙ���oRT6s�ƃ�s����!�Y��
���7��iX�(���&Q��c��4��h�c�-z���й�>=���X�K��ym���¤� ��160����⫘���X��W��vx�_�[������m���F[�T�,��"�Xb���?cF7" i�i��ϟ�_�:b�f����]s}|R�ώ�:�����?9�D%�̍�YH�kN"�2�-����qs���*,LX�)Z3>��d�����PP��(z_�E`�mS�{�0�c�˛�����>[�\��Ȳ�7��T|��^�����(z�ْ�{�]��Pi��T.�&�3L+�����!!�ii?j�ZZ���{#���澨��7[<n�\�襡�C�+��E�644�K-��]����G��q�����qm��'�WW�˩Ve|�޸t\-&e��w���W��<�m�G�� �h[��)�"��Bn.��l����ss�`!�8�4�{ɠ���T6������I�x��t<e-S���i1���Z�����M���X��,���o�~ʃ�����ӟ�X\�4PHY�٭�P�Q���?����ԅ�<� [n���FZ,������Y�)����1�����&>���lId����c�10�}K��1Z�%	��f���}hc֬A,	�~f=S�a�S6~��9���6���g�
��N��c�%,��Wh��i����x���*D:b��'o���Z��e��Y`_7���Mz� �%ge�T�w%nr��4Ӆ6ѵ� G-����!��YJ�����;?�	�M�<M���9�x�-��c�>�NbU�D��K�n�'+10$;��{]Iu�q�f��m'��*|C��,n��	il|jrR���`0�rm_E�	�_�[�d�h�0�4���쓿��K'�״�����/��>�����c=|�!��o� jܫ̇`϶�	Uk7cc*���t%���^�HO'5h�*��ΥI;WZ�66u-��+b�JU]ܡ�ͻ�ϟMM]���Ͽ��V��H����
�/���n�%��@��D����@����1�q�,���B�%��ZZ)Yr�L�r��_/��{�#E6�H:�ةB$���M�"����o�������|�LR��Lii���sg��\��r���͋��و�@�B������%��,K�J�^�5?Ϭ0ZV���j��+;����BR�fR���<2�?��κ����s��.�Ʋ����?����,�)A%׎GNF������P�������x��=) ��1�J�{\˽[l��whO��-`N���.����L��¢J�E� Px;�������ʺ�٦�ǉ�lN�Ny&�ic��$�f=2��N�����DDħ�\��))�x�->�R9
�n'�}���U,�;�r��Y�W��a)�<=���[[�͖_S�|:���Amg���QZ]���SG�e3+��p�̛�#%��i<�ƿ+�2���Ϙ�1
@�'A�ɀX�|`��xq��WS��Qʦ�lJ�����v]'"��������䒆fX���w�ܭE�6��(��1>�Q�FYZ"���_$��� ���3&x�S���ɞ-Ak�����F�&'���_�b��,�����p�G4��R�3�������88���m��gBB%-�OL�1^�&p��XZ0�ܺ|$?��2�&󵬱���;?���4�[$�:��<ML)&�O,���:M���U����ja;q����^���zx{7O���aq�m9>vH�Z�Vj���3*;��a�n�d�Hmp9(`��xdPc�n�q��\��H�<�Vn{�2J�o@N��U�D�..�4��)<:֖���x�OMMw�=�T�t��.���Z����B�h(�-p�f���s ��KGP�#��|Y/�R�M���n����T�ZWx"�3����<�nЫ��K�m�Ã�)�te����2w�J7/��m1M�+k��'׶��zݞ��|��=&�&P���WT�L���j��}�E������^�]����ϧ��7�V]rŊ�2Trr
�3��o�	�Ӣ#D��V��&lG���L�M�ttPs��3���A���!�h��pۿ��Y��w�[J��v�P:׀�����AS�߿���'D��)(�����X�UT�	^��6yLdX�GFFڹ��jz�\Dn�B���l�
�S���w��XA�ɫ��2��3_�g��2��B	����粎������N.��ch@MmҰǈ>����# �Z:xBT�cm;�j��d������tk���Ub�H����&uL��9���%��b듦sK�B��&?ѓc�%�Hg��q�UcG0󛩱ѿ�F�]�{�����[��yVm�hu`#�y�E�=Xk��h��sl���0�������C�}p�*�Z�L�\E|s���;%77&��ϰ�q$Tt�o��O�ۦ����#Ҝ���}��'��V%�/nO��d����Fٙ�,J������Z�h ��4e_�������z���H0�j2�en犒�9�A��!J�P)���,����B(ge�d���QU����\��jp \�����n����#s��|?�*����x������fo�E��S9��� ����|�4��#c�}��ٱ�b(*��Dg3n��pgB$�W������=�`1×@�0��م��&F�v�����Q���t�ɨ��G�<�\��nΉ'���;�;��H���?v�LXZ�:��ã���>]�&Q�q����pbq�g�F�����bӴ�i�& 0��2x���d�U0l��aP<�ϕ�_K���4���p-�| ���Lwߦ�Z��t��mhX9�z�\��^��3����~lD����APAA��|E,��h��x���k�p�����i6c@6d��a㭌�A�4BY�G4M?�4���^���idV���ݿc���LN�>�w`��E��Çx�Yw�7H,R$�`&	ٜ��P����$ ��|���C#&Ҁ�A�K*Y����0\������%�Y.�r��n���<��ͩ��q����u�ڙG<��D���e6�
iM7$P�0jT�j�8<�Z1
�Q��\)�Y�ױxN�r'[ƻ���D(���P���%B��23����K �é2Vd#�"�۩j���6�M＆�TU_��Ed�S3��$ �u�dY��я;?22��Јۢ�n��mzZg���C��$	j�7L���?d�<�:t+�[6_iy�Os��kx$ k���@��f��2��U$݁� i�e�? m�O���:{�s�ͳṓ�q�2S�;ܥ�
�K�_�^��vI�w>}��������w�W��ַ�a�R���q@���RU>���3B������R.�����][v�y�o�G>|��&H���<,:���R�\��Q���`a���]3����ɶ%���KE�`�k~Σ̰�x&.66��v�gNq�\�P�~Z2Zt�{��?�ɝL�y C��� 7���RR����B�z1��]���Ў��tN�덉�
ӏ �:�Y���i���=���0xv�^50��I,"����U]q1�|�5<�t�'������y.�ۉ�y/����<�%oT�益r���z��AF�A�J�b����;ո�,�M�~9Q�m�u���>g7
�#���;!�B��Q���{t�G[K��浪�ü��\�D�'G�B��9�k����T�!�����P����u�����g���l�ͣ�H��z�:L�σ�,����Y�2`��s.���C=�:����B�뭮�A!&���ѡ!�H���V[>�����g�߁ܖv���8g���.)������d�Ŝƶ��vMj���χ��~�T���nEw��TGx[�T��+;�4����-��{j}@��R�F��{lw����W��yĔ��e��;#)^��U��焐�7���5!NT�l�!�F���ϓ��֖���(�23�E�`p��Dz%A��4��6##�rl�q/��LrZ�wbQg,��f����D���d���lJ�a����+��|֭(Z�vyHv||<
?;55�X����������	D��_��[�e{Y#�� Z�����I����n� F}�526����
B#-�I^�qoBKW�Q���@8p�u�z>�	D)�nr��'� y�����ڴmpJ�%�@����F�QO�Z&v�o�f�ҍa�-�%=���|{��mra`t�M,�����3j��Ń�,���-���������i^������e55����V@���ӳ��fZ2�$O:Q�-"/?h�CDL,s��a=����&!-�=��ʏ�"�B������y�%�c�{G��b�m���뇩����*m�F�����^�444Y��&��F���_�����G8�op�'��4��v>�i��d:� ���xANX�(��Ó ���\����F�E@�Θ����َ�3���{�_ �:�EPK��}}}m'�wx�8��}������9�9�8*��_ck�oxzy�T����SU�z�B��Sn��OGOߞ:���`����$���������nw�jEu����;R�������iQ��>>��Gۗ����wװl�"A��b��;������ ���l9݅�g��*{)nӣb�K�{5�3�/����>r-Pg���С����n�=mt�K:���;����H����<me�Aee�Wfrf�EE)��`Vb:��l1��̲�����ռ�Q� *nk�x����2�A*K�iUAUeA�0<����Q(��T�4�JB�sZ�i0�~��54ɦW(?��Lм�hXx�(k���E�v؀PM���������fBg�jG%lh��k?�����zTZa56sm�8�o�B��t\���ߤl��S��tm�a�l�<�f�+�Z���p6W �� ��@�ժ|��@�3+��h�e����.�����xB�>����d�������o{ٓ�|.��rB#����kk��b��+r�<���v�Vn��6s�2�\�jBwFwlE���ۙ����3
,hi�_�V�����<@��Yz�3w�h$6���q2�X�L�,1#v�sNN���d��Q�{�Ue>��"���2�33���ʈ�fw�} �t�@�>b���n��Ny,����1���Ӫ�Y�A��wCp71�.�U�x6�� �k�h7�u��1��㵼����%:�3�]��]jzz�"����Yݍh�'�K�蔻l@I����PI������FU����j$�����=͕=�+C8t��;5�0��V9����̣�Aឹ�c_'H���>j��l]dSF��T�X����Ӳ�L���k~�u�2V�H�3���~�J�������w�����v~�scRgw��\;u���4-Y��u��67���lW G�po�����r�)�Cg\����C/ʽO]��,�H�T�L�ڵ������f���ӭ�K�[���(4�nP��ȴ_j�X�l�E�,/np�|@�O�B��Y �b�FT���T�b�������be��SD �t~e������n�J1GMS�W�����&ˡsf�l�/�k�ߜ��no�	~s�7�F��d�B��Ω6����;��4�g4���`�ﵵ 2b��j���+v��P~%z:�6qR�GZ7���ɛͤc9a��O����Ԛیn(�E��8�ߴ�����5ɴTT��w�b�&�3�xI:����tC�g��D�������`�2N��-�l���3`�ax��SةUis��ct���;A���O.n�/,��\������ޗ��#p���o� Drv0�}AV��7y,�U�DXᓧYc36�fk�{�Ϭ�_����E�)�a)��*�;�� wÀ�K�g7�����2�N�DܗJt�=k�u��-n��|�Y��,��2r����7_�N�I���:QSWZ&�����ҙZ�vvh铥J)�$��َ�]�Z�g]��oUs5PU�=���������^jQ���� �s�{�����>ɛsuʭ3��j���w��Wf�S�=�a�Ճ&k���,�
�#���Ւr-&�T�Ծs�U��O/�މ�E0�+Әy\t4եD����X��{��|�� ��aq.e��J���k��=���߫�["�7��d%�?z�F�;<�$*���P����g������=�0�t��I��[&�b^FF�\,�|%��?@�Ѕl�ߛ:jWYTuL����|x?s �]/��솳���&(�za��ug�1����TI��MڦV7��^mVT�it��V��wq!d��/l�pd�j蛍GV�2.Qk�ʳ��u����g�N�;`�4���`>7�v�p\"�ps|�촭��#g�p����F��$�!����ZjXC�\�l�/�m˵��gnRx�u-�`|$���P������4>�P���B���4��gʗYPVP�����G�S�4�Y�q�r���qp�;+�&�,�cڤ��ʬ�Xo��dg���*�jWgy��8�g?�G�S/�_��a�-H%RP�%� �D>_�ϟ��W�
��G�+;^��F쀃�6?<J�,r��t\����OE�czyj�h�u˭����@�R#S�|N!�K�<�� �z�5C�,Ǔ��ʼ����H^��f��y�omm�fbw#�vO����8�(D7��=3�\����d�6A_~��w��-+�0�ig�Q�9�����2�4t(�Z�����>"~��;���Q� 943J崍3j:%IRrP�������I�|���T%��f�C|%�6.6��~
n�o��A.�O6(XȄK-�QI�?�)�8w�Dj��}�cA� ;Y��M� Ȭ��Q��x�E��Ф��{j*���c��mӔ�	`��a�vz-�;TPe����$�v�-|\sҡ��XzZ�䛋���8S%`l0@�QB�o4�����\��w������	��t=.(1Lڏ@C���`��ܜv} 5��q�Z/�kRRn{�P�\��q�ӗP�ݗq����||�/�b�-�Nē�[�F���z�4jɭ��{�	��pс��xI�x�ip�*���M��<]999���Z�'�?K�ཾaǛY�<��[dŠ�7��ÃO���l3�qx�do�Ս1�
ЉSaP͉פ5��w��
����*��766(��=g������Y-Z���=��Kx��������pDN߫_���t �1�����H��e/e��8��b/��H��	�a ��lh����0|�s�:6zJs�Y�����n��E>��fa��E��2������o��Yd���¿`g�3e⋩^�� �x�Q�uw����Nd�� ��m1,��47_X��J�9�
�p���aJ�&&i�0����E����n"���v�	�[��i�Ƴ�dh9F��5�7)�y-?��缽7���H���<.���g��A�w3?V�&^-uJ6]�(�nU�75)h ����$v���T.ޱw�ګ��2�vo�ʇT^���98x�����s����ٶ�p����!�Ys��G%
�Q��a��{�´ܹO#���ٳg��0�����F:#xa������.��N��kj:��Δ5�.��FLz"����F�����"�
W��//����v���GF����܉w��D�}���Q��'��ٯ�B0�60�K�J$��@�B����II�Iu
>>>Ѯ�@2���ֲ`#>��ۓ�y�����n]3s'��`�FWb~�?+���2�����ts�A��ž�F��YR�x_J��!&f(<
���|�f`�״���1~�d2�����sч����S�\���Y贆"���Y3]�{x�U���¼�Z�s��dH��?^��ǆ~-I �Yi��%��ՅW�Vw�}b���{vnc����;��=m݃�\�_9TT���:s>���E�p���$��z��6��
��f��Ғ/4G�M��l{��<��4����Ӄ(\F�_ccc�/If[�'���J�v��⻍6I�&���\\�x��@�k=�X�K���^c�dq�y�9�鈒�'ۖ+�o6O)K �O�G��TIңb��..��G7�#p�=�� z��m�X�q���11������ޞ��o���q1���bF|�ҁPψ�##���sX�榫x]�B�i/I��Ҩ��_�2���_��l�/�����.�g�� J�xu�x��N��
�W3�#��V(p������N7b�㦛S1���C;��|ެN�`��<�K��~s�����oq���k�����%��� A��*���&�-l��ٙ�7��;U1Y���]u�I���q���>���), 	��f�73ZQ�L�B���M]8���8��j6*�'�n�����S�_}}}F-��T�7곝����stC�kN�bNN췄ׄw�yEE�Sg�����f�wR\w�;�D�D,.�qs���Ohk{�M���Ⲡn�F�O��tX��鵕���FZrr�2���WMq1c&��|G�˫�wKF��?�4N�u�(0�π����pޛn���\P�j�uX��j��w"i��$�[j���E��P�nu��#.ݧs�=��fg{;M�zp���:܆�j�ۢN���]�V�JqaZ��X. ;�SM�gj�H䀬�y�Ze���U�/�z��6`xSm�����+G��I�����7_~VRRz�G��3Q�K'Ä���Y��.�"�0�=�OsB(3�>���RZu��-w*�d�g�a��Ae��KkkƧM� /iչ?�9��|Z'N�{N̛pz��=ٟRl1CW[��Zy�3�ƨ�����c-�>t�{2�5���:"ݒ���[1�QЂh���M�:���	����@��ٓ��?1��ܸ\;[-�L��������,�M'ה��P�p�x�б���u�F���o��J��
�v9'���H�e��D�z�>#��ϡD��������Ww7�,����o��7�����[��8��#���RPR��Kn��`�]G�w�^��E�ӣ�ļЮ�d����+���]��>% m%n���KЄtG�)��E'=l������|���⑲׃��a1�R��8Ov|���'��D�nK˴�̝t�� ISZ���� #'�v��oii�Б���2P�����|����oy���n�6�����zz���dy-?>��E_���gCB��;k[��"���P��}�ޛ�4���B\\<� �L�&Fz3�3�L/�c��IH"Q1��_�|����dH�D'f/�tqطU�݇;�0�阤�<�̬,L�Ǥ���||;Nh��L�W'xeG�����uX:�k8Cw�i�͓�g�Ֆ4�LOҽ�C:f���WDo���l[�4�e���Ǽ�'��vV���;�7V�v�f�p5����F�2 4�I�Z�� ��$s�rpr���c:�|�u8 'JW)���a�_/�g#�����+������_� ������7��&���G���W77+�����4��_�\ѫmg�a/U����ÿ�"w0з���.vF*T566����Q�8tU6]�ߖ��B�7^�±,S9�Դ��P�巗Tŝ�H{��35����?�]b���Շ�nnu��Պ��fV�6�cx��/�'����vww�陳>f�)��56�3<8��䐍�aQe6����{w�;&���8p�k��K�w""٨����k�kk�ġc�''� 㵵��l�Sex���u��/�����Q}���""݇�Z���4F���7$6%%P�f�;+�Jy��K�us�CKg5YFb*�L�#�2�h��.x��J'�g�2=?����E*�e�/9���X�)���5�a�o/Ө��v]���4W���n���s=\��mθ+�2NZ�{�-B7�&"���'s瀾RQ娕{��,43���4��|���{��y�L4�O�F����^�O
�s'�00��p߸���64���<>�-Rk&�������7�J&$���S>���F٦�'��J�����}q�2�A���"�t�Y�m��\�G�����ˬ�/�̒�������0j�$�)�������߂]��!`�DDD�~?Rz�P��$W����6��t�E��t6�ߥ�Vdt����fTTT�շ��t��>R43B���6�����)�](��H�p���d�}'K���R�����A�J;��^?����nmy0ᛷ�ɐ �;tu�����6&OOO����"]���]�X���^��	��x%����u�������-���hTQ��Z�-L���omlJ@/S置��-�?]��J��p�_��밖T�s@��� y��� -ߛ��
���2ig$1�a�����qx�X�I��s4�n.(��˦�R�N�wM��M���j�ccê6���b�[Wg'H���EE�1pqݎN�4��3������h455��Nd�GZZ�7z<����	mx���o]R� �7,��r�������R�1�F��A����|��v [g8*a���뭴�]fwD��+�:3C8g`�%-�ׯ�%���ϚC8�*z��[
#V|���9��99G<r2�IH�d���^XHo`�@�vBd�`�o��֖��o�55@������/������w�vE~ �q4�9������F<ݜz�e3+��\�F��ð�<��۷pmmm_��@U3���eeeX��@�(�WT�8I���"F�E>1+
2����dh/��y�:ƙ�q	������_��u� ]�s4���_�<Za>���x� +���?VFCC���J�'K&$���珖;��p��=Ǩ/�Ffs���ʕ�ETO@�[����jJ
�0$��͐�]@��`�*� Żn+M:�WtA�-��@�z}�}�o�� �����O6�sv7��F��0C?�p�u��Q@��حF_X�TuD����Cc��5�tU⏨�dEGL�Љ��)��&�P���&V�~wĶ�y� (��wy�i����w��..��_���n����/ P��sP�Q�6�6��,
_�=;6^���������MIIAaJ}�Ow��X�3�ޔ�}���>L��,���}�=��W$@�B7���
��i���D��f���5�P����s�����d�w�	8,�\���	���a�!ƻ3��'�c�l�����\
�'U\aLR���z�.�pr�rD �!�a�|�;s�������w��x�|�^ a���dy�⧡8�aa�/���yള�w�����-���%:U�л�&ɕkg���DcE��)�D���ax߅�P�"����ii4~45|�M�k8G�#���-:FPcW�a��<�.������Zy'З��ܯ((���k+�'pO6�
	����hňƐ�������� P����񏈐d���+Mgnk�^���!I4��'�W�5�Ш������/5��:�X[Z�u+&�f�mp�΋:��iLd��v�3d��gO��*�~���u�H�6<�Y���=t�n��J0�mxaXX�t�৏����G����\����4�q�xW~�Y���Jһ�n���w�<Y��3�۷z�?���������t���r�����ƅ�.Vn�$�f�|I�vy��9�͖�x_2���ݛ�;�z������oH|Hْ��V��ٽ�����{O���X�E��ԙ�#����O��/�G�y�Y���CCJe��	����%�����K$���ߚ`6X�n��0КBI
���A�l�9m=��I��xL|Oԛ輫�j��ho�
��2
P�s���*6�w��3��s�P��6�=�PG��h��7���EI�6���c��b���˿�q[@�F�>t�6�Ŀq�}I����g)5+�K��P�m U��
t�իW U-�}||DE��,,R	p���݀�M��6���J�1k��d�
�zxdiJ#�ʚ,��5(�DFF��^��,�BOK�z�kh+�з�P����ї%%%�{�����^���N=��#�Q$~~~���(I4�Lj��%�V��e��t� �u[�12�(nM����I����K�h�����7���p8���#.���\��d��mo������Y!Ao" ��Ѷ�������@��
,�7xy����NVV����`�9����w,F)�}IOg�q�B8im#7�<"�By�ZSP���(�Mo�V�q�<���`�������WQ{r=����KrCyy�T�j�d�8�б8iS�H�����*��C��"��u]ZVRX����hS:��c�R�5vpdH����F?q~�2�<,� h�O޼@��������;/ⶄ�>H��_>b��X*be?r3�,E�����۱w��G,��A�*��`���ֱ�����1�yiu�3t4��XDA@ZZZ�n-���>�4@,2�Vn��N��@�
�֩)u�"�G��"���01i�S¸M� )7\�v: �Dނ�!�#����L���U��psrr������Y�������u����ڪu9H]J��G?��Z ��/�sb��s1݃�];��u�J'�V��?�����I��͍���a��� ڟ>e�g�s��>kO�m�
���%���
	x����M�itt4��gO���i�iaoL'6K �
X"����M��[S��+V*�@􈈊RF��|��������~�.ȓM]��!�Pa�Y� )��dy6Sv�Ԣ9�5��K�@S���ݽ�kG���8��WH����pn���:!a�	^��z_2�
� �%�~R0�������ީ��s��8[C�rd�sձ�oӚU���1yo���Ɣ��^����,ɹ2�����\6 b�Jm���V�F���4�ROٖ��~�=�ӊ�w� ���Y-%���|�H�P�c�b���[oF�ީR]�Ƴ��k��UF+�¼Z�1{u2X�eZ�Q&����i���%	|�L��
� |fU�?a�`i��h"""��|����*��( � ��?ň���,i���?xKAA�����!8#n�q6d=�W�4���@!�m�4��G	!��q��o�F/Y�^S7sFX��ζR�9���s@��*ыg�8�A�����v9�*�l�#�NgI�P����V��$����92�0AB&�0��wVjZM�9*��N �N�@聡ea���'Ŷ���'po$;%o���+)ʔ3����4�wu���_��Xͅ��2���~!����M�AB�	�����s�tC��p���Pf��;����*y{�Ma���붾�<_�ZpGJ��a�vg����k)�dA��Tv�J�ѧ'7h�@��UWOħ��m%#�*�@j�^Fǆ	�A��<K�gڪ���)X�5�WlTTTj�N�_�H8��%��g/�!���ܲ��[���c�N4�m��2F���� �L̏j�b�i_��s\� �������%��j^!�c��,W�	7==}�ms�^��Ix�;
��L���oJ^M�D�~Pƚ���026�o�u-Lv�d��t^�}⍈�����&�އ�zF�4�=Ж����.P���I���+������	�f��0<�w�¾�(�Z ��Md{.����C����]jo�%�t:��
��Tf�jq'���e�U����S��E����v�d���oo]�J��ɡ�@�DK4c��ړSS��ߺ7�O�� �*E?`{s��A�N����e�w�F�1 ��&����dάnl�p�R���f�x]JB�6ۣ=���'����1밦�A��R�P�I�t�mTM^Sք�[�Y�.���w�OZ'��T�2�-@Eˁ��v�.?�����2
ٲ�A�^�b�u�����,����c@���j��*��D�!{8T��'�矆��\��	�jj��֏s>����������:ա	�
	�"��-� ���9����t3��`�̻	�
3䓩\x�i5j��ف�/�]蓁a
��oC�����(;މ]G�/�G��Ti�_�4��~�룽��n;��is2�����}MH�J�L�ii;�*L_~���K�Cf񇺺:� UYF�P���GH�.F��{n��PW	��
�]x��O�P�a3�����m��s66L�����KK�cא��n�hZ�jpa�!�U**򪱑�7U OE��h�����P���Ђ��W��� l�Dw�{����u��;łw����0���x��@�����W#h��7�V�j���>.�Z0�����Y��p��)ާ_�^S��>Χ�ʳЗ�� �C|-��m����O��R��ѣGf��Y���?~�3�6����Q�d3�� �w�U���.��6��ӪwB�ac,Wzd�.S!��X�h���FE����������$s�@�SVQ	������Dz�ڈOJ9 /�&2/g,T��Z�Ɗ? ���_�N+U�Q�X�RR���Dd���I>-�&���)�>�Ȁ��ū[�rZ�#���z�?U���8�����n"��|�FGVd��y� ��#�G Jp��*�#��TJ}٠�����ؤ�7�w�iݶ�D����?ʲ�C�����~�杪����zb؊�9���T^7L���t��^�AX^��a��ByF/X���Mɠ�E���gl\\rZsR?\��$%����-"~�5;;��ٻ��iM�o�s��&LKAZ���O�6,��9�			���.�i�ZH~�/�f��'���ݼMj������uNNx ����˗�k#��.�Z�&�J��8��t*ԕ��c��:s#-;~���h	���󉅮׻�����D�M����D7#����ڷ��g;WlP �x���O��"� O ��iM��C�UT�u]��n)����i��n��.)�ni���o.����{g朳c������X!�s��R�U#}uyMb��$��4�~6��60���NoK�������-@�|��D��{ "R%�E�{��d9QQH��#R��v��+ggN�-n;cd�Q�^}f߀�v n���Vy���bҳ;0{�|�|���a�3p�����
�d����4_QF9����»��T���E����U!(qd������2殞��u��s�<�	��p���X�_~��(��F�_ݡF�O�X!�Qp��y� _)���\lV�F~~ua�\����#.)IJd@�D�ʝ7�c�)�&���䄲,1)�m�������)8��kF����oBRRq�xvFz&&p����Nȩ�`0׏..��*���D��I�ґA3��z#gp�!!�M��X��u��B�	f�C�6!͜��~/
�R�;.��4��2ƕ�U���F�*�-�^��ʶ0@��nQ��Ɯ���z� ׷��$rqu��(T�b�<�)+c�akc���L�5+=U�0�l	�k�;bu��Y�ϱ�^�������X��j��'�p¤�������~:ff&�;͒K�����JHP&����;�9o�$ڮv�9]Ūy4���#ox1�.����0oW,c� !���?�$
���\{��򂙏/���b9d��qi`�5�ê>�H��̽����W��{h�577�B��/�
(��h�,�\��т���X�<ɏ��@/T?d�Y3 гx���������۫�J~��q��S���ny-%��@Z-�������?*^��D�&
�l��-P'y�uj�����#s{����_�G%�m�QN�|���pλD�f$i�n0�ޗ���M�"�~��ٷ�"�|2%�1FD���:�������ϝkjj���МFC''�NQQN��MaϏDv�9�T������9�ɴ�����z|�G�d8�R�g�ws��j����r�a�@�(��o}=w�'ӟ,FN8��� Ϧ�ch���m�'��:� ܱ���_NC#$g�lD�:Sƹ�US��bl'��e�=�� 9ʜƼ�f�oh�b��ԲLv��ggf~��^U���� S��;scm'�@͊	�sė3n"���5�0Q�K^��àK���	�����<n����KG$�/.�B�:d�����񱵢�1�@�K�u|X/LؔK5����^薓�ej��[�&'�;���y���L��MFX]-Ck��jqss9l��oo��x����4�o��6�w���a��f������ׯ�Q��5����&Q
�@�*��M�����Ghf�:j�gf�c�������. �A+ԏk��l���~�x]��3����� ��jK�pϓ `g�i��/����a;'�?�C�6.12W�=uZ��l�$%=��`d.!aW��ȄuXZ��9B(���z܅��㓓��+�#�0#M�h�,	ډ<\���g�+�C��ބ�"�v*��d}lMI�@!=S!&�ȁq���_�0��s���ܩj�R�d(�-��S�zLQP��"�q�#���g���p�dvC�Bb��
�+߾bڐ�h�C�e�塽2LN5=}}��+h�?4�>��c�����ɮxr�S�YuԐE�n���ͻ)I"4"���q�'$����cBBgё��g������y��EL2�������������Xܹ`PwFO���}1?��SG`?�J\Z�����?b�ڄ��CJD�<)� ��T�{MAp�TXH�����d����h�M�y`1})�ִ�����yyB��Q1ř�����>ӆ@�����*�QE��j����زΥ%�M䃃��Ώ I�����N���m�����>"$���)��8��x���i�..F �|����L�wO�/mս��Ɔ�V2ו��������A>���Ŧp�[w�v�#���x{_��{3���kt���h�����C�$��U�/}!s��v4=�v�x:a��T��/R~�ڧsmcCWV�o��<*
5s��H��	))"��x""_�kQD�DA*��Ύ��wR�LJj�7Ue���������'g���iU��4��r���Ծzlz���f�5%�n�qK��r�f$����G��֬�
�ٮQ�dK�����Н�y�|k􊌾#�M����!c��n�p�Ma�e%mC /���~��#cm��đ��F�����Gs���hwcccY�)J�RL��I�Ur�Q^����!c�Ɣ�onB۫Q���S��>�r�������_�I�L�O{*1L�Q@ �3���\߷�6�݉L�����ܓA_c���1�*����Vi���<��e��� Ĉ��P�fy�6���
s���a�N��L�dL($�C��?�D:jt���UIq[��~�p\/W"�L>�pکә*������i��H��k��)�`�54��cb���^��̀�EKG׾ ����ly���)�߸ �m#/﫠������L�h�ʳՖ�l�<��H�G?ɱ>	|\I	���k�2H� pK�u*<��h.S�dhXX�b��r�=��C�����"�(P&�pr�(b "���27��UlGI;Y_X̘+c�c2��j��:����h��x��}�o{u�������׿��lmm	HJ��0'J�̼J�47�M��������>;�|���������py��RHP�/x>mh6r� �#;�`���0�t_#�h,1���{�:�����Ȝ#d��6�'C��A�|	\�%T��cGXz)nZ�V�����ZaV��;��RQQ�l(�*�w�P�8�V/�''���w�ˉZ��#���iQ��7�_�i�! ����`�9�ٱݰ���_�%ˮɺ/�ǈBJ)��Rjy�S#�h�h넱��XT
 �����om�+��m!��	M$��e���S頌R u�l,,,N���-|����S^&&�"$��3x��q�r��M���3�x/,hC��x)��R���$������2���)	��+g��k���Y2��kiYc01k�Ad�r&1&*��L�}Z�J�A�?icii�����0{ޟb�y��r���� �O�13��q P�?]A��"豲�BY����\T�^����N�}t�$j�b�@v�t ��R+�g�u5�����6���i-�m����Ţ1'�>Ev^+ϛK=�
q��R.o`X�F ��&��U� ����|�5j8>��FR�o�U�Y�����Su�,�(�j��&6�, ]�H�}{9�Ο����}=�U�ՙb3&.���㪍��$��%��ǑqqP����쬵��Fnn������������R�L�3���III�c%�1�J�+�&AM�C��Z��t(0��7����cOܐ�f������gb8pĨܷIBB�1��ޥ�
�gr�rvJ��
ƾ�^\�=1�:�_����������j���huӊ$���
��+ͱ�uq))_�{��)��\خ�N��ZpĲ�bW���N���R��biTZ�^ו44����`b7�0���7�w؛|�q���z�x��_��]���8��<6��ԓ��p�_�B��h}�W�=��"��!�[�44�%�����H�mlЂ��?�݁�FE%�h5�����}�S��ڈ��"]�s��y��������/_M-%��U�n��H��un�����=��������
r�"���'z���ふ���ɡ�0uDD~c�q%�Q3o?�Q� E�73�4s�����n�a��P���;`�cm��0f4��}�%A��!���������7�L��M��3u�H�NJ�W&�~z� I�J#���UU�r�^��E=ym���'�;�:���o��000��̧�v~h�8�w=�[�h�ɚ�N�PJ��r��`c����ƺ�2W>���޳y��v0��x��dye�w��HS�H �D�6uL��0IH��s|���;_�jA�_�����@��aaHs�w��X�An��t�ZP%ʻ_�1��+FbT�&J4����==�w��ţs��ݜ\]I��浶n~�rww�IO#*$�r�muuuJ��B6�ni���es�z0T�X�E9�D��.���� _	{��0����.���xyC?��GFF�zL$��Z$����2+*��	����mmmM�1�f����$:����צm�O��dCuV,F&&Ԋ�&���
ڣ�㐢޽!�Z��Á;;�"�:�#Ͽ�qpp������Cr�������]4��pc��IQp��'}�����æ�TM��&q(i�2JJ��y<~�B�@���)�<��{�ɾ_���g,�����:�W���ީ�2�Z��g�0�r�)U���+�]Il��<��_���m�$C�o��g��o	I�?��_J�����KC�TQU3� ;.�fe�Gg0搢	
���5����EY!��ۦY��o������eė���P�����e���J�<�~W��	�o�f��^DLc���2�|�aas
��#{�q�*ޛ���U��T��K�6< "������✞}k��j�ڝ���
�R�? ������I��b���K�6)
L�5���N�,�������
�h ���, p��V$8&�Vj�����U��el�ٺ�h^:¬�v�_V��t}{���fS��5���Jlq��B"���0,��-Dl��c���D������*��/om���sj����#%���9���Rl*kjV��Ls�J5Z!�_�g��~���;���0�g���Xe��������UC���v���a���(�(_�A���Gϲ���[���E%$����5
y����/5ؐz��[��+Kt��bbkgG� Mo߂n0m&��o���Ȋ������h㊙��YD���|���l'��W}�4���k-���բ������R�ɕ��(�\+Y$)���`� �)=����� ��_�ZTX�ԢN���׼%�-�fot�J���~���c
*jNK�Ko0\\\��d ��ӝ`ǕW�֕�<=��D�Ȯ��<�%�Eld� ���i}0_9��q�v�H.�9^O-R$ 쬸耒�0��8�������%��
c�2;�S ������&�_GI�?�C��șE�����iF7A� �$k����hi�2�Q.UEH�O�jjl�,��E��:��==7�n�[�.�� ��[dn/e�[^�����*���6T��9��e0\T����MMW��G�B����M͈���&B�(6u���4�[ut�*@*�R!IT��9�kR{�!��"	:�^��ʴ�?}/u�M~3���*�8�pNJII-U��X�F˾������h�[^^V5!��#����y�ਦ@ ��5�x������k���<���kux͟=G��<�| ��`�?�{�ܖ��a�EΏ����&���륦R?����4��`�5�%a�S�n(�J�t�.xܘЬ�$<�@�;G����Kw�����r+������Ƹve�M�M ~A[i4Xߑ��L�$��Y���2h��B�ʽ��?�p������<��^ #���#=_�z$�W2��$<���t��@X�0�kW����_x�F�@׾�`�R **��"}æ��%�):���j�����ȳ�/���)e�އ��W,���V'b��,�(ѣ���������%�&Y�D�i����UH� L��P0(f;�wi"�����\�67?����9t~���Q���M���ʀѸ�\�T���<��c������[��A-,,��t�Lu��������y�+���W4��c��C+��t���'��?n"q����j�4$�����������ABDLLA��|�cvmA�&h ���˨J�Uo )ao�,4׺n��P&��d�������l���L'��K ���I��23[�=' ��Q`C��j�4 �0�wǰ���a�r*1�'�A�B}+�A4HH�k�(�c�o��6����72d���������F���$��i���H�t.}u	�4$�}��н�bv�\���q�.v�zBHo�,#��#�rff4��ﯠ-衞�x4xoF���')��4�Ã��_�8��mw0��h
�9 	�*�/�s.�,(��utgX]ճ4 �&��e�����Ucm9"[v��H��h���5�%ț��م�d�����0�{��%C�Q{��½����N�5J�(s��d#+�V)��)�jjr�bb��C���裶��,���b�?Phǒ��gms��Y{��t@�J�P����!O�fHR2���`�ʆ��s�=�KppTL�*FV;�J��Q�w�/_ ��;��1'�j��j���� #!�]�g67�ư:��t~g���D^�WI�%F<'' ��^��Q2 D �iǤ0+�S7p�p������G��3d(}����?m	�/�_��V����?����È��b��C6&&ow�:|W���!��wb�I �ł
y���5i9�u��M�\�B֨�fz�]]]rZJ��f������ �Y6cɯ���%���+����ʒh�������Qxb��W~�z~^���7��2�u6��ػ��mmm�icx��u�l��Y9����	/i����w<��(�v9��(�@j��Ba�&���.���̹K~"W<d��%9	U#?��Lo䵔�/��߁~
g|\	TA��Y*�<u��Asrq�(,���f��y葈1����� zϪ��Cd�Mwj��SUU%.)����)��5<::�q�X�R��~A$���]ny��v|���������E	;W'�x=33��Y�]��.M~---���q��Z����.i��C<?mȚ��/�ɝ�<��r�����~K� �שK[�� �}_Щ��Vi��~(��" pZce�S�>>�!8�`�0�ng�~fjk342�V��2��w��tDd���TH��?��gQI@O�{�0Nb*.X�xo'd�)z��)q�C)��W�pKIf���_&ğ6�,'W��N}�ÓTT���ʙ69h�P
�H�8t%�Ba�5�t;�~�$��@L��sڡK�Q�h���-�5lb�p�~w2[@^@�l�a-8$X���ܣ��� �{�t|U�(w��(w	Ro���o�[  �С����j��ޟ�����	�$D��eZ�eSC���{���< 4���7ŀ }*[�x)�b1Y����a��Db.���*?��r
�RMo� ;�GN�ӓ���4� ��j���i��
�޸�����>@���;�B��m�OyDpL|�3ź�����*^Ը�8�8���C�ɖϷ���}�������M��c.6��G����"F�? k(���KLGv��տ��y��g���ӷ~��,?'�D��?e��V��#C胷 \+z�墘��<��W� K�9a��k�?b�0]Y]-w:������I�ٱRS�Ť�{�f(�e
j��� ���5Q
P�	����J�`^X���1=W`%�@"6�����h�g�?0P<���3��A]�^��7ͬ�+���X ��� 5: :	�cB��*Ő���=a`>;"ώ �W��~?�B���֏"�����5`���]�"{8K���Ck~����Jn��X� �}�m[� H8H�S�2b<# q����|��Ą�]wg���tE(b}�tYDh�_ٞ��`�w�UC���6�ș��>Q�Y�to�4�l�zPe�V��Y�v�r��������Z��z
(���T��\��>�mJ�<���+k���BH�����Q��f�À|���i�DX���s��#BM�aEBC�.����@.������B�f �&1���}�8;�h��O���,k�j�Pk�Rィ���g�f�|?7���-C��u�/ʲĴ��aR�� ����9���^�� �4t`sB�LPޚ����hzLg��ۑo�"����'~��N��N-�<I��f.Ƀ\` �f�7���h�_ *�� G����ъm�����I�Gpla�H�W��B�H�Jt�؋R/7L׿�NC?��>��"��4���Ш���C27�abL�)�_H�J������yJ�ŅȮ�##m=7b
6h�Ԙ"$�œ@�p�:��F������g���,�?}j-�5Zlr&&T	�*��?m��5}C�d���ՏT���@���ޥ����b�nD2Z��ܜR�rhq�p)����Q�4�<�0RY���c�)C�����1�[��$+R�� �fgo�e�5�W"blL�Ζ��-G�T09�ce��##Y���w�0�����(UU JJ)WX��M�,!+`%���tpp_-�WVV�PET�Qۅ�m��ǃT���$6c3����������p;�Dqu��d�6����7�t��e�!�)�yR
�� ���w�	4*�Z�Hj��c��L���:��,O5`��k���&��%������?�F%+��A2v�H��@������ X9�!���|���B���W�,F ��n��l�<����{���\�fA�`����H������� �%%!��/$�Ӯ���Q`�L8�������� ���:Qn(C�Ƭ��!���S-;���:8�Y|迒�R�r������$ѩ�^�%%H�--�@���<�� ��:AM�ZE�B��/-��ak��@!W#�s�! g����,��t� ��"<|�W��X�ٵ9�\�1���z�g����w�P�XuO��^p��!RW�577�L�����% d�LJ��8T�s<`���N�~~B��{n���N��*T��ݡr��\������-��_�
�׫��f&{C>ϴ?m���T6Ҍ���V�O�D�u4�W��k����ߡ�b����
�l��2�(}�
Ppǚ�MML2�ʖ ����4|"#Q�s��[�<�vF)�&�u�ǜx�G�����J�4^	�bv�	�ObP ���ۋt�74,TA��s���.�l�����8
�eO�����ܪNbXKmmm'6OdB��O�M��~�)��f��-�k �W���4��� F�sbC�������������Y��������7���5=	Z���͕�u� Vƣ+7��rPm�)xo���޽�)N�<CF^�d������HE��0��f�'Ibœ�V�e��o&B�=�����N"�74�� �̈��u�S}C�Ls�<S������ ��t_���g�^���J���	'_&UHH����/���Y�� 3�:w�Āù�;���\�	^^&�����	M�Bӫ�����,-\������@O��i�pv;�I���=�p`lL�r��V]����1�J����\��lFH��3&Y+�o�;�dbfֽxz���_2� ����927 ���/_PQQ?������#��L_����K �y�'��'=��,,,���
�8b_7�T�^�O��E��@f����S-)_�Y=&�� m���:�a�Y�\̕��ˤ-����?H{��'ږ��AAMo�l�hE�<�W����1ߕ6� ^Ik7��i�T��.rZZ� nh���_S�����G�0Qb#/+0�&Bp�I�(q�;-�h!We�O�'5��s��o�)�:�Xu5; ^m�mx{�ef��!i�I���s�v5T�4�`���V��O�}i�_œl@����F�Do��=��;C�ͺA���Ê:W��1���,�M���j5�Vr��gJ�u}%�� b�Zm�fz>�5פ5�J�>`H���q�����;:D�5�s����>\#�.�->��C��!2t�5pp�Y��H�~H��k�|O]uU��[��/���k6�M[��a��gȽ�{I�4?�E�����ƀ@]s�����[�1C\�G����ԃ�oj��d\bdL�[�+�O
����BҺ7��cD�d�Cױ�PPU1�SKL46��.zA�$��Eဗ0qs+��q�X�,et]r,ʁJ`2_@j��p��J5�G@��;�/�� �"x:C���Yk���~������C�w{�����z���B��8��@�E�K�d���.�c%WE;o��~{��qjl���ؿ���9aJ��pӦ&�o'���
%_�s��=�?r�~S�TAQQr�ٿ���i�d��@�=V�����}|����JJD��E�i|���-�=\j��)x�ŭx��	����~CV6���(Ԝ��d.�Јc%���5Ĳ�����ד� ���	� ��5V��[��n��3�����*���w�UV?�8�3� �*@���p Ȝ���Wn�������$2�@�ǟ�mܑ�SQ����M�C�l�Z�v5�_�C�*�~qj�zK�phL �Q������6Km����;��Ƨ�$?�l�����cۗ�
�F��4w�����{��!�M�<rAAJ:�ܘ� �~�H��q�EdT��;J��iw�z�@�$&"�!�[y��r��l-F�5��+��Z��\pU����5>c��'Ԛw-��3�B�����|pɃ�yKI	"��z����6���|����P}�q	��%�n��+��C|~�Ʀĵ�37��.���k0	X�W�IRon�o���#N�rdO�h;�OM�b���-Hf0 ��%&�t�w-6��v��"�z�L]��������T.<��
�r�n���h\RTR�	�.��a	�ζ����^��A����%����Z/$wfY,�U��P$%UI&&oh�%��Dgwv�F?�[�vD֍�УD<��[�_==	J�,��_N~�hV�g�v�ᗟ&�S᷿��!W�Q�2ȐX3~�ծ��ж�p��*�p\��3�� �*#��=t��@��Ì	]�xkI��ys�
��ܼ���<0��R{[�A >��)+G ���E�7�?&�[C>�S�m�֏����]%���Z�[L8����S��{����������Yk���^IqJM�&%�Jn��/��.uZ6�p]���p���])Ho�5p@��<��J*@����:7?�ݜ�]NUQ�Z������Xn��_"����㛄$��U�|���Z���p��`�����#�G߹����'�e)~�f������4�qg�bhƷ|8 q�����a��sp����QY�q*�/R.6EVUn�?lܡ-�۞$x���˛��r8 ���Y���!C�m�ë#gP�|ה�!���l��׵�~��c.�º@���0� �D�bO@1��D����+6���4��ݮlS�QWT6��W`��Kj	��o�<��9RO���5�Ҍ��=j_����fM���+�+�����9�btm��付;$�`ܰ���$��Sܥ���%dI�+��� 4�U�Kl7�V�.P)�)�����? �����W���T�4JL�tޟa"�'�@�l�-]Bf��at�[�y�WL.���^���tl@�Ο����:$��XTʹ�E���j���ܷ(j���da��#��\����'b{笑��B�2�h��P�T��9h)T��]�;0R����4"N�n�eA�]˂&���Iv���V��E�;���4��s;=4]l�/�Z�:�6EOȵj�~���[^��JS]��b V�9Ml�S�[t	�.@���y�����tt���u�z"$�~p���?/�����z���v]v`O����Ŷ-)2��R��@ǭ펉Vرa�z�n$�����n;�wE�P�p�bf�2ف�G�?��~:��5)���[S]��Q1)��_^&�X�&����U���m�466��2��m?��2����#�w�2a~p���7ɽ����Ῑ��<�.�66�Z�^�5�Bχ�&$1XAJJJ�@Wa���c�Sx]F6�]�p��������Ɨ�q��#�űGL�k)��D�W�;�=�����4"�Z$����*$��o�z�GD�R+��\�(a�^�4R,�.S�S�~%�|�o.Z���j���r(F�����>F$�Y�죄?~��nJ�V:�R�u����9E�	q^��x�%���[Y�I���!�ם���J�1~{�s��b�����Y��_7x��8��M��\	,�b}����U7�Q2(�S���/��w'�&+��7Aa䛂^`&�K:�O��F�5`��%Y�<��l�c�z�e����(3�c�+���֨,�NY��.��c
?g�ܽχ�oꄆa����=\ 2A���{j��E�"�A �)�YZ��E�X gP�} �]|Y��Q�,�M�5T�Us:(��a����?������Y�pE;�A�E�˟��N��o�'G�j��RMy�]/����ٱ���ԥ����
(i@/��8K��v\ͼ�B�YѺX8π-��f�O!�A��y��y��������m��ǧo_EXL��6u�(���z�������]�Уc��W���ʯ�S�{[��v�ـ�<�g�ui)���������:�|DSw�i���aL,n_j݁�I���N�b�e��Sb�c����v�OӺ�O��G����~��;<|���'<�d��ҷ�[���CanŮ��3O˃E�����vB� �
�QH^10��F~%s�i�>n�Z�=p��k%Z�C{�z���
& ��jA10�p�f�� ��W��]��o� g��J�dh�.t�=vh��`KM^����ɭd>�a����:,� ���M�x	A�4-+wI���W�j���[Xu��|S�쬔�`3��8���	���%�de���5^�J�?d���:"7g9���bM��ͷf�M�ĺ�*D�[q C9r��X��b���s��a��1��PU)���^Tll�eIT�_�o{���?|#$}�R%mo��3m��QK �Ű�i��IR�>���V/�"�@�g��|�5.�w�>�\]eV6�*�u��!,\�k\�!��7��*u�{���4� NZ&c�^`=릻q��~��y�<��v�*Ev'J���wu����� Ẑ6`5����=�������qv
خv!�ħqآ��M�s��LG3#q���7	���7�;yzܔ腪�7�ւ�ɘ�oܴ��������xۮ��¥n2H�x�D���Jpp��2/�)D)�4Xf�:���orM�=3^���I�56��ğ��ZV=��l��矗*"�]M_Y��x�Ԭ���H�}��F�u6����
NNN�Mbdh����MM�Х��W�����}�ݡrE�}菗��s�A�X�E��P��o�]+�(���]RUiŜD8w��Ŭ�R�p� 
�%W�ZZc�]]]�e�ȄWH"��t�#|Y�W�ٹ:FggC6��s`�&�-|��O]`����g<��`���7�[t#��p�v���-���O�h[{�3��(�\��Cm��!�T� Xԕd�i_Pu�.��Y����n:l�k�|��I m3iQ➏�,����@����� Q�J��Ѩ	��)~��))2^.V��-;���a��曦�:y��xkn�&�Ԁ���� w:�mR�a�|z��t,쨁����ɀ����{G��f(5�^��N��~�ӱ\v���%sXd����b������-���Vz,�{R���~s�UF����4�pv�bpK�/X�y���WD���( ^'6��oJH���BU��\�KYDY3m�� ��T�b��sm�[mP�<`N�'��K��ոs�!5�@���9�@��k�<j���;Y����2ܗ/_��jF5�뜎Ib:�C�xп΅���Kߜm]~:�l�������Hv�QTYfA����4��|���t�o;�����y{���;".'���}/����߈�oY��n���U�A��
e5s���٬ac�I�������������Y�Y!���J�\�·� �U��C�J�����JD��-u3�(d6�ΆOH˜�뇯�G5]���0ķ7��e7���a�! #g�8-�)ض�v�C`�i@�#^��C~.�	��Q�����_������C7<����W�o�y������(d4�M!C�N���7�)L5�g�NLT���gz�Yŕ��\=K�M�9M��S�`vv>HQ(�o{w7d/�f����B�Ҭ����\�Z��E5i���^7`L[yzd"���`![ݸ��^�O�>|�����9�{T��9X6�۠FMR>��
g
���_g��s�iݞ�g�T�庐�zz�o]�H����ʔ(��̴ܺ��w�777�eE���*�{FGџ*��Xk�%j>hA�W�UM��.�p�s3tÁ������f|<<��>5�_}Tp���gG����-� ��=��w~c$�����o###�*�S����F�ۃX[!Y5WŎ�ED�S��w���|o�_�s�m�,�Z��E��h�La���5xy7_���8������M�G9^�vʿ\۩9��#�w��X6*�Y#(��������ȅ�?W������T~^��&��X�3��ړ�w�Ϗ���5�����Չ�GP����{�{��e~��=�vV�%%'�i��h�q�L�XPXU��=��Brr�$$$�e�!�0���^\��쌫<j��T�<�~���
e1C�A��X[���0����E�$G�˫��@���628Ԏ8�.k�R%fdD�ï��]���n@}��c?��s&E�>�wt�W�Ku31)��\ᑗ������Ĭ��}Ee��ؘ�\���V�y�)Nvtv&������	%%f,�Ħ+.�;?( �#-L󷽱���B�/���"����7`ͪ��G�R*��$�Z�P�͛7C�aFf.��i�U���̭�<�` ������q���J�;E"��>��4K�Υ��##f�X��������}0k����Dx����i:�l�Aȓ����H�md������(o��qM:o�ǛW��I�����:����ޖ���Gkȫ��j�tt�ΌP�*�h<�I�.�㭇��(�zP�Nv?v{-\4>�b�X���'����B$����g ���m��m?��($�:�-���ҝ������ry qw\��?��϶G+����VWV�C< �����.w��o ���EEUX��5`�TB{��X�e���̼1[�l��f��iB&�������p�5660+r�no~3��d@�j�^��Jg�[lN�_z��ٙZ���f����IE=�������Y�wQ׆X�gȫ�@Mr���rt7 �P_�{6S�t��w�U�NC�|9����"� @	�J�lğLm� �w{mԢ�Z#+�ub"���[:_�<i�/&Q�>�7�=:�к����Εw� ͓/���AZtTN��Su�>kТ(�E_�|�R�r;m����Y1������''�O��+t�39�oҏ;t�����;^\�gj���P��oh6`��o��ݩ�7��b�������͟K���Ύ!���S�8Á�Y����O�X�*�X����ʥ�<yh���4*&E�zcc�oϬ�pc���3��g��[Q�����\�~
��<�ma!�ǈ���l~g���f$�OY��`�c�@}ϛ�U�1�L��]�����������::.'?����r��Y�y�.;KA�.�H_�ST���[���I'�yD������]8�N��Z�k^�z�p�C�D��a�)d*�z2��]��[3!1�u�;|��OG��Oٚ��G���Ց���ӝ��p���J�8zRi��:/ �R��ZjKK'�,�pSu��R�U8��=�7,�A!�n�h��NЄ���aC֕_��bx��=DI���9���I�i3�C�,�����{�ʷ[�N�(Y[�:qRӰ�7��l������X:���Ǎ	�f���(��;*�� �s��;����nX�qv��mii)�_e�8'Ȩ Ȥr�ut@Ъ��=��ʹ�O�s���&��'��a�Jc��<��Br?�GF�}��Q�������OA�_k�{>q_�~���E���k��:������~L����h]z�|���S4a�vLd6��������O���Фn�cm�#��(��ɞ�g��I/�u�Ј�A��/�o���-J�ż��b�8T�����f6��i̚�X��o�`^1S�<y���",hSEL2kj8:t��헗�Ar2E7i��kP�[� ;��R�~eո'1��"^OA���@lr_��t,晳��ҍ+���^@̾�  b�3<_��]LW�>m�6-Y�M�[[Ce#++F�Ƕ���b��Syp�ug�
�%�=�x�ֽ�*�R��i"3�c�fryu��$�i&�{��U*��Ll��+���	�����t�:��x9̳� o���oW�g�6�SՄ�����.Y��Uק�������O:`E�Ĉ��I�A��Lx;�-�(��k���Q��s�	��Ɋ¬D�0t��
-(2����{x�e��|��wQ���rq�.P���۠��(��C��999rI��tBc'뜮�����`�yo=������dtuIbLv�*��L�`�h-(�N����p�QN�j�ݱI��4��T�x�hվ��_�����}�ɍ�$������3�e��i�M}��̗�A�Wܣ0�Г��<�KeSP+��|`�Jـ�ݧ���_1�j1!x�����a��Y ��À[�X��F]ഉ9��J}�Pt��ixr�_P�~��+�� u_�
i#s��w��%����s�`�[?�������\,��>�2��1*�Fmb���]�#�8�l��k3��|��I�ҹP�qt��ΫSjAߢ��L��MQ?�n��9X;���8v���N4�hW���w�"i�M0Wqƌ���)�qq��@@A�H�i�c2U �͆Y)�?::�y�]�9�R헞��2����H��(dY���7Ϥ�/xsI���?��ɡ�.0�N,��?Wp�d�:��42.vܛ&p.�[<��@��})j�[!P��~Ɩ��Q�q�@�P�y�a."�3�c�K�����-b��b��'s�ltK�C��s���l��͒��7pA��M� ���~��d����^%f��w5��t�1W�'G�4dR�0ͯ���e�lZqJ
�H�o߾��ȵ���O�?9�֤�^ߝ�{~��DI��#�:��cf�4\?�*���ɞr��b��r�c�-;h���g ���@E*�T��cS���� _��U���&��7���,�2�S��ZXh��x�?|?QzCNHb���G۾h0����H������1��?d5g.�7���F�?���Q��w*�or�|���{�/��z���\(֧�NӇ�O����o;�f�I�c�ݶ�rЫ_$>�:��B��Ю���R�0�>������|�R~1i�v��������tH]�S���t7"\J�����A���C�I�������{����眽�^{�3w���e����-8��8��_�C�F�X��m��˰W�w3w��Jڪ��z`8��͵��G�šV.���Jc��xm"ȿ'�~B��!E-�"jk����W��+�5�D������*��y�P
���1����H@+�H�m[����!uS?B��?_�tp0��Pڅ ��d�Y����{H����,1;�oµ
h�A���-���t���1YR��,��g�e}"=��<����>=����^@���d��DW�2J��-�}�����\�o���e�`�����N[ƽ�\N�R�_D2&���3͹Έ�Ӳ�|�������MRi���\�z2�e��(�F�B�?���FTyT�n�삤��0�����2�JB#_ ���v��nߟ�{���ÝA�Ÿg����;:�����/�`R�����W��U ��[.���I��`�tŰ'�s3��[����n!��}~�V%����O3ޖ>)�����C}?��B��q8߻�C�{�%��Dq$֍��Zy�b�w��A���arO�Ӫ���eM����76�����h�vv�\�)��ȼN��%X���2�*Ex�c{�@���
ew�Aw�UdG�"�Q^I�2��b�e=3#CFAa��l��]�g�Y���[��{&��s��:�h��:J2	=�xU���vS"��껟j�6���N~�?�Sr��k�e-ә.e�s��&h6��i��%�k8���8��E�Q\R|X�[�˴z���;�*�������A��;���S�j��F��&z�,)a��j1	� 1�\ZZ�	4�#� �`�xP�}|s�&q?9�uP%����ۙ#�����=�i��"k�j�DG;)S�F��ӽF�������)N�������'!l��nBOu��3Js�?$����%��i%���X(E���ZVK�x�t�r�752;�0�ۤG���|t͞/�zs���kx�M��ƖB���+m�8�>V�;�%!1��~vc��U�U��ێ�[n���I����T�t���?�M�*)\G�	�o
3c�h���84aR��ʌ�wR�dw����>	{�%��X��������e��z���[u���.J��W2�s!6R��@�1i�	��)��*i�q������j��d:�.�$�1Յ�5�x�"Ump,�w��y������`ҌA��բ��6z����� �H�Y��[�s�F'���B����T@� ��~�l��oV�C�u��Q7k��q�vtd�G@�ՙ�ݲH��/acS��Ч>�]_b�N-���0�e�$���*�>\�gʻ�i�Wv�HJ4��3��WGHuc��u`N��w��}BҼ���c|-�ૅKG�U�+�D�A�I,�����)8�hl)e?g�E�zη`���	�3NU'gfz��2��O�3k��b�5Wk�w�J������L�t���D�S���%R���0p�TU�~f���&����@��%)kF���/m�xoŏv�g����}E�׊�A}R)���W�9���:˃Gw����9X˚i�Z�ݐ=?xِ=�K���Ԯ9.��E̹��jg���.<��������r*�럟[?����&&T��fԙ5h���qxa��ז�^�V=I
Rƴ-�g�0�����E������.�{q�5@�5�fw�m��0��Y؋ &���X��bI��6^����n���ꭒ����j+2&Y�Y� ���4�������m��`b�{�=��_H��fz]^��ݴ>��K��`�[���0c��Y���mo��E���u�{qZ��*���O8�:����?ma��B;�1�^�!�T�pE��c�G��t�k7�F��Z����`�+-��~%����Y|���^Q���O:VVŽs��C�fwLr!�۔�����o3�(��rZ��p��ۺՌAfuֺA��z���i
7 +a Z4+�H`���^��c-=�7Wa9mw�B����U�=�e�+ã��W�u�#�O��W�n~�������"GIgZ_�D�t�<F�9��}'ݤz2�۲��a�Κ?yT�A�M��jdD���RN�fl�%!R���<�P���
�]�!i�c�l�	����U��T��5�v>�V�R�)�5#F�}���N������@m9������r��^�`�[�9"W����c�lq%y,ںɭ]�ޟ6��s��e�2-�'7̍��#�Y�ZB��;Ы�6��M7׾ �|�b�W������j]�ܘ�H>t��
9��E*c����f�r��2^�N�t����g�O�D��yK�V�����t�`����ի���'�4iiy�K�Zs���;
Y��N�������j�IK�����N�^�{� &Z�BSSSe�{�W��?U:G�s�U
��/]Yt���l��ܯhӳuԋgÖ��:9q���+��l��\1�:W���z�x�}��* �?�}Ê��6��#�����4�{�Ib�1f���2���X!�X���Ցdg҄ԩںS*�MǟD��4�w	�xQQQ,,]ק�
��#l>tCy��L�-�$�upbۣ���F���wĪ}��}n��tEs�ŭ���0i���?�vSW�t�D�<{#l�W�c!��{�_p���<��M�5A|ʷ�����(R�7��bBX#�+p�M���y�lu_���±*�V�aҧƾ#}�I�-+GnȼY�L��zWU�g����?.���Q>Xh���pZ����}��uܥc`f��{#���4t|:t�k�ɟ�=�����^�C��4a��K7��bݖ�A�v��t�U{��r�wqz �X�$�A�<�F����ܖ��sunl#����\Q�� ��;��a���|���H���پ�$q2���6��X�����
*��\Kk	qq�%v,g���0��>�CO��4�lg��7�~��ѩ3�>��pd��i�xT4���k()��p��Qځ���Ԙ������h�i��cH�&L4���h�R�H�Ѵе�����L����s?^�[����xt
���O��4b0n`[�ޔ��B������B�U���/5�Yn!�'d�=���7L�ӆ�����v�Nb�J"ߛ����}���e8�{<��Z; �0�8 �{��j�� 6�����[éa�<�i7ϐ��M�`i�:ðև�� ːL�S�����<���e��R/447i�
�E菕�u}��|��h���Q��H��`b?�*��
G;aO<R^뮡��l�pl��G�Q~�%2 d��&�AU��e:�?���/�º�́6�MM���坓�C	�	�]����j�]���M,r��z5��.
��Fv�i<�mЫ�joP�#�ON��'��:]wpxD�^�}N�z��)yT�jE_��j��G�(�4BÑ���>��x�T�3Ģ��T0v#�;]=Q���_�x&����4&������%�D8:�.2y��Q<����_���Q�����}���a�#+�/�?�+Gl���u6<������jƸ[�ylf���8�+�w��jj�&z�Jz�Ovx����bE��t��Nt�cw�$�������9~��E��b��F{����;� �\.��3�+�% d��ȍ��]|�h��w�&K�7|��H2�����"���*}�)���t��;�֫%��:6ߩ���j��{D��E7N��.Ӧz=(�H�UUq9l�<{�Z?"=!�[|y��
 Lnv�[/6r��../����6��B�!��.[�bOa(�Q��fR���t�[���ᮙ�&��_��g�?���3Y�J��v����c�<��\��}6��P�V����Q{W��^A�X�����pg�kH���P��(KZ+̡�!1����b�C�F� r�sǫ��]J�������Յ~o$\Gv��8J�����=LJ�����}�{-��Aȕ�K�\��؜����@����GbN�\�}k6������a&��C���,J�`��%)IIɁ������cIU3$�0]����(�w/D
�U��l>�Xݦ{�h;;���e�k}$5=alP�?2ש�lܷ?�������J�����Pq�F|����-����6<l�N�jAF���	��6@)�9�ܶ���߃��{�7Ʈ�1�~��?7?-;o2E�C��_?5P�%�%v�_^;m+^\8��|$~��Ș�N��_��=@0�K��J�V��<�����4�:
ማ�-���d��4�.�H+�%�:_�*����(a�  f�+C0T��侊Q�]��gw�n��;y�W�<��@)�MԴ�ɼYN�Q������;N>��t��f+ō�7ɱ�ha��vS?j��`_gD�����l��f6�����}��"@�6�f�7x�n���.H���kZ\�w>ę������$���h*���o.V�i��GL9nU�@���O��P[�cn��e=)@j�[ւ��Uf�r�"W3��P3��9��hf}��5����A0_HH9|���������+�%|��УG���K�C&�Mb� �#��#c>=�3��{�NԨ�j��<���púh�:j�O[N揩K���.6a����*c~�3w^^^����o�^����|��O*�� �_6�vm�x�3/�I�����s��mQN���/���㼼�y���T4���>6%��&͔��C(�Մ+�5X�^!UVS?]�uC#D��2�)������ē�^#�1����t7�՚�x�7��ps"�ɋ��p'�����1d��g�N��������9���R.T��,�0e�t8��7r��藟N���:K،��y>G29E��Vk7�N�sv]�L�8�L����b��TGh�:�I%��
��q���Nh��_`��"DY�(++G��j϶��Ul�u�]�ox�N�������������AUm����B�P�XN��2{��K�n�dx?���eK+�N@#�O��/֮��r�X��	��9����ڼ� O6i���`c����2@�^�8���H����y O*�g0w�@�m�v�Q�a�%�D{hF�^c����;H	V�A�*�Y"n&���tA׹��]���Z��W�����6�ׇyݲE>� T�FQ�{��4펊f�(����M�Я_��%��^��e�RR��������R�-��������2v+׵rOޒe!%�n��ނW#YZ���'^H�(�I���}%_�=�]��%��㝝���5|�C��**�'�l��/)��k���X���`6���2o�ɷ�[�6�,$�2�������}W0*.DK�����$O�֣c��ٖR���&ڢy6�\L��~�m�م[~�������%%�����6s��pW[[f�L,������Н
f�4���\��?4��6/���_t+��3��W����B3ݜ=�ʞ��l�L',0�:�h���'K�B�fA�ϊE=/j�EhU���O�l��[�@����ܿ�~Z�<E �U툦��q���͍w�L/�sD��k��YH�^F��h�7m�Ƙ~�?�F�P��z��q>�k��t��Q�c
�P��*Q��5��~���W	vx��O��Y�67GކzN��!c?���-,X���oښ�ZT��O8w���3��Yc��qxxx�ƉЬ�H{X�֨������䒿�=�Y�_n�<��:<=�K�.���T\�۾ɌM���'�HG��f!��lH,��T�������é`���`�/0S�C��$ ��6�:mPH�1��x8+w3[���@	�8� �Zկo���4}N���;���k�ԍ��ֆ��	�,V!S�3������7h�@��&��/���t4̵��@�@�|�w�I	��l�[a`����ˍ�dk�#
���(��;f�� �����y�xˢ_�r|�ջ6� ��W�#�i����ۡ��tv����X� /�(R�e�jA��~�Ύ�=��E�W�qPӯF2�L���ʜ:.�k,�|������=�.wLjɫ�zՒ4�/��a�Y`�RQW���/8�}��3�T�W6^]\[Y��潖,& ��B�bt
o�*���xxys[��t")�8�7��b��c�닏�5�j� �s�*��lSe>C�'����iűi�@�Z����-l�M;����)� Û��f+|(���4��u!5��γ\�<��yW��ϻ�/��: �2��z��Yt��?,WS�%^�fy������@%?ر�J	Zw�2���G�#"�u��b�p�5�T 1U��/�����jlߞ�,��~,����x~���qJ��n�p���7�o{>�^��
,ыX�ӆTV���s'�$4@�b�u̪��XFOo1�+==]��۵�4l�<Dh�|Ȫ�iõ9�.�n�3�t�\�Ю��zW9����؈C��ȓ�<β�<�R���5EXYm)��OO��^���4�?6���>��o�rp�3"�U��c��\C��`(5*���JA��+��M�N[#�k����䘞u�N��`�u��.븰}[����e��Nm�;��_�������m�����z�I:_�� 2������Đ�b�#?7�=R�{>��j�ב��I�����e;@�3���%G�&a6��.��&�8��r����{$������י~���]�W���ɺ�Z���t�
%�%������a��8��ä�����3��}H�i)���i��� �4��D �n7___��Tb�*��~�.����=%Q����ϔ��?���%�4[�ٱ%��" �0����t�,�ֳ�C\ݪ�,������U�l����O�NJ�2k�����p���.ߩ��{�RBK��'] ���[�ڏEՐ6h�~'���֖�p4��4볩�w�*�|h�՜݊P꫿���r�p���~ш�rx{󍅈�l����%[����KKK�Q��ƀZS�Դ��ef��X1O��HJÜ�l(Vo||):�Ѻ�����}�\e���D�����ѳ�[���%��#ݣ|����q��6��
$�	����Z��Be"^۴]�4�@=����x�	��߱j������	 �����l�#�m�C�q����xc����H}����j��U_��v�+-�Sa����H��q��&�����;��g��a�k�WO<�Xm݇2@p��*��O �?�t�
�
�����`Ij�څ�?��8P�/&��V�Z���}w��w�j��� ��S�
�S����Pf[D�'͢�
ˋ�#�<���q����^�䉫�>�����l��/�;o��x϶�fx���0;��Cѝ4Sgh��	�߻T[�:E��b��z���WA��J����Gxi�K0�}Ǣ_��e�f���RG|����n�jOTgn�����*��L��W3���,���ƦW��M��j6Hm�������v���k?�{\}�S��^�����1-��1���srhX��Q��5�"H��1X =YpE�(X�;��뷨��/s0U�F�7����S��l0��F�������h� /]�לoQ
��|w��pL窽��̲�p��#��;ѻ]��*�w�k�]�c'	�hP�K�n(3�_����#F�e�q�%9����'uzUsY���Vi�Q�ّϳ��k8\����Ϻ�/KW����G��9�[u��jC�����7��*s�G`�S_/�1��p���qD߫ۘ����|�ǋgW�G�|#)�V��"��ټ=9qR�	)�s*j(�(v��$���.�|���C&��U���<����S:�J��b� b����5�;DV����e5;x�]�}~r�Yk�-�2���g'p�a�GF"n6h�u��q<��\f3����.d�� �(�����!�V�{�k�P�h� �7���'�g�����U��-^[++��'�y7���0��3�N1��TAt�Ej؄���"(eR(���8���dB_�0�#3'.���T�s�a�ߴ��X�x�:92u�:\��[��yT� y`P0��D�#W ��ۡ��2YV��^�𲖪c�a���C�
�}��XÕ���#��U��������(�i
R���?���6����6W�.'��ȁY�~��*�_��$������o�m��M+0QH.�9�${�p�� �,kw�D:8�"�
ׂg��Қ8��t��#��nu�K�	_1R	��`���!�&��4��������z�u��r��%
�%F�V��&�	����[����\zA������g�F����:s��=$��*�-q#/�S�)���m�mR8x�ܗ��a1=�+�^�!�6-�p
Z8ȝ����Ht��˧�N���2�l������q2u	8���e���{��R4�	0��B�EA ���'i`q4����Ӧ��Wi������7�2�t��zڠK� u�3�2�0g�FtP:H�2����ߣ����w�IiD�	h5�d�E�Y#��FQ�O� 3�ƿI�<3��i�pl͉rO,���l(©�F֝�z����u���������g(}��H�	�B1|T.GC�ޘV�s$��e�a�+���w�4��ظ�v��/��ϭ^1�9eD�Mx��7ެ��G,�EjB��|r��H� \�Ϻ�����j:��܍M����>��7���(n��/�l�a��s��1u�Y��\��`~��뷃�O��#A��Β�%����5^qi�ɺZ(ziۄ�~��C�SR�^����U�\��I��<pK)��A������O�
J�[�j_����o�O���?��8,�5@��b�������0�7���0���>MT׼��hg�m��rB�Ѫ�4���|E]�8�0�y���	�d���A��(<]m(>^�3F?$	*N^<���NVE������bJ�:��B[$��ğ�G�K� I�Q]�@lo���~QL�p��K��=M�&$l�Y�z]0���k�RJ���� |k~B�x�� �y��C�Ba�Op���h$�_Lt�t������(]>mdb�	�w	c��DȂ@����]K �WP},U���������t��l��P� ����%�6	�X��i]�>�e$H�T�CQ�h_�ˡ�����[+ex:��,��kq��#�tE+v���z~le��'>�A�-{���C��n�I�D�<�`K(v��k��͸��隓%VW�0(��
���'�-�ɴ��oّY���*��9ZA�z#`O�VG(��}$5��!5�~�'�+j@�-,����v���Q׶�:J�>�Bm�#�^1���Ԛӑ*n��-U�emw+*ċ�l��L)�bE�>�.^P۶y2@��;8�֏'���&��sד�Eߩ�O���d�5�t@��~�B%XZ�pӆ��?��vRQ�5��(��:���U�8J�x+v�O[h����V�:�"��[�ˣ�3#b�P�+.4!~n��xt���CP��,A&.�ʥUZ8c�|j�h�~l@>o���W�"�a�
|�&@��0RG�Li�l;\+��;�[���z��Ci��e��5�Ƹ�N�/WdX(�L�l�Bw��f���=�m���Q'�h��Lp>���;����z���4��զ)�SG�êv�x2CY�*��w�P���QG���\��ty��u*�7�s�;�O����U�/J�0(���������G��9�WO�D��.�H2����u�v��0�r�@,�u�{f�4�O�w-U���y ��zy�{&h�n���j���k�{$�5NT7Nkh��4��5�WETt����P��yr�7�
����3]M��%���󮫴7�L�ғ������H���ۻ���"�V�l���J3�v(��&���"��q
����n��7"��-����l��O���V�����GrhBYKŨ٩�����4TF��^ �iB���+ili�`��ͮ���H~�Z�VBqpY�I�u� nV4�XSlG$L��3���;ݮ���H��܊H�J5P3��?�"���Kt�`BF�
3!�߂�搋�3Apvm��L����)l��J	��)
C2a[�J�h�Xa�|J�Ǳ"�?@��YΦ�[�|��M�̳4�G\�s�����@���zz1p��U���Ԧ(V�-��;*��F�*�y���z=�@<}�����ƙ�!T-�v�j�� A�i�&�w�8��.�ʦ�@���N}hZ���`�`2��I0��5�Q��#�`�X�p4�� ѷ2>G�	?ƅD���T��0y����=~S��+�n;�m����j��^ )r��r'[�'W�Z�%����4��m�"n��%$
X�� Hgd��x�\�Ƹ5'CO�U�n�"����.���)�YKGUq�!�@0����8��YWK��#���4�	=�����NK��s�:����� �"e.g
���LYL��JT���O@���vGV,���{��W�w���TGM�5��o��п�Z.���2cYV�!g9(���G1���Lԣ�T]�q`��L@"Y���P#�}��G��=�]>彣���l5"�I't�PZ�ٯ���ƽ�$o�I�o.�JH�?�<�&���yqw-����ÿ�'�}�E9��~�5�g�U����_�smv<W+,m+l�5RW����`Z{��qkT ӓ4�es��#�y�VF�do��b/���ۋ£��\][��=lW�U�b F��"R\d�'�5A���	V�j���ܱs��+��]����3�o�BJ�)�mI\�:\�&˹��;�-w] Ê�'&p��ـ1 U������	�T"���Ԭ�2��>t�;�@��#̛^���{��LD�2P��_���P�����Wv��J��A�,���d�4��u`��a ��Y;벽�~�@�����l_��9�.���x@t@M���f��X.�$����~�'���A*z(㣒��e/��K�Z������%�eW�B�����>��4� ���6���E�	����P�4$�.Y��z.��;ѻ1,���膉�e��~�#���\�E��'s�d���=}�OX� �lAWq�˻l�a�.��G��!�a�؋q��W��c��6jq���b���#��b���_� 1�l?DJ3��xR�f�4J���v	��Ct:�['3���[=n8UHf��e�5�V��'Ҽ��4j�'R�^�Z���ȉ�YI�Y�HD�=��$r��b���բN�}��T7f[9��= q��t@�!k��}�U���^�����S�5�Ǯ�0h�������k�k�`�@<=�xQ��0��ƶ�l]�Ȗ�e��i0@d�n����z3*j�x��= Lv�L�����D����}}w�` �ˠ��0���.�P�./�a�(/��(Dۛ8��_ ��+4Y���w���0�^����*�X���VׅZ!�[e���JXe�`���
i2z��j3ļ?��k;&V��h�	��Z.J�{�����z��#a��E�YI�0�pXc�~��c|RF��݂T��f�5�sr��,�GB�Ǐ\�Z���Բ��}e1g�3,[��*w'�EE4X����Vb�Ezh�Î#�ߛ��h�����p��"�x���B(�ZV*k�Á��HGܖ���,�HC
�-|g�}���ۿ'Uh���䭸�3@�m�N�)�JC��%A��"�����]n��UELL��(�H6x�'�3�Ą`��>j��<��%����wC� ŭ�ItA �2�R;֍�0���A �n���N�00���Oݓ���oL�����'IJcM�W��f �D��Y�����v}�Zw��4ZS��(��F%i���uXR��/-a'ט9�0�Q -H����G����<�
sL�W4���UV2sR�R���<���j�!�R�d{U�jt�}���>���JM�k�ǐ�Y���uW�� L���M����!磡//�."瑁���
�K���Uv$J�0�*6���y��y��(�?%��q�/aD�O�y,eW����{�P-�� %��� *����(-�{K	2��/6���L
7$K�̵_�#<� ��"��Ֆ�t$��+~!�Wt>��r��\ja)f'P�C�ӀN�bT�	[��D�0�3&���5�����V�f��Gx�6B�5�)+[��g����?���c�£��.a!�`c�#��Ϝ��d�b?����j`������^���/	�^p�&�
��>0j���M9򜗘��� �a�o��������}	�ʔ����%�p���D����7�ŏq[��-�()�Y�|@��Xh�d�-��u=,�'-N�#�B��@%eE͈G�:�s�p3pb��9���L��|��{2y�Cb]^��'����	�|me<���i�������#a :8W�����w�_��u$|�f#�>�y0�s�(�9��;�H�d���y�����f�=)�����\_�,e���Z�@��NX�_�<�r�l`)x�Q�k���1ZҀ7�#����B.Ed)bp��B�]��%�(���yK�6}��/�o��m`д&O_maqm�l�����-�)�⵴3�����T�<��:���5�8���V�b�4(O��8s{)p�.^�E/$:�0T�Ƌ�����}!�#��ER\�p���vऀmʐ�J�ԋW�H����c��Ivpz�7.j�)�4��;nl����<#ۧ:B���O��/�|�&��A��NS4����׾����*��5��ߣ@�ZU���3�;�[8�c�}�V,���R�|	M����U��[��0@h|��}#�>E-���'R0��=�CI<.����[� ��|y��e~p&�nz=�Ǉ�����C�>0�����ۊf�.B��x��n�l�侹t���q���,7=F���ק��� ̰��m  d�|ݲ����%����z{fE3 9Lsx煘��������v�*��˨ ��<�7�>�C&nՁ5� ar�@(��a�Q�K��G�k��<����#�%P�Q���}i���#����ca���������%\���r����\O�b�6�󻷵3a^��EV?[@���J �#ܞ�0�B��a�(�(Q��n`m�Wwԯq��ل(b�&
	`c��(._����8t��`/~��m��1\&wg"0��3��͍}Û4�"�J��U��Xʱ�4u���8Y�vCP�l�2�P�&
H�"Y����{��Q��p	[�{��q5Q�(���~���\\\��:w���a���w~/1��	�� NG	�̵�y�J"� 	��K���@v'�?�"��D�J�SL�J���L� 20�vC��X{��a�	�!XOn��{`���8�D���A&���������һu`�;��m� q �����'�4���d�����Q�������#�<�x-t�+j�ut�=�h��37e�]�QT�	u J�������o�f������T(�X6�'r�*�b��}X;�@]�r����]����P�L�j�����}�Ѹ���1��ZQ�c4{ip+uy}:(А=����^�+�����sűa巧B��څ�}�V7ԅ��PO��-�|[)�-���1���YEE�j7F!�䲔��TMX;U�5�g�k�r�[m8γamZv8��Ȅ$��=�_���y�.�`�]����p)��J+�\�a)s;vK@��784����{��e����U���~-5�P��8�p�� R,�#�'}�(9~�=�� �P��`
@�#a?YːܯE�x�[$��{D�i!L]�7ֱ�=KЖB��9�;a~�5BP{=	!L�{]���5��'��S�R)+]�&�L���9�����z�YeJ]EȆѨ��1���Y�p#�ǡ��u\�e�ץ}�7S�|;�H(F�O�%Bô�Ko�Ŵ�mh�R�X�_��d	��tuvu}�p�%��~qy�6[i�@c�9����f;й5���wB3q��7�\�
�t*'K�	�B��"��2�Eӈ]r�RT������}n��E�	�\����36��^�p;ۅ�*Cpm-p�Bɔ�\$��s���X���s��E��&ȁy���5�u��;GG2:::�g�['f*����G=����{������ʍM��O��C322���s�566�MO���H1L-ûL��G���6�m�cT" SЯ�~�ƶ냖_퇱��˱H��An��,Y^�E�y5u: �Y�����:�Ņ��vFQXX���@��}
�e@�Z�1�&X���ż�Џ�� .���Q���#;�47�3�cS�sW�ۉ�;9'�Ϸ�� �@����H�'n϶�9�[��
x�F"@�|������{ֺ��E�A�ք�k�4 G<:�̀v*m����غ���C�RZ8E���MTShэ�$�a�5V�	��i���qX�QummN]/������K_�����|�hp8��Ř�vf�	��|2�H� ��u'���-��Տ�^d@%�1��Z������XYY��e/ܧ�y׽�� �S�}�z��N�f�L�3��COOo���ϝ#�ZX"��~Rm��S.V��u�wH�ߔ<ȼ ��>�9z�j��c��a��9~�f��	�ą������{[M�0ft�_C&  ����W8���=�>�¸�@�oXJu�X1���Kzyyɥ>��k�����daRԛ�ᥐ���[b��/b���U{�� �⬷��?G�5�T��`�q>Т���9;;'S�$�[1�����ȅ�Hihh�*�$��r�ڙx٣�n4�d<�����f���Ǒ����a~����7t�B"����s�&J�@����Z��6땐=?��ԧ�$×(>�z2�U �&:���aU�~%����0l�����M��' 4�����|�?��1��ٗ���~^SP���3/��0���J�@���n;�J�=�+3�:1!��ǫy����|���I
��d��%Y��}�pqq��;�s���}��;�Q�3\��v�{�D_`�ɓ��ܼ��M��rHT'�k�ʍ�\c�������4t`�����6��r��fCt���Ո%�v���2$2I5�8�~%o�����h�f�����vŚSq���~Hq�@�9�i:|͉D�P�[Hʱ|f9ί�̙&�G3/��	�e!%�XL[�KG���i/P/�X��Es�A� ��6Ns�gT��VT�ሜ�l3��BMLg�]z�Ǆq,MWݵ�s�6o�*�HU閼4�-wO <2�bƈ��,�J/.��q��nD�N��,��j��#�Ԓ��EZ�HN4�rĨO�!go�%��y���H%%�6�}˪�"�6�)U�s�k!�@m4��l�A|^ҷ��Aϊ�V����|M|z��K��8�ė�ؓ�j6&�N�mL�LZ�]�h��?<��)~�x���^K�ΐr���`�q�>��+�@m3�|v����\M�̀�b���O�V$B���7���C�kWLQ���$Ԋ`�~j.�!�#֬��Rw��`����衯mVC�G8����oƲ!(@��>w��v�3"<u���0u��F��:?�x��p��R��E q/�3�\�5���˲�~#����P�g�5}����~NL�0I�9Pu�ҫ���e�&$&�����4���LS[@�y�AH�Y�?�p��x�H��ok(Q``�5vs�<�-������ݏ���ٯw��"6�Yg��p� ����aw�\+#�5a��)�6$Fm�g��,m��a5<Q�[@�nC��=l���N$Z����#�
��Խ�{��䵫
��c�����s��H�B|�Z=�bh_�(9�K�3��n0�����im�$�d>s!�IP���9�u+4ǣ�������>c��Y��\	t����[�[���	�c�|p!{,��"|���0���f�@��Ɯ<���\�F�Lf��O�����t蕧�g���2@7�b��z��9>j_�wJ1/"�1;ȼZ%��FSd��1������a��#Ȟ���i37l"jٟ���k�(%*�h�A0ً��`������7�g!�F�s�U�������R/��3
aM����7�p�}���P*�����5����pt o�H]����K�����_cMr�w�{�L,.��v�\?���7��!N�w��)3�rU?D�$6���Ek�q�=��3�V�Lj����tz����B����gl[�D�����-�#�'�3'��F�M7y���] }��w+h��*��Cz�l�ȫ��4��l��V�����`\���-����g���1R4�eB��C����p�N#q�sOpR�� >L-W0ȥ��_:������D����ز_����;���,�
q�t�Gڪ��6�@�g�j�1��|>�A?�.�4#�wk'o
�����=�#؆g�����r#�~�mgƻ�e
C2א�?�$�b�^3����D/�����x��,�{���d�,����L颇��T��p�鏜@"X�fb�U�|�5ݽ6�-��c���BIIik��9�)��W�k�^��W�C	��4v?"��}��7M\��w�Ɨ�2�l��:���+sZq�������ĉ�@���l�Ǹ���ͺ�|.p��w�(�l�Bv�l�!{r�H�Lr8�6��0�����q��c��a���������x�f��Ә 6��Q�5z�(���#��(ů+q&�ָ@vR�b���\�ҟ��ƌ��|�0�.Q7^�{���(2H�x��ن�H6�5�eh��Pžܨ2��n�4�ZD�98���>�ON����Ѓ�P9z)��+����C 7�N�`vq��o�a��M���O���RÑW��A�����z {%L���A�iv��5���,Z*�^�>uuN�U��iA ���*���/j������~�z�)�A����t4�.4�bb��du��6��x���k�"#�1g�8<i~<l��ѝ&~����ꫣ�z�v�n�a���cBDP��CB��;D@DZE�k@�n)���N���w׷�]k�������{�	�й��W�y� ��:M���'[�@@h��8Z��c���.ڟA�4����.D#�y�=�7-qo!lFW.���n���neh��Ț����|I�IH�y=��]Aei�1�v���r`�3GWc|y�,��j���4�70H�v*M~��
�%��8�
}j<�p��9y�U⨴�Y!���A�`�IKECC~�B\��^�*��j.hu����jD��e�҃��|!��ou��5��I�����i�y?|Q
sX��mw�� g�s����Xv���1�P���kO��R�|��9_��\FM���Ѳq�K�)�Ѽ'`kzjٗ[~�u���8�!\N��B�~����{/TOwH˂�2�BC�'0��P��Ki�$]�ͭ҃=A����\�g�{��A.ft�	����	my��6Y j��W`F�v���G��-Y0���19�W��;�wi���Ţ���g�v
|���焼����hI��鮕*��&��4ՙ�q�Ȭ��;���t�'f�38���b�&��y��B+	�L���hc
���KR��4�31[��F��ihC��2��y����I�
a l��xa�{4��  �����G��A��������' T��$���x.�LH"�2r}����=g&�~�C٭��p����D��E��-aYJ6.��n��G�K0$eپ2��@����ٿ<�����$@3�~8��zv�=�T-xc�l�_���w m	h�Ȁ�VG5�B�9g~i�� ƀ�Һ}k�,��wXety��xbhB�u��5�ʵ	�[`]K��� ��[�%�={�u~����[�%�H5���`�+ e'cW�,8�>���?Y�z�n��+>�L���6+��Q�*���R����3��7J�9ˇ��=4%;h\&ig���gY�ՋG�?��ˤW(.�m��y�#�n�!�������`+�S���K�k���"��C/����Iq�ił�p(U�H�;��wi�jL^:굈�C+UB(%b��z�!!���a�A�4ˎ�"�5��\4����PJ��������6��x��0Ⱥ k�;��%�WL@�eg�a��a����%+
�[}�j�u�qʹ&�~�+��>�A��Wd��O����������-;���}���ղS����ؿ��m0�*�4��eE���>`6�7�c��������x/�G����3�/^���s�7�!>/��th劳2�Uf�
�X�H�Ѐ���`�"�c�Y줰��?�l���.A�=���7���u�&foU��C�*
l��JQ��y��{t~zN9�#���1k�E�6V�D#�<�����?2�Ɂ� �(�Ι��m�Cޗ��XX�ڋ�2��!��+.�z���w@c)1��μ\F繰�C+$��Ze��X���𷴍��yQ���{�B���h�K�'��M.+4V�g��	yﾳ�{���^��~	!������>���u*�[�	o &"J���{�[y1J8a��Lw�O���.��Ek$cI����;Z���Ag��t#9�@��U�HZ�̕q$?k�c]#�@�i���U����K �u���7T��>Ŭ����$�|��p�31�y�v��6],�V��(�=j��!1Q��BW��5�yk�!v���j���4 A?�����أ+��������D�}��S�9q&.Boz3�6f� Cm����N�(��;��R#L>�hB�Lc9����b '�+.܄�$�`��-oq9ǳZ_W*;CT�b_��P�}�`�߻R�������yӮEլ�>�u��R(|֭Å��(+�p�u�f�����)uA�Ǻ4>�z�[a	@��h���%�GHD]�0�R��G��s�����Z4D�_�$���E��խ�VT��H~�81p�z�Ll��H5S���W:���}$�!* >�}`�����x�
�-�rV���ſ2��;$C���$���C�@5N~�CnOPe��\�{��%c��qS'!���һ��Q��3ς����S��R���t��9�
/!�xiʕ5���I ��<�B <(㎂�if^}t& Z8[����S.@��E��pn`�wl�=�E�&K��9���㒃��1�w���T�}��QS,�"8��3a�9ˠb��.Z|�,�j���
q�6����k�u���`��O�s_�g׀dY�c���;���WFuP�ly����š��C��E'�O�SVg�3ڶhB����1ЮzJX���PHwT���;Q����~y��pk,��*�3�X��6D�$L9ǧ�V3ն7�	 ։��O9�G�3�k|>�	�g_��Y�z���������l��l��X�g�	ܙ���RG�N.	��
��6pZ��Z��nm�@%�(!b	����A���4�Ī��a�¥��"�QP�[����*ۡZ"١z�x�I�A2��ϛ@(-O֛�!dgL���N �Xbv���i�vR���w�B�&�3T���e�s����*4�g���bC�b5���Ĭ��� L��2EV���ީ?���\����L��yzci�b �<�EQ �ŚE�>���xA����Q��!g�������$L���_8#	g)��T�T�aK�����#)UB�MP���@uJ�7�?�h��E�w�}"Bun��z��]S���������N�-YY�7n�p�	���A�K�C0�0&v6V(*C#����{iq�������<�j�a���S��I��RxS/�������j�I7�ي��.�L�}��%��z,�Wj�a��cv�����a*T����
C��gB� Ŋ�r���c�)�I<E�޶Y���1�^� ВN)P��� ��Ys���NB�`� 9Q$��=��\V�$}��oQ+����1�"@R��s�Q�=�D<�^e�~��;����^k��Z��;q:F�®�rl���6�P&��W�oCp�m<����Fg)���aI�� yG3D�,��8�����,�����SkR̮K�ޤ���#9ʄ���0|-�������ٖ��_h��V7���a�W	�7��K��eW�t�P��(/� �Ob��?��iB��e8�U�vK�1�sq\SIO�hS<Y��o
8�����X����fjhT�Z�(�#I�l�J>>毙�����ep�/T�4��P���,U���f�͟[C���IQi��W�.��E�FI��C�2��'�7�y�0�1�%\��ߥ�W�p��hM2Y�)e�3��
K� ��ao/Y��B��8����Hk�+�M�8=g�T�'�1ә��4��D��%�4��i�,�+�W׋5����Aخ%ڦ��&�lDZ(iu���ۅ/_����}��|��,�\Ql�-x)-0�_j�T�Eq�3\A�4>?&.TT��z ��WT����ON���k�5�>O��}^����iFJ�eξ����5��ڔ���t���;	�������&���mJf�V��� �y��\O�o?w�PG>e޸u�n�[jNh���JI~�˷U/�U�<�Z�����/J��紧�x	��*�)3���Ya%	Ơ�+�C��D/e���7Ss�Ǿ��%�ؘ䒆�����V��e�+z��0�#��gKdNw&�X�?�T���޼G0'���a��5�	��	[���BO��24�>�uP����Y�I\D�܅�^���D����>EO���s�� K���h\ϐk?��q���l��, ���H���%����z�k�ސҽeE{���8���h`=���Y�4'�	&;=ﱪ.Q��J�F��U�ZqH6%�i�6&�|�g�.�m����p�y:�D���������т�GN#k^'Z�%Ӎ�}��lJ�Mmؑ��� C�_�A�.����f��I����gw@۱��yb�����%��_"e�Ru�}M�~a#�G���CQk���戓�t���|�X�
��]�8����vXX�{�RO�(eo�*s�n��g�%�չ�[���j�=���h����itf��gژ�흅bƅ%ۤ`�� �Z���R��	B:���p�&��b���
ݷ]���g�-n�s��~��T�����Z0]t�B.��9Ĭ�Q�Qk$�S����A�#�3�zƜ1�7��tD.��b
K(}�c_��xE����#�}�.t�~�)yU &6�ૂ� -���},�'�[u�*t�6��y�_.)��f�Q+��G�◾͜��5m'�O8�%*5���,ez_�{7ǜ;��ǯ⺱|{!��D���Bo5��$�]AjsxD{�_�@�Lz~�Pm�e5���������.�I�ۨKEH�c��$V��G�:N%9��pM��JOcp%���>��s�jr�	O�~lv����X�$���	���R�3�w�To���/]Z��(gQAzPi0mT�	��F1#]��L�ֶ��>��ḻ>:�Oql��hmf�ԅ�K�\7:�20�����
���OnM������5b��ɫ�.$2�o��n�i�J��UN�Hϫ��>0؍]�g�w�h�
J�>_(�73RcB	N�;k�b97��=\��%)�jg��ɹZׇ��r�̭�$�	K5<�g��5Z�rM��CG�-222�^nV�� ��t�1��]!�H�zS��U�bkH���v��P�Ծ�\�����M�Q%W���+7Q���?�4��5��Sx���R��dF�'�HhCH��yʝ��9�M{�+��ǅe���Kg�w۵u�:�oK޼Т�a,��ybN�c���Ki>\�N7��G	���I�������w�h�ou��H��2G.�B�X�GZW��ʪ�Y0��c_]y�űdPx�F�Uդc�`â�����Ѫ[�7���e���Wþk�R�n�x�a�/$���X����V�&�[�h{�5��y�����!�:�T��*�#=l� ��#{?�w�۱��x��F��w8K���l����]}��d��x�x#�ҟg���!��P�	y$ﰃ=��v瘘\��=�[�WL���ThJ���F��$�!�s\U<;�t���M����t^[���%ݛ���_&I�nB'�E�����0�&C}�8�-+��S��Hh4�)u[�9����%�c�c*Ĩj:%��3�����k�����G�����D���m� ��`^�OfZ�$t�I���,)Ӡ������R�u&%2!�����'5�H��9k�M"Ju�Y# ���a�_&K���q��&�xI�F��}���Xm���8A!���E/dc+a1v��y}}=[�	�k��ֱ������;}���P z��6�=S#Eho�����% �S����W������<�p�e�N�,�:�*66v{ |�=���U�!)�c�)��� -N�jt�dU���ŧ������'���6�3Ϳxݛ_9�ؔ^>J�fb�xj��
�l�m)Bo��(*���z��*y�F�+Hh%��ը:\H;���}M �)��	p�3�7��ڗ�:�}�3.�G��ҮB4,f2�;Aŋ������ϴD����Y���1�\�q�>����^�"��]� 	����RL����*�,�����E0s��}�Bմ��;!��l�c�=8՗�bd3�C�?���;^�Y�\ȕ*���y�;�O��#hs作r�[ѩ�}�`^�#.��\G��T��I���/5�U��I���˿��(NCHj�$�Vc���N��dV<VL��u�fZZ�����	�?QHr��$F��7��$��.�#��1����NC�&EL��%k�D�f���%D�Y����Y�h��C��u��!����i�=��_���^�4�Q�Ҫ�[��?��#|
u�����U
`��o��
�o����ߴ)���û�u{b���Àx�
~�䃊���t�O���r��ow��(�?���&��Ƒl4a�8�:�3��(��Z�pp������e�K�P�O�ɢ���et�����R�OO!9�X�:��'�ɣ޻+XX�G�b7ONӇ���\�)�n�:��]��8��n�<��v<�����ۊ!Mԍ��=V��&@�y��.�:B�/���L�"9ʸ%����X����-l�0���s����c����kh�ƹ����$��V�T�ٳgJk^����p�TF߾�?�`�ȍz��/5����9>�w	��,�����Ս�$k?w<��G/�h��Nɘ/�J����cǨ�C���<y�=�{��^�JxfZZ!�2U�� �֖��6&HT)ڀ��->����Q,	�t]�`.8U�{Lz�4W�`�Fs�k���*]� A���������t��_c8pg���Vzo�ta�Ys:\Oz�4��5ۍ���@��˅$w!ߊ���x���A��C��\��o��L��&���m�/�tgJ��e���^�%1���'��.9sXs��=V��
u/aj�M;�E���?x���	�a"��}�~����_j�N=��{i�p)�F8�WC�e�}JKU��_��"+kz�G_8�:�Ӽ �C�0=���|�3Ւ#�����m��ep^��d�&�C���m�b(Ku�~U�y��x����4�|��:�|M��i��ق�J��V�(X�����X@�T��-��3��I�cվ}��Tj
ڹC����{~�Č�&��5>�G�Y�����a{�^����~��8�9�(0B���+�#���Kӷop�s~Ig�譢���w]d	,�H'�~���K%v�4p �w��UB�Y�HN�El�]�1���;l�?cD��q4�*ş>E��JA�
Ʈ8��o%o�:�y��	��+���50�����obl5j��T�f�}_�� ��"x���h>�ٷ�&欉�W�~���J?���X��`HEA�n�Z�0��n�+j��,F>��o5����2P��X.�=��Wm��z_t����!�+��u�1�mϞ-EL�lH�a �X��P�}M�)v��$T�"�;c!a_�Js	z7�y^������0������ˊ. zռ|��[�����n/28F���ĥdDQ�f'm^�ߜ�4���֬,���6�Ti�Q�5��,��Q�����'��)#���i���v������z���#����g�h-�>�un�.x�����U"זf
�BHv��$���;r�����@ g��* @��)�0���7�?�0RM�N��n0	���). �!�[�|� ����>'��{ׄ\.�<��]TUCC��Ȩ����bɉ?��/"{),�!��кM��� ��BYY1����;�/���(�\胧��ޑ9lBq����Sz��e�-��P{���S2EM1}�v�%��wx�g���t����ȱJ��r1gK�E��:�X�����~-*����-Mڲ�?�ӈ���-�1�Qc��'ҫ&�e�:V�
('\������Uh�SSS�"""�O���Pn��}0����pr"䪵4%Ө5�$Y������6��T��/��H��� GQ:@ Z��b��K-��`8z�x4����kاjfJQwg�DXX���-q��)��e��g�aZB��:V�O��]��\�p��n	��������ƶ����P>1�����Ȏ�~S�b�ݧq���J�g�O.9h%��?�{m-W�A7���a�r��$\lc,�$:�tH���y��=T�F��b&�+}Q@��p�6_5B��?��*<�Pf���Ӏ�@Eﾍ�o(1��,X���Ƚ��~�U�r��cP]ՙE��b��;k\�0	��R ��nX��W�^8P��K�6��FO�W0:�m�
�(��S�y�ĉ9"��s.�C�ڪ��j����1��W�2p�m���� i;ͼ;yPn�Y��$畼")T_g��r:~dD�q�U5�9�~�����kb���p���3��I��p�Kw�'�@F��:���n���0�P(ˆ)P(g��a�̂���]4l��Ch&�/��Mem%GG��`yj`O��)� \U	hX�!J>
%|��.��f��[$����������*cdd���� ��9�%��<ŉ���]M���"���U�4�u�=�&���������+����!�g�9��̝�2q�V�;ŝ�(�i&��zHT"`��7�a�
.0�W��bW���U�
Ǚ{Ec5)rh����m��S1l�C�y(7�	F��DFd|��'^�]�5�XQ���Cmi
��1�HA�ڼ���u�70�Vo?�!$ �?�.�\��ʐ��c��?�ˡr��3����-�($z���;�nb��k�Y����u`kEkρ���V!9{�{�?��-�xЊ�ohs ���4�9��Y{/�^�C�h�Hz�L�<��29�=����`��*`��X>¡�v���J�����2�`�`rK=���>j���M,KKFHG�|D����4Ӡ\π��O&��"Go�,GѸ|���N5@R�,1@KAj:%G����}$����6�GM�0)@���Mi��*����L o��7 ��|�g��!���w�V�ϳh� �k�/�h��yu�/�y1%�+��U�%����y�!Ss2���;!$m)�����/-�������������4Y�Y�Yn� ;Z6����V�8獖�9[& ����E�&!�����d\���U8a��е���ۗ�k�Ǘ_[��2�{��9�k{B̓�+�m�4�fxc��uT�y�'w�T�3������R|��'[�6Q��l�ۋۻ
��#�l���la���Q{��J8��GC����,Kͽ�����5��� ��p���B'Rz���5��	m���VKv�̂<Ov�٪�M��v=�T�P8�al
%��F��.37PĽhܰ���z��2�Q�;�+�[E�ccqXY����|kʹ?P�Y��� m�y�x)k��2�P�޻�:ş�R��`	'm"��<�����>�!��AXg,K G���b&�&�%w��>�Z�5�X%�d�ܪYgSJCD�LdP<p<=�����x���VZBv�Xv������lᓈ�Η��R����&�����{ө��[?��'���,@׬�!Q&��tZK��L�R�i˘"G��θV�0R�u�{a(z�#�,�%��Bl2rr4�s����=&-њ�cMt`M���`�(f:rđÿn�Q��wH�Z����a�3r�mY����	x� �*D�_�A�9��M��	����VO�]
j�<� ��g�(����'�\?J3M�BѨ�?KK]Ny��=�_p�-�z�)��`:�)5��ʊ�M���Ty;��58V�����n2�Y�V�����p ��-C6�)��2��3Gm��<7�Q��<��Q�d5� %��UIQ��
<����r��}�B�b�+��_��I����q���9��>As���g���I�%�r����ʂ�>PK
tHj�e�f�
,|��#F�zb�<�Maǌ�X���+��)�3�_�~�Sq7Dh!#ƴ#��_��#]PS�^sC�`�m[G��1<�ӽFg{ʾ���'�
�b���'b�^a=)�6�H�ˣ	�C��)�I}��y�n��9��cpCz:|�d��"zml�� c�X�D�$8�s��*f��k���~����
�j�����O�&t��8w!r���ڡ�u�7
/�c���h�`)�
��WԼRK�<ovC��a��G�"�S}$Ih�מ$H�h�<�?W(�cw�\��;f0�n��Q�Z)��W;Z�J��hp[w@bWq��B�EkY�C��
��X�o��7��h�cg��.<�|)pO���,�6bAduƙ�]I�����i݈>ev�>��s1$�1XB�!��'�/�;�-`��>��L�o�';�+d9�NqV尫�h�����LU��]~]����4D���$-|�L���t�|o�yV�"̾^�7z�ѓ��c�g�ѕ�N?3U�W�]���m�g���D�mbw�˃����O%��B@��m#�[$�zCR5WM���_�,(ދ�{nmv�r��$��i��?w�n �]_d��D�>u�՞������6D�����Ap�!�[�Y{3��,�|2��JR�L��=�ި��EX���,�K0h���q��!��ZE��n@;f�/V��C�b;}53t�Sz�l���)t���0������35�<߈������w��,6���O�&*Ϳ�\TS(�Q���Tr�i+CP~ŭPn0�݉1���,8�{�ը%q�}�1C��p�E�
|=�5��?�j�0?�v�mҋ�6�#��b�X�0ګT��$4�D�Я�@�������tGɇ5�I^ne��祈O��H�+����b*���ma���ZmZ�*�F[�}ۚ����蝆���7�J@+֋������O����k�/<�LT`��c�6g�﹍Y�����`�R>�cB���׃$�F�{a�3!W� �p�s��d�]����ⵐ8�Њ+6�>z�ꙧe36���L¢�0�%��>��Xu�:�=�g���єG���P�5�]]3'�C�K�Y��� ���0�;Βf�*b��E����<����.;]��Ir��n��0�&�g�D��y�eX�{� e,q���[�3u��ux͒ǌַP�7�p4bhQ�� �E�N�����l��R▋�t=��D�=�ZLV������ �es�HD
	��F����O�Ҏ��C��0�F���Tb����e* �"[��5j���2�<ѐ��y)U���?�������D�%�R�A�z�Uf��<"犿?cmQ�e	����d5F�!�h���w �!�ˏE��G|����k���`�&��ί��/`�9�u���m;.�V�m�����Iy�A(��1��y�#R�O�d~�C�%����A�I~��2���9�d��'�Ѳ�]���+o��������`��D�OL����X���ܿvRȩ�d�6� �n4��2�ų����#S~�J���εb��v r�tu.�{��O� �A4��r iF�o�X}&�:u˯$��n�^���'s�w&���S�Xz,�4�� <=��x�	�!�M��Xw�;|��^��u��2��:�A(�Ä����c
�z�T���*�8�t�Gqc�
��� �@�H�!���x�Fȶu�u��Yr.�е����P%�����:� ��Ѕ�#��N�X+��s^�}.A�%I뫄6�r�C8�[V��xi��N���CQv
>|��>���Jbu4�ֹ���ua<��-₽#p�X|!V6���ބћ��`��1�	7��kɀ�|��g�dyc$M�N[��p�����%-���g-p�z{�C��7���K��%���Bk������Rs���Qc'$�I��IXAF~�{�K�g�L�G�V��8ş5b�9�O�3װS���np�L�q�q�4�B�\@G���k��s/��$�m����}1�b������/a+c�.��hT��=V��M��v���)6�����y��%��8.W\��0�\/�k�7� g)��������I��X*��8��!)��[�o���|t)V�-���O��#�w�������*�*|z�C��Q�ķ:�̧�#����W�@�Ś3��2~i��X�}�������i׏'22\`�ۑ@��itQ/)Q(�Ug������oa@�/ U[{�yM�\��-����2��i
�e͙x��K"�g�7�7+E
����'o�v�����|��w����Ӻ&��z�	�	~k��KK�&����w�J'�}���d�¤h)L�)� ?L������&��� b���k��wP	$���t[߯SM�7p���{� JA��a���\\!gn�Kј�uǪ�{�N�!�V+��G��~h�����f��THq;�B���s4d�2�����@ȋ�¼�`ȇ���.���_���x������`�%�\�z�lm����8�F ��|����TY���4�  ��q%�F��������u��D�"�s�c�F�~R�_[-���3&Yu��0V��8h&��+%b?�^����� z̪��ֿ�7mnA��7]$r�8$*uD� �E��BCm����1g�zd8 ��ܛ=³D,�
-���qH��N��;�߲8Ce\���/�o�t�Ӂ������{g1Hh��sg�3�
܅ѓB�D֒�b������j
4��ϱ���_2�Z���
��\l|����7�ͼ������}6��)�x�/�+6���=��aS������w�WF�S��,#���6���g)M�n���X-�|��|-i�0(��y��Hј�ÄNq��ؠ�9�/s�g�rQ)��&�-(4�, Z"kjk1���*4G7����(�w٘�#��1���V�&��m�!��]�G�)
�Y �5�lG�_m59+�b�Կ�1��J��v�;F� C�@��݂��[y��%q����R~�g�A��1�"���������k-Cq�1�ے���x�jn|����<\��F�U�}�Cvv�L,�80>��k��iA��'Z��ۖ��N��ߡ�9��3^��f��֦�A��ޙ��I��&��	������"�YE$�_��?*�$��a�:	�Ǒ���T�k�:/��hM�<�����6Q^AxCμ��� O�R#�$¢�7{?g_d+�|�*x� ջ٭�5�8%Q2T�>��2�BD��H쟯h�N��]ɣn�6�/�G.���[� �a�5i�j~޴�K�tO��M�r�䍷5��X�J	��ζ������ ���)�#IE1���7�ub�#ڑ���Q]P�q[Cn�nJ��W��U�~L�)�� �8n�WoA(�U�&Y�R��N���"$Wd,`܆�޲ۑt4��(k��V80&�Hr��bޡ=��C^�'��g����nh��=�I�w-��W����N���Lz$�[i��lBq���VI�(/�a-���]a�!/51я�������鋎![�;���q6u:�uJ������jG�j|m��-#]���'S����g�*�y��H�{p r�����<��f�����%�N�áU�=D\������[k쪝l��O}#��&\
�G��Z��Q������� ���q��[��H���U���!��ۇ�����m����oÙvBD�%��{�cK;�����ɇ�bM��t�`0�$�r��?vǙI��!oNV3h!ȓoUJ�������A�A�HXVu���y].&F�I� �ڂ����
X��,�D��e�<���[ħ���0�ҟ�s��s�o��;E5\w�8f�[�~� q�ְ1Z[S����Jπ�:%�����ʃcŖ�=��y�#$���'�R��y�� 0��g ؎�\A�m�'� !MN�����0k���@��~�j̒�����.~u��,
Z�-� ����5?м���կ��?v?��3�����.q[�~)u��|�R��թ:NI@�@R�#��I�Qqܹ�4�;���"2�e�h����q���D��H��K%�]��-�r�������� 3��W��3qU���s���ℎ�?М��W�R�~r	d�-�����}c����}��Th��G�1N�~:��v��jz�D�&MC؎��Nz�)���HԸ�x<�JpV]qFN�q���)oz��h�S��G��+
_�+L�w�W����o�#$F�wr?s�O�B�/B�c"�x�;b�������D�ep��r�1D��qC?�����{U���͑o�f��3^:Q��>�u����>�F��&Y��鿁8���8C7�DC�xMD �3O���P��� 7-��mխ2_��0}C����*tt�6�����~��~>��t+c�y@+�̋V�/X�~ո�(b�*O�9������}��}�|0�@ӹ�E������c�3꠯L&L�v:����g'=�#�R�S�{�j�l	��¢������F(�]Y��� ����tG|H�����{ ��Oe�;% �=I'��"��&F�nD��'O��행��w�Ç�v���~�ӏ�e�GHy�%���eHB���+s~r�3��q��(������8��(��ض�>`�(��,�so�&m�9�}�X���.���ن޳���/�!��62�������"�\he�>��`TO����$���H�}�Xy�;���}р�M������u��'���ۼUE-7�\~O|�W�����n2���a��Ȗ��ne��=�^-j��m�����
R������\��qT���#W]m-����"���$%3���a�i-'ϻ�c�9���k���'��b�����5���|�� $������P��⁝���6Q�����c���W Q;}s�-C'��]��(!�E�o����;����o!!��*.�h�0Ƌ/��Y�*����}�g�6-8�V���6wb��5�0���ʎ�`fƤ��P�+��  ��h�ii�^o����%����7�jlw�@��~U���;(�?G^�5-{B���	6X�P�;H�l96�E�y�u�����1����4�)�0^_V&# �.b?wt,]n�[{�Q~�?�e�N`��U����A�ցL/�����ڃۿ�D��-Gk��ޅ�x�3ݔ��ֱPv��^XR�����<�b��n7�!��3 �B�*�{l��GtU��)�0�(G��n����L��o�/3E�{�'O��ovX�tK�� 1.5��dJ@������|3�Q�e��'����$�����������р'��������w�צ��?|���|Z_��~R�H%Y��p�׫/���%~Z�g�j���O\9#���"����e��0~����=�a6 ⤧G���>�p��i=]a��҄PhȆ�I]��;���N8��;�Ib��*Ե����w*>j))�����[�b���rnw�|ƭ��|f	�9���<���]�i���}�:'^�k���ӂ���t=����[�6�5:<ܓ�jer:�e�Ǐ$���6P{����ڣ�s_\�G@�V7�]{]�KIM� Ӿ�y�־�ѰO�c�)��ԙ6��з5#��+�\_F�BE����p���-�|�ҷ���[Gǟ��-i�=UlHNNN��m�F���uB�/�mq�Z�|�P��U/g���p>}��k��bo��|sWܼk��a�u�j�[0y�Jb�٨��C�ps�l� s�F�sA����G�`���߈��h�N�����9�<d�+X��̏`�㇤��{��p�I�o�f�.}��땛l6;�E] �Ì���X�������
���hXkWXWF�^ ��%�w�r��SeO����L���C"�xkN@���)�@\fR�_{|�p�%���s�>5�g��:H���2/ȓ���C��㟠��x߽̓M5�Ҥ<�g�{��e�f����m+����6j��?~]������� �c�ڬ�_��L��g�ϾFa)�'﷐/�V ��@�,����s�֜�?�i$�ٝ���P�_Y+L��o~�V���;��U��b.ݍ =6�"��h�̅�5?�?Jf��w1���TM�sp�P��3���+��i���F$#`+=���%�b�(��|��m���1dX��>S�%����&&"J�*�vb�&��ue��'�>���%�W�NDDt%F���bӒ6r\9+���$'��ÞUu�]�7��ůtyi��K�w�?(�@��"� �P+���<=��z��[TTUU�?=�S�5[��!Q}�(�!6�s�e���>)���jw,ׂ~���B��?��P�5��0�
�
���y��?:�׃����˸�{�c��@]�Q��ű@zm~=�jo��sW�Q�E�����Z���!�}���i�o*��6���ORs1ρ4�pE���ĕK=mQߏ~:`p��fz?e|��O�W�'�.�*�T�_sb���2�)�.&���>����N��C�*
H���$`Pi�����N��Y��,���7\�DXNp�d���w�gc?��a�,//�����P��O�wD�qT�G�q���4p�~Xۼ��hܺ`_P0[�Kw]�ة`9�k��@~*.����4���}O8�����͓�95�&���x�j����ն��{�o^�����'9�>��
��(~*�W'�T�f/M(����AwA�/_����ӓ��7_������k@����/-��UU��M��̓ *�k��m��%5Z�O��ڝU}�D�r��W���
� I���{�{h$=ו�\���2pj��tߴzكJ\��u ~=��ICe��a��Ύ~�l��|�'=c���S!(�9E�S��(0(�~��NQfTK���i�V㬳��6���˥Tr����-	�P�n�M�G�{(��W1��Z�n]�t��ɿ���� a�o-�K����ⱒ����L��B��"���˜7LC�K+p��������'i�ΕW��u,�e��t�����`��Vf�H:�ť�y�����u��䚟�L��4-�����4"v�;ؑ�Ġ�WMy~2���4�}�%�?�� b.����s�.��?�E����M1���������	a�k>���m1�k���!b����E�_gIMȄ�+�f7^�waX �} �g����: �hk�t����]R"( �!�%��)��tww �������{��Ο:��9{���߳�F!IM��c���F�L	W�U{�R��mn*����/�VxJ����o O��V�������G�����.+�߼����Y٨9���L����Ń'�U���	���54@��g���6����g���Oi!Cc����`�=�`��:�ۿEA�6]n13���GŎ�������P�V�@Ʀ��E��0��/�"pR܎��$�c�eY�#� T��O�e�*�(����y��#C9�uy{SE^bW�)�M=�?��F}Q=)F55Q��ھ�A��p�T�o�3Sl��������0�g�z�5�6o����(�?�d;'i��ׅ��?�!�ά��d���:��x��aWw���A��J��/I���l��=KI���+8mS$��6���� 5x�B�V�ށ�ΰE%���o�"7k���f�:X�OJJ��+0~�ջ���������V6����Gqi~:[[��̍����m� ?��{m	�<t@��f���ԴT�8��7B���K�G�"�#8	�ߍfn|�7�����P[����PvJJ��98�(B.X��B '()a�ei��u��<�o��\�<�����i3{
^>��mU�щ�E�0e��\�	�p�~����*���r�_$҄��i�������E|
{7�4�p��v��@"ѻ��%7���(���v�@�X�����VX�X(�T��� IH[����4�+2ݺn,m�繕�z��ϓ.�����^���#A[Lj��Ŭw��rr��R���.//?�e�RCBw4�;��&44���*@����������K�������8j��������,Q�aa��Et��7H�ɯǗx����|��il��_!M7�I� T�>,��'dC.�
�����N�0$+�C��Ť�P�=��3����.�=&��v zp���"�l/"��}�Ru00��P�iBgR��֞ިy���F�-���z{{髕����@ԯ�f��!z�簭���_� �+��0~l<'��_@|A���S��k�7z���:"4�E�g���)�kWkqq��Y�P�]\!�_�FHY��_6�4� PQ�nηoݛ����\pZ���	0^r6M�΋K�\�g~���@�ʩ�A�sd����P��ξ�c�355ͫ������|NW���w��@D�(뮧�+5K虙�s�$~M�}Gy	Z[��܏����B���yUU�
�៦?;56��i��p��#Ɛ�ll�OHJZ��g���jf��Į:7�s���!q�
�h�*Y�j�=#�:L(�oMk}�	�]�jk�ܟ1�.N-D-Hʦ�I+�7|�5G��7����zOv�ף��_�������'���95�֝��K�K����/<5���{�H����Vu���U;~a:PD���Kyہzy�G��������%%SN@$�@"Rq��]���W�8/��Ƀ�bҖ^[��@�Sm(3�L�<���笯v ղrA脙C4�k��V�֓ �j��˟ج�(>pns31��N/����wL�'L"����ha�uݹ�e9@0i&5�!�C����M�#����巸�8��P�Ģ�Q���G�@��jٴ�|p C$��%��Nj�C!hI.�%�=Dg_�ƒ�*���)�^�T����?`�ʝ�6N��y���mX�=�2.K^��$�|8=�!��Ƙ4zU2���]��g�,�JD-��U�r������6|4z����F����E���Y\WY���P���+��a��d9x�����7�[�z����]~����Y��ȗ	��?����#�?���3�V�_�^���8��8� �?k��*z����sw��j�s�;|�T�᱒/� HZq�x�r�}��"�C�����Ra.�*��]̒���F'&Pr���D�ϟ?�;�A�:�;���G��CY׫'�;�OR�1�-˚�.���n��F�}�#7�<�wc���g���WYY���)04>�L��o��w��5�|�
Tt�b=���<��R��}_!���Bݾf��K�78��O�H�������:kky��*�ę变M�0EΐZ�/��/��A3>D�y�����%!�t�D,��/ ]P�?6x�+ $��S���>j�k;��E腅��=��c��"�wܫ(�DH,�D���䰘�-����;����ߎ0~	��~W����3/��-�d(N@��CNE�"�����i��w֩���,a=ᧀ��4�����3�U/`o�0��Wv�de=�l��LX��C8��b�=�zB�g�^�����π6�)�ӅUc6��EU�ր � ������5%����o��-5�������gL��{J���t��d�KU\`�Ͽ�;��:o^��Z��%��\�@�.���D6���vHW0ƾ�X])M-$��&'?�V!��^7cW644�s��6�u�o�����K��1/��	�G����a�);D�b��������[#���F�h��3q����b��񄅲�+�E�c!�(�e�k��;���|�0��´4�/�_��E�������[v���h%��wv�"�����e-�;��B�<$~�ht�rk�ю4�R^��|#�Ԉ��{�c-,��E&�t�4k�>}���Jah}
DFtFR�c&iv�[���8E��Uw8[s�b���{cww~֖����Pg�xJCEHT����[��7��#��{���zǦ~)���t4hΪ(BN��}����E��|��\7E�i�gA� ̙E���AԊ~����r��5���s9���A�'����N
�c\jj(���mn��XY11��C�F��i37���7��

���5�@��9�/,*��Z$�~	���T/S��Y�:\��n>�#�`
���'�������&7.�K�`�	o��TZ�V&�����O�ʱ��s���*yjUk+)�RF��x	�pH���$k��j�3��6�I]}cK��56���Es �&L�E���ambF��P�c�q�`/�ɼn(�m�c��i�t^���j. �~�B�<<<t}z~�\�/@�-���(�.Ǻ\�)������I�%:F�ٻg�ǵ:8 ���[��rh`21�\@���J$`�����	~�F�����Mݜ���
�ǚ{��k=Nl�44�{����'rG��掵�)�a6�}ۓ��
 �)x��C���J�6w0&Y�Ȳ;�j��Ԣ�W ��7��yu���Uxu�\�?q`�������\��P�#�����2���k)��N�:���G���Ym}+Y��u�.����؝pZ��L�L�V�']d��Z6��S"�w�����S���9q���w����Dw��$�s�jF���VU���\��������J!�����(��͵��a��E�}�������"z���`��Q�;U�w�cL�f>��*��q��Z������WLg���n-�:P*��I��D���7���t�f�<�~46L>�ûn���,xz�1[��΁��e���V1�'#T�	�[[�f���q2��p?wN�y�@�3�uX�Ff��b�:\VL�1L`H����=0 �+@�QB�������i�u+�TG������A�#I##XP��|�(�п�w�uCh ���K���g�d��-��OS��2�h�䈮�a���B\ݨ�B���
�bYH�x�	�O?Y�[�gH�iG$��-�9Ł�# ��""z��B��
�M�Z#|��{��#�K0�hh��w��pj��չ���@A��p' ��˸�� } Ox�7e4�8!H[�UX�ڊx<��o��~�F�;:#iw֒P�1���R�IJ_�T7g��p
0HÒ���OԳ�	��|=�t46��J��p*�̵u����4�Hi��Æb�Pӿ�4�]����K�45;�N���D��Y։�3��|sPDݫ��F���\��5$S��G�dNRCYqD��w5D>�I�Z��F�Jf�*=ә-��wp���:������S�D��<�����nB3Du<fAYe��ܺn���f��d� �w���no�|�����|�̰�Ut\6������꣓��9:�)A�\SSc0��Ta<�k��F�����n�/
4s�pA 
�]CP>�*Dy ������Osۣʕ������YB�ma`LeUUl�`��Ga<*L;�{D��Oc�A�w�-�."�_̥�8:;��x?�ܜ��n��/X�'�"1��|��Z�)˓*~�v 8��?�xN����
Ox���T��S=��:3�WG,����u�FM�Y��-�����ù��Ox��c��pp�!m �ZwwB�z*Sf9�bl�E��qI�z��Q'	�� �3͢p?��rw(v,P�*+��`�)�G'-��Q�k{�LQ��S#�>]չ/]�7���ɖ�4�HŅ���O�L6.`�直��}�0��+v�#m�Lk^�M3-|�$�k����%��lf2Je>	�⢢.�h�=�����ނlﰃ����	�b�_�0^@
F����O�#dGv%�̛~�GO�Φ��N-��jl�� �h�y~n����������)�6U�iz�z�٣������ݫ�l��9�1>�&S��àQ�/����^
qQ��hN
�^-1MP0nD�|�bC�{ur��ۓ���	����7aΰ4�~��v-��{� ���|���9!��H�|w@+V����K�p�
r�����FҸ�B١l�&�v�x�ُ�	j��sɿn=�2�m���i��N��e�+TB?;8^�����!(�j���D��Tn�;fd��0[��@t�R���9?����b5���5�҇�-5�\�����6�9!NHL�M&@}������Ҧ�i�JX�h�;��:�c� %���Ǌ'����f�R�d+����S)�F�u�K�|z<.T��k�+�v�W�(�?���-����|'7�t�c��� �a�pY�m`^K������<�.W�ǝ�w��aI�}H֮��H"���:�e��f�f��� ,��"����6����q$��9���v�[���?|�fQ��Y����E��x_��wY��Z�BVnk:ܯjy����j0^C�8���0���pX����,4��K�?��t���e|�ma�$�ǋ��O�$�K��z	J�:���-�X9�K�ds���$b�;22R��*��X@Xs!�j�O�2@�3 �� �R���'B�w47s:.�>k�7��tM۠��6@e��bbcs�����u:�adb��{�)��#hT4]�р��TEb�Vһ=����sNS�����W�Q��C�)d�p�y3�像aL��yї���}٢���6f@>�w���IJʿKD� �؍����I�@�h<�e�C��Bw�2|>�j��o�Ia��^QQQ���!���ʛ�W���r�e�|���c���"D��D�������W#fq�v8:y%�I��XAI�,�ko����ʼ�6*�� ���V ��C�虦�}�.�?"���w��?҆������M��6��'j���S0~g$��t��m�!#��N8g�N{o_�-�qN\y�L[|���@��/q�W���n*�<rq1�kr~ޛŰW��Sƀ���MMO7i�y-Ө�5S�ׅRz�=�h ��g�1�Xfi2>��U'�~�]�eKg͘�ԑV����o�I�q���0ΈKH�o#6]LV��`5:2���X��j˗M���v0��}IDn�|��B-���Ilm\�1��?D��v�u��M�����p���������ln�aj�kd���Eag�P��2wo�S:�\��3ׯ.��?R'�y�]��C�����h"f_��d��c�j((�h4�Ӭ��
֭�P���.�	�:ˡڑ�o�NN����u��r�[/M�W�-�.e�4���'6|���e���7��.˾T!�Մ�����I�d�&�����(�Q�j׮);��V����{� �o�r�ɔaŏ�Fµ�5�V�%�O��4T�_T��E��{�lnv��p��ҿ�=oC�F���&���Nu�(�7܆*�EoXN��7t��\U[�9����O�^���>�lWp�F������B��8�2&E2{e�č�ݽQhZ ��`�Db��,�������-��P�	���d@e����Z'|��i�r����13.��̂���j_��*�0����.AD�l������nD��r�If��w�jR||�d4X�;��~��8�;;�i�[�)aVx���(&t���#=c����M��AK�a�2��1n��-:� ���6����H�y������>��V���O�|H]����C�]�r��g<}��%�7���!%�R�ǁ�Y6#A�"�a�D:S��̂�+<���/[��F��8�N(4+��п4��,3Q��c�_v�F�;T7cQ�����_�{�!��+�ʄ����j�1E����V]pP������'�<d�@�����ؓƕ�@T����;$�l2�d�7VWWO`���32$ݥ�+R��T��X$�9ꖙ�ˬ2z�1Yl�߽{�g/��*Hz�.��O��L��xDTV�n��!9V�)w���JI�Ϋ���8,F����"�ܔ�뽑D�u.l%;�~�,�DDR��-0���O��Յ.�Q�|�h!�K��I�����y���%Y̑��T���5��5�O��O(XXR��X�����VW�}\��~*�0﫶G�� ��0���<��a�ɈCS����FmQ�(�G19�^JwO�kK @���ttvĲ6���k��`Q�%}f��||�0�?�dUt4���y�Ɵ)GCh_*���u]cOR4��İ��񂙓[ϐnJ.7v�IH��(|��I}f[7n&��=!!aw����-� �/&��n�i�.�]d"ڮ[��U5e
�u#'$&q��~����p\g7uu�=CE��߫�����P%�H��א��R7!��ѱa����rnAA�R�����r��*j]֕�%����ѦL߭� ����i#�R��'�
r;��nA������+�D���s�}xdǑM4��ęE;��.mX�
��ε��\b��ҏOE�$8�%rf�)��r���5�x�?�|��I1�����fF���󃉈�̭K΀۷�}9mi�,�h��d�)���Z��ɇM�1e��N'��*iQ�-u����5nθ���L�o�sӫK��\'�����`�5-�%-�G5�Hi���K�����91�����|Y6�j��pbX/X� =�~^�n>YG�x?�g-���<���EM����+kE`꧷��/v'���q�!�-D?����X̑>��v=t���0rʢg�.�<Y�) (p��C����?!͊ML�!�����.��Lj�'A7�������5:��	'�̈-@я��������|��%'k��Y(r(4�8������g'7+�#�{������s�8��߾�17X�	�Z�i�,ۿT�J�~uᄺ+�� ^l?�����A ���0��E�S�ez�G���������L�މ�,
R�ə���+G���%Ǆ���+�����%XƧG~�&A��Ϛ�A		8����7' T�r�1�p����yejj�rQ$$�G�F�X�"n��$���#��
���Y�:e���+�f�Q~6���L�ug��`�?8D<V���M��e��!�6�"��%��!;�o^������r�+��}h�kN��B�?
%�nJ���Ad�����9�������BZ��>����	��s!�����t_6�=�*��S{�sY^^��?���ޞ�jW~E>;;��&����]�mra�����R�����Oв�T�y����66dGe�z��h�ֲv̢i��^�j�����x���?B�����<�.a�nF�El}�v��l' @��xs�j��h"�WD��5���u+��1E��Y�3�Rm�������|6��gJ��S~r��܂���~e ���?l:��.⡹�tٮ�`bcbf����JiLL@����`�]6"��rC�F���G�v;ww~;��ܪ<l��a��(��s^#���2�ʪ*��~�B�k��@�c�w��l/�[{8jx�=ҽ�q�k�v
�����䶖b�1�#����ru@0>e�õ[��*��v�p��%P����o�H��|�����lӚ�����Y;���
����;�.�w:��T&�����b��� 3.���&UkmOO.�%u�{�e
�F}�
��i������;��yN�.�˴�\�K�R3�b�Ǻ �)�ؾ��� wb����"Ep��~K)P<�W�k^&���օs/�N�3o�R��R��T�WJ
�d���>9

���:ͅ���6
Pf�T����6W���m���5�+o7� �fI����G�
�3��wt���VoV�<b����,�.�*��#��o��y�
/:����4���c	���b��~�=���UR��@5�B��5::F?6����}0�D�Rk}dT6j�w��׽��<�)��?a��*���Af�K߁x���?��T����G�90m�/,TWW}���\U���R���;B���������Ōxm8$�
�8�Hl�ʌr�P�G��K�)�����\�nD@9}]�P(��X�K،�����&5mi&���#f_�,��i|�`�]�n�$>�E9*�&�P���A�`�4
i�Wt���(�V��	@�/sh���\V�����T�@sD��ml\�3tՈ��6��yA
V8�e	��O�	�8UΣ�}f�>��<<���N��ޅ�WXFE�I=}58���<�9� ���yrbˬ�A�g�6_GM'�߇ |��Hcg].`��Fδ��-W�t�#�*�X!�N���ff�jm:����B|��G�| "�Ѵ�G�{N/�Ό��(V�z���&VVh(n] ��]�އr^��vg�#�
�(D"3[8!̬ y�����O�w�-%����`�����H � ��G6�z�:&G�����C��]��v:E��~h𣖖@Q6�d�ŕX0b�F����ffcF���
<ՙ�A�K�O�^� �g5ِ|�'"�JKKSVSqO }�����c�EMc��򁊲����eu��Zg���8!`V[�ھG�ܹN�8(�x�pF��'�H���^
��{�W˩Ț9����ssr(�j"_�JIr�
gc��F���FSۻǿP��HA��5�e�c��룦*~�|,�� ��Ќ9$44IK�"��)�k���2���%*hr�_l��0�]_��*�S����n�m敕�u��^�,.�،���?����JXJ�q�V�	њ�ߒ�RcIi��o6ӾTlrZ�_ƿ�0M1��	��WtR�z�����In[8��Pm��<��.��&2�P�����c�՘����~P@��.sc'tDQ� Q��a��gl$R�ѕ<O�����֬_�~]��d�h=�v"lbdܞ|@�G�)W�L�jy[HP�|�����ZϴT���h�P��v�Pb��˘�r�9��f���c�DL��i;Ȗ=��ֳդMhu=w��W���`&h���.U�o����pd�"ka_�2#S4��:������Q�r�#���/><o��h��v���.x��p�y��ef�܌�u�z?9FV-�-:�W����tBv~��f4�Kw��z��1{48�'�ˊ��/�,"ǐ� �3v`�g��'l0k��O>���"��"�@[y3y�^�[�Z폥r�/y����M�a�a�}e�O		�:�̆W���d�݄�M�;��Ґ�GI�.w��� �`�(��ro���,.K�vl_��;�u�_fu�E�?��%'���B�.u�n�z��;`� �G���Z������p*'䚫��V�=0��&3#�oa+agl�rM�YI1ٚo(%�Y��F���koe�Ʀ�������;��-`㡻��1�a��mл	je�b_���k��	�}���L7��Y���QS3���
4j�T���w�lTE��D�Yzݗ'�U�X� &�Xkl�zl
���Q���wD2�i��B�JJ`´fЍ�n�KA~xH���(�	���1�{�����<���&
_7�K��Ʋ�p��;��A���_���n�a�ɜ/AP����Ϙ�a$�!V��X���� 2�+�1"�!5����97�N)�Y��JQ���;m`����B�k��F6����Σ	������Hz�f��q˵��Ӯ1l��<d1H5����.Z?%2���8����u}�W�
�2>@Qv\嗦<���8=Y�g�PMx��.�s��R&j {	Oz>�g�� ��?Z�����p�<��D>������9X)�*�����`N�[�>�\GS�������Ŵ�M_���wFǆ��/��R/j}Ȓ'��Ȯ���SЗ�V������z������j������ζJ�)\�hx��F�#��А-�D�������4h �U���0��,qݏ�q��g��lT󃧡�����#zt������z���嬪}�����$���h��
���g�'������l�g�8BiQ:�E"�!�4(@��PƝv^v�ʿ�a1�$���/�Pv������tU�� T���v��)��<��+��XΞ�Y�.+s�����Q�����u3' ���t����S��:f\���
��
66�R�6&�#�V�g�]�}8�d�'2�Lv��2+|���!0ɜ�����q_C6��:����j����څ¼~��;p 	��F����ܜR���=�!��Pc���.�W��t}%�g��|�����G	.J�^��_D� j5�=>�a���RzϨ��#�=�H���ޓ�}XYy�B�i�-�{����z�:ĒQ(�dREP�rG1_�� 	��H	���j��{��"8&-),300"7;*
�g��t��邬�
;�_
�l�q}||�'>l�_{gkp
	E�`w(�!c`UˆuS-ϙ�K��Tɳ�ٲ���ѳ~d'ܼ���k�6eo؟6�s��K'$:=;J6ͼX�79�/�l��Jii���E�>_f���	{���X���#S�jy��]�=�܀�TfHL�?�p@� ����}�{���A��W��P�6+���x�������`���En�b��<dGg�	����ږ���=`M}����̲����c����`/�Y�%.!��RT�F������8i1�i��
��@.ET(�����c���p�;�$���8��uJ��Q	��)5�����8Ɣ\�8#�����!o��u>~���599a�)�������6<��AB-��m���c�R
b�nt0�ٮ���<��~&���� ͱ��cc��>�������Ϭ�[R"o�u�u�Qgg�r>�V���^�3Â0���n�<<>>~w *^��u�x���+��%�,�8�tt����D��N���كdя������+�ppa�<Ŷ�GԌtab,����MJ�Ŵ�h�ˬ�
���RU���-:=��#�Д'
J�j��G�Y�@�l�u��L�l@~���&�@�����ܿ�������K��2v�N�h*��}�J�P���c� �M3q )&-�o>>h	퐉�XG/��e`�-,-bSB���S)�o��ͬ��$�H����Βg�6���B�3X��Yvݞ�)@�Ǚ^���&#��2}�C��brfAb�D���M�ӊ
��3K�,�ɯo�4�i��x�=!ƞ2V����~��G�z�Ѷ����Y�
T��9�!�+fG~��/��n=ao4Z�����3^c�"��^�������YXZf:�����JJJ��Åc����Hd��]�Y�Sqb���a8@m�\�	?4P��ӊ6o���#0�f�|��H�I�;��z��&����F/:qY��$���-�;<_L��l��55��_ݕ�C!����p���t	��t�T&���� �xh�gw� ��U�����V{���e�]ޔE��qK���׌�|�i���''lG8��YCt4f\\��ׯ�z���Y�~x|�����O}����8Yn:��zm~U���W&�ɻ�����$�B
`s�B�aŏ�|?�3Z�o�\J��6� P�鼩O_���6M9W��V����<;?X�0�<��I�f���+��^��x1���K+q�c$l���ι�S��L�¤i�uk�b@�TV���ye8��Z@�<�.̳}��>bB\TLY�nd3KX؏������QI6�N�j�$>�)����v���B0Y��2bbIKy�nCܳ�3CCC@�Q"��е�b�u��W�~��(J��R%ZFŅ{� `�?���R��X�{���z��c���]/�jN�>�Q�)*@���	�54��ϛ�i_��&+D�V�)���GC�y#7>7�{��U�ƕ!8�;���������봇S�{(�#R��۝����������dw���^�|Lrv0�)�~S'���EN�9ϲ�?��m�D�NV��<�ˬ33nM��=��=�T�c�%��@U�
���]�s1�Ţ�C�*B����M��� ���g��{j:���!�F�F1qi0,389�HNR���h��j~̙��KF���Gm-����+���fX�f��q�h�^p������z|����=_�Xw3��a�Y�r������ש-5,ϩB�?<�F����B�߶P4*�6dsm��(Sʰ���j�M����&��W�����ONO�3�!��0�|d����G���63�Lܒ�'�VPR��ad/���R���b>
���}���E��|�/vvv�L��A".�HT���@��Q�d���=��-AFA��$�^C��lۢT��W�j�>�ݯ��<�+��|w��=]�n��w����Uw���{� �WAYc��������^��ا���L�C7*[D_`~�\��4
��]��/���]s@l�d͐�J��9Β$�����h�e�r��ae�6����)^���%��Y��� ���	�%UN���e�T7�Tj5	+��np���)J ��t������ϝ���2Q��e��+'�}���?��*�};�k��>@�������L,��xB��?NNN���P�\�Į�������[2��Έ�ŧ��J��M�����i�(�0�Z�؝�'#�pGx���MeBR��im�F���_�.��=�w�YΔ�%.�mT�
;�j��3��Eb���Ok�o�&�gx��H]⏊���_�i�(%��M��Aڜ�]�++���/�J��U���l����o����Y\]�������%�R518(')}FA���&H���Cu�����]���No��U�j��f��+���Ci*ՉfH��������Yy�3�z�Z`>Q���.aW�!2P�����UD���&Bd8�	����G=����O&3�N�9u�Ba�os�񡔈E�؄�جtzi�rCڻ9���8H�&��2����?݇r'�C�=�Lꥫ�F�P5g���mh~�Q��F�_��*��.22�a���t�{��-qf\�	�@q
C#�z
%�U08�E���hbb���
���l���Ҿ��K[f���g��!��ʛ�	N��sHh(�����Dc�ؖ�疖 ���p���200�q��K*�;wºh{ʺ9x�ًf��R���2$:����t�N�s��nꂍ�d�+�=��Z^^�Ж�7�L�v�����ڡm�_K��'L�@�WH][���7@
i� �����Q75�~�"􏼼��w�Q�RҊ���?Ȓ������IG��,����9�m�	'�J�v~aa��p �r>x (�Y��װ���?Ҿ�l���ʌ���Χ��bc_����YZV8jr6�n;���?�]����b���b>=|_Ⱥ�$!�q$�䘫a��ZRFbH�z���v
$d�GXb���F����҆Dm|AT���=��L[	rW�����e/�e�PWǫ�$0�V/��K;�v	]�܍ �������YՔ 8��Yݢ�G8���Ofm���?E�R0��Yg+��Y��X[3 �!��B�>��0N�)ۮ���t�"�n��ϜΟ?��K��[�>e!�բ��� K�=��(��R2²���GM���-9~H�}ɹ]tX������+����-d-e?���=���a�D���}xd��y�䙁W��#44R*�(�u-2i
� W|=�d��k}N�p�@�q���P�"Pec��+�k(���� �MG<��Ы&Q��j d�Jlm�]����O���$�z��5�J�����}|�s�r��#�+��,m�Pʈ	���}#k*I��v:��B%��j�Z��VO]cp����R�;�x�S�m���_���{*66L`Xݿ9�,��iiʅ���Z�\��éIY�G�T�1���#�{Yse?�!����p�p�����kt4U�U@�ঊԢB3;�^��Ը��(a?Uv�/Y�0m�`U�1����KP����?����X�m�%~NʎCSK+�5ȍζ`����޻
�
�b� ���+�E��k��]<��h1�V�����Ё�A�R������`��/%�2�.�#fhHi�x7lV���GQ�%���!'�?���r��j�z+嘵p��2|k��Y�I��bX>�x]/�����  "���5���`�	T3��2�?j��`%�l�
�+�7]~P�_��j�-�������ޮg�N�H�S�6�W��!���m�~{���w)8�[Yoj�>�ӵ�BN�a�CP�������BϘи;`Q���9X/>�Š:�������Z��D�ժ9+ދ	W�X�51666��R���.Ʋ�Hg�g��ӽ=fM��#a�P��5�(�v7��j����T����aJ�ӽ}�z��w���bӣ�Hpz��xy�9�}J��!��0����@��Ϥ>���[�> 	�g#ư�r���� q
kE >�k�RUtz}�ǹ��hB���_~�rs���l��095EE%��2�>��
����Ҳ��XOꃙO��/j�������˩��߿�i��渃W�NrsЧ����\Z=缳R$}��f=����5��MgJTo�b�(����7�	��������9��5�����5vb�j�y��D�����Я�X��!�v;*���o�YY`�C��:�D�$��$&J7x޾۲���i�3ve	��較�a/P��2)��ř�aZ�6�3�����xɧ�p��՘Eu�������_�8;;���^r?����R.U���J�������Ҫ;�6��. �syg��|,�5Ǔ���]\���0���"0DL�W���O�����ՍQ���ݝ��ό�H�e:MAp�����I��=ڣ���ц{s~yO`؊�x�������h���{�(���k�@�$�����fp����f@Tƻ҃Ȇ4����cD��j��{]�D���I��f��k� v�p� �]�!��A����h��5_v捇T�}����D/�7\������3�u+�xl$�M���Ҏ?�}�VYE-�F>�%d��9A�t����#?	(����Ȉ(��-)Q�eX�#������At�N�&���%��� y���aœWY��3OH�8��(����qg䨟_��s5h� �T_�m��|�5t�1O�*��F�\-Z����������))���Kl�ث��EL��S%�j�-�g��2=�yy�3�}>(��р+T� ��-w��4����9��/6+V�����r�U����I?���˘�ט���\�ܿK����_��'1�y�u� �2 0�	I��/�W]�~'2�(�BVn�l7�����F$�;$*�Zޚ�)ޫW�|IF�a1�e!m�ٖ������!�,9�Pc�]`B�~6�k��4�ZҮ�����1�(���*���2� �Ir�یw�ƾ���I��CZ����q|�0�b!th��PX�p�
�ňA<Gp���?�?zeywO�k`k;�t�L�f	.Aj���ӧO8@Y%�Ѧ,(*/���R��d���"�NcȰ���`�����Zc2��rS8�n�����rc�E�j�aUx�����n�D,�`�@P��R���
%6�+��Em�w��|�����,�(;ؽ�"=��Y�&?�1����Sm�x
�;8�/z�����D�P��-���L��ժ����HQ^AU^�L��f�x�2������Ƈ��9|L�h� �Bz�&���]�b����ra�1��μF������q����$��  ���N�i�ۥ�軄vvyo���%m!�pxHc�ڌ�n�
��5J[�ǧ��wB�V+�}� I�1-��XFqj�5����/�mm���e��A��u���'q��yCz�����!�`��ZZ ���O&[�=ȗ*X���0�!ȧ��IfZ�{I�7yK��h�3��(`��x��<��[9��p��J��,������H?�())�x��T�;&E�'Ue�ɫ+N��iѮC ,fy��� <��R��#��{�}X����Z�gx�G�u�e�o϶��I1���t跋� VK�G��`�j�'o��[KOز��H�c6Č�� T� .!�Yr&r �-߼�X�|0o4g��D�������QOj6��e�z���<��&C<��Ci��`���!]��8�G�������*z���Vz 2 a��o�����)��:��I`�1�rTUŖ{CSl������1Z,%���|��i�/�pn���� {��2�ˮ�N��}6�K%@R7i�_�����U�]C�"%Y<q�~h�uu�����6��Fn�5�&��tpXmmϽ�b�+~�C���8����� Z�3n����K�.T�l
�l�&p�*ؿi�뀺����t\�8gT��
;4�j�I~�wLP-$2�����MޕZ����:,�i��tw#!�R���  K� �]� ��-� ��"! ]���}����������g眙��{��.l5pC���\�T�B��]�I����6�m�t�LK�1u����-so����>�X�����=iH@ ��5Œ����1:&́~� C�T���0i).3P�2lăp��iA�sEx ҁ^;v|��Ȱ���p'G,�~�[�NS��������yDooC�������F^Ak�tG��$�$AhD����\����m��)<0�A�iFΗ��7�x�>�.�]���W�%%'G��HL�`��8������D�*�8��J;�P�t����&A�s-���(�1�Vt,�R�Ғ'Xi� ��_�A��˃���e$�9��<r1IH�z��Y��ܨ.M�Sz_z|X�mU6���
�&������z��Y�puI�3S"�a���O!;.`���W�h�����!033���:V��K�������=)*, �����J�}�taƂ;�WV"6ʲ�f&���V�#�?u��^�#���P7+��=�C�p9u�3g�ߒWZp���C�ݞ�����'�=�V �ɑ��S҇@Q11�����@n�$	Xx;��6���1vs}��@Qi���`���䠟Q�-���P���
�	���j��"�����r�Og�|!,:��+1IR-r�A�(  ��4R.�W+�d.g@�)o.W���r6Q:6 \��HHH��٠���͝�v��&\DX�@;�����ȡ�փQ,���u4�|888��-��q!?�c���uNA�����*X{)��@�v��n�X%8p��i�k�*DC!�M��ʠ&U#_q���8:��Y��Zw5�����"�eV��<�xO��=~w���c�(���ӯ|2�uAX%;114rU�{��۴a�ݒY����>���gl\�;_��Jvy}d� \��W�Ø������`��
�7x�����,_{��@����t�bL0�l������19���:�{��uf	tѨ<���|�'�9�Ӿg��[b�$)^!` ��HeeQ�In�㑒�s���O㻇|$�mmߛ���k#`�o�"������/��`��f�t�
���O���:����	��ġ<BBa��ּ��#�#�<�e�8xQ��ֳi����q�ܼ)�3����� �)&߮���hK4'�ۤ$m�}%징-�R�p���Ȁy���·T�[s���dQ�m�O	�G�	��x��D݋w/�Bl�<Ľԋ\�@	�*f�����ꚭ�`Uq�#��V�L��S�w��Y�`��P�u�G�>iS��9��M��zc�#[ �je�W�Z�6���*����C��{;fοo�lǦ�J�1n�����q�����"���s!v�����3+���	����ef޾�i�.@)0��L6��.e.�k��
s�2B'F+_6��u^Y����Kp�I�@t*-���Z�玥�ѽ����r��� ,��e�<5� �M�e�x~q�c��C����Ӂ,���]w�/K�u| �"!���u���w�x12���`�R��U���5C \��j�h�Bs�t	T;��Z1�v�7E�Yq�L=泷o�>�gI�ܜ��zG�ɘ]��B���m���Բr��O��!( >�P:=�ӟ8J	�_���`!��,uY,�x`�0��D��X��i�B���+������r�2�3kۏ�P�
ݬ
Dd�5j����"]9[�22~�bS�Ҫ*�i�1��y&�g�Qd�6�%�Q1Df$�������Tb�E�Z6�z ��4leG��B"G~矎P2��,�GNf���3��j��l�)H�L�EE�Nw���O� ���z찾^ɳ5�$:zzDҨ��7���щ+��I��l��8M��z��žW�������ES"�_��u�ML�n ����s wk�7�5��f���
"__�%;�x������1h~U73>iM���>ln,���8��W�~M�Q�n;�	á�N �t�n巾˅�Ͻ�"��݁f�v��ϯ�����&��8�kyF�13UBrrhB{i�M!��N��au� �bʢy�ZR�S���������H�����ӕ������8$-��Im�İ������F��$��w>7*�+{��靊�7S��<�?4R>).����VB4[�P����m#U����ߛ���hh hj�e��#��dx�P�jD� ��,&O�р:����;E�-}�����s\�J�G�*>�5hu;!;��aD��C-{�Z�##QԾ�%f�	���/JH��%B��z�qq���4(���B$�϶�E�X�g$�lˎ�t�@gNdĠ��$m��jn�)�:W�e`͂�0[�z����q��r*js��u�^^D��o��m}SÏ�q�Pb�z��zK;;rT>�1������?�|7�:'8���D��87�؟������-��;W�.�ʯyo����A�s#����V{�GԋE3:�XR�'�lb7Ic���ٱDu�&����E�3��UT �$)9�@$������T�	g��L�`܄A�[Xn�+���p��.�mG)++3�<>i]� �<6�7L�h��B��������7�ӑGӋ�����u>O
4O�ՠ���$V�$�R�~�K������(�c�.����*�O����ܵ �C�p׭�� �/g��|4�s����e�i6W�V�)G�m{R���V304Ӵ~����~����>��v��SAO�?,�HU -U��E/Iu��i�x$�JA������j>>���g
x���_|��5
F�FA�l�-�7C���ݞ�T������U�6�P�
�lǠ&�8߇���R>|�?��6YS�%�m"�j�hGBڐq�E����V�OGG���>���͐�j����rMM|3s�W���f�4����Gn+��sm�e2��m|���ͽ�I��͛��B��i.c����N��~ ��@�JQb��ҡ��U���3�+CC@9sw:gt�Y9�5>1�>M��u��)��������I��`�
�L��������9
D܇���j�O��ж�/��z�!�3�w�H3� ���\��.���j(��M?FbzT^�����o������� ��4�,tqqћ����j�Z(hV�u��p/^m��>Ԙ������WP��[Ӑ%>8:��ʘ��;Q�>wզ[��+H+?��P�����ZI� 2"Ӏ_�Zhz��[�%�۬��ϭO�=��n��!�[ C[��q:�:飖@��fHK��V]}�]T���iE���Uk&ĥ��-#��.u|d`��/_l�3�I�`v{Z��쏀�D�5���:�ov�ohh@ ]�����p[dT�މ�����.��>��5�;�d)�|�ޅ�����{���js�f"�=:#�b(ݎ�ףa�t�����iiRVr!��[b(�H&ʅ���9��8����*.�R�[���q������Y[�ks���t{s#Үx&�Q���Y�X?rpP>�� 7'��
�5 �W<�Ү���4�$������^]]9��h�]��U�z�(y�>�yO����Zv��ڼ)�{��@�E�b:��t�u�?�}�P�L��/�N?����և�ys���1U[�_B6�[�������l���a`l�?���2p,|mK��D���+��:�ŗG��������bD��.�^�����J�QQ>��F�ӕ�4�h��<>���bMEY���ʿ��t��^ThONO�X��&ྺ��[����d��o���U%�1�7��~KZdɋ/�����%�B��߳�|��k�9e�ФSk�V\��@%�o:D��a��(�伟
KG�c���C�,g>6�\�#7����B]n`��V�nOhϿҼf"U��	�s�&S�b^G��� �|~%e��J�"�󴩰��w����9C�d<��3I��K'�5q�/�9�<��� ~���}1w��I:��i�����VXD�&y�]�c �Q�c~�Kp���&vv�F����Lб$Ʀ/����б�d��a�{����䳾� 8��R�F��E�n� fi��͗��e���a�o��++���R����Uؓ�zo$LT�5�؝Wu�Q�y�U��=��!$($��Ё]%K<
���^A��0���X��377gJ����9
gb�;�B%�JP0��Jց|YHCǃWPPл������a�<��5�Z/�RRBW|v6l��h����L�y i5d-�G=M��9#d�2@;/��L ��ʺ��_��skJ���3�eI)s8I��kg��4z���6��ĸ�kK��A;_eS������O{�f�-\Z�e�j�°^ZkR��Kٯ$jdI1b�ć��}.�v��{���k���%xW��~U�M�ѱ�����Vc��U���<��'�:F�J���K��F@
8����S��e$ ݪ<"|��s�H2�~	n�w��1%��c��:3��=����V�ڗ��?��Z�a�'���e�?S�Vx�X��ojJ���:v-lt*"�K�Ƕ�!�Q��Ї�St�_Y�~�i5e�pZ�-^n�]�O�KKK�Y�9��7�6~���S���Pg���p>V���I�i=��4e���r�����` �uv�d��<���D�f�.kqe�SOO��*��g [z�Q!���hM�d��W�'l��'������h�t�-D�LL��nE�/�vb�.P��D߻'W�����'�UO z�ܜ<��HA��v�-�>�e&��u�-,�LWԝA�%o���`�w~�--N���Z��V&v�R��|�	ʿ'��9u\n{�v^H呺dr������eZ��s^z,�
={�u���rz���1����;>l�d p��?�8HJJ~kv������W�	j� ���
ǢS����ݷ���}H��95hܺY3.��Qґ1mB�B`W���=6�x��eA����.#)��ݨ=З���OCCä�D'F��7�C�@�S4p�����/���_|ϐ%i�FR1#���M�v�E�\d���wQ�8���wF�3��%=l����k:>����oj"����@��@��%�{9>/���c����X�|U}��-`����WW�o(�����㔝/'_���bL���:ֈGm���G+��9��M܂�0pu��)����r����|�DF�"�믦��>��3O�2pت��|����"vKh�f���]���[������m(����F[F�u*���6>K��9'15`̺��(��d��;��V, d��w4r��	D��y/̃�
4}
tYE1�Y��J.5�]�����5�|����/0�噦���6oЇrP'�Co=�ku�N�K�&�k�ZG+����)�a�D���/���G��r���Ͽ]������zP���Xh�힞&��h������ԣ���_�)l���6��aK3�8��kH�Ǻ��?U�o"�����,hz7��>�	+!��z�憥�|���>22�S~ENdlp0�����?�T�?��և��F�!F���������v偓����k|��l�����.;�f'wB�3HBB�^AO�W>��c3d�X)�������@Q��N�~*����+Y^���`ұ�3d\q֏.��z�ml�<�ng�76�q�g�����6�ڀ��}�(,�?C�;s"��f	y˒�#,�w���E�9P�ց��P����������9Fb�sfV�)?��e����}%�*�Zj���	Nnnn��i��'T�dI� [P,�}����h:��]�<��:���Eڛw?��t6�<E)-\��ۧa���q��$�T��2�|2���/��mhpDF��ü����oّ건)��se#j�}	�G�+��=*mM���' [�W��踧Ǹ���M�� ,0�z�d���)Qqy	4�)�_�ŋŻF����*d�����A�솿��7��\^�X��_��9V���z�H�v�"�� �Og��2��)(d��1�pp�M�((0�t�+�!QP`���RcF?sXTV��JN��-��?�H5������ �l�A$?�����^GT-Q��+���"�ˇɄ�T]�Ѵ=��Kn�� C�m;���Ѩ�? � f>@��iD�[f]�zj� �#���u�s��h	wK�7�9�bS	b	ٞ�$s�%}�B]ZF���+�#;�u�����)N����C�&E`
��܏����RC�?�7�b����7��U�J�L!�/,���઩)������y�D[��z�����y�.��>0���u��AC�K�Q��X�_3���P3
���.�(�E��Z�#�|4G��B�����d��@FD|C�|�es4]��|�>������b��YғZS�Va�����`���X�G�i55\�ëG�W�@诨`öz	�k�e@��q�=���cWXa2!;�v����E���1R��+Im��7���k���� D�2	��~}�'Iyt?�̔4�w�>�HA��f����t��W ��y	���I�8���a͠�m�E�ܵ�i\�f{~�����h��#i���G�F����?�9d�H!���vRgy2q�3_�廽���usmu>��}�RZVj�/;�}����9�ڳ3�4��}g°��h�F����hC�hYʟP12*n��
���N6,;i�LO4j��%z�R$=+^/�����Z���l�ůƥ�Xx�ɍ�yCz�ZQ[�6�o;���LE���;삣`%��z��G!=�p�t||��>�.�D����vp�n`��B��	��y"c��{�ϖ2=O.S'5�?�ۜ9s���w�\P���Ll�;�,N�����\�?v�9C����̔�KM2(ٽc�Ar��ڰ��_�ϯ4,>��� ���2�wr�|�q�F�f-m�-ETttn~3�rT�"  �^T4lwn~�B�5�Ji$IG�^�щ�v��_z������ȎI܉ַ�WeU�hr��}CU�mP}T�Ii�����zS�00ԫV�y"��i��u����1����=�q;=���ցtba��'E)�wN�.�-���<{n����a7h���3���b1��q5�t�#.x_�Ue)��5�2T��(�x��sr�@�#��ĳ��O��=ۭLL@0�?+��d�#�z}]cf�Q_ϻ+R�h�@�4��Y�h�p�]e59�3��_3�}vI�PHI�Ct�޹���dc��1�t�)�)��T6�;W;�U+�?�Ɂ�A�>��3�HHgc�T_/O���t�P���Tat'G
��J�먩�c���h"���(�ᨱ�N�{�����=3k��A(��_�#f1�4���=o�z��a=2��=��rf��d��J0u_VN��X�mqq1bK�{�^���U���/;��ߜ����9�=���h�R(->���f�~ �LL-�*�����!]L�c����=s�� ��B���5Y�m��ݹαxǴ�Ð��̏�e�x_��P/x��zy�l2�F) �u��V�?k��.�����)���;�o+��iOC���h?�q\jX�~���1����qp�ц��a�������O�1���}p�����`���Y�'V�������/6���eQ����z�e����1��j�>�6l�0���=���!X�̵�>�2S�3wq�eT��MG���vX)T��z~�W �*1�S��To2��ml��]���cx�.;������hn�(�W]/p�Cѷ�+r�J��:��5߸[]�i}�욒0O)�:t��v����(��ag�f/��5W�k̝�3s��'�	X��|�<)���B��b.�%���r�R㜰0��0���6^T���Y����f�3��5{�O����l!=���g"�ʴâ�l����?M��芟춍�mGek�+!�@�s�PL�v��,����a��^a�Ye_oo `�����ZJJ�5b^W��U�!�u�:�=gӕaѴ�S6�ZZ��s��ceG���H�pv���/3*����q��N�M[OЭ��jxH�B%}4X�=.nM��w�Էp�(m����T%k�� �m�ש�(��A<Y��;�RJZ� �hjjRss�� &e�ա��酧��{����g/�9�q�$&'���}�Ȭ�j�n��>?��$��?1��/�
/kh�WQ���1
G�Ni��W������V�`2:[b�-9&�"Vb�AWC��Zܰ�0��Y/��y8-�lHHH2r8��9mmd6�@�]�=>��z#�|�2�"�$1��}��cICuux3ȵ�33��ñ���5�=R���9�9�<~Շ�	z�uM2tĻp!��6�6A�e}��/12�#éI�ME�`�H�43�`����w�bpu�nƎ���Z�z�M�S-�Wx٨����4*Ex��A����J�W;�;86,�<�[��o4�P�B;��No$��5����YD4��� J)��L-���׋^��rڋ ׊�ܶ�xJ�wF-]�)�,.��䔖Q�cnNV�3?қ��_�M�`.���2h����1���X��9���p4+�iT��R�f>f�l�x��Ș����U's��9?����]ZU����6�fu�Y�*X���� ���b��=�=6��/,DH��y	��/>q`����٭��gߘ�gpc���� �������Uб"r��%�1���0 ���#Q���������"�dG@C# q���_��
��&պd.�o@=$�����w�����S(`���3u�t7��o��9�b��.j��x��EG�����qqsÞ����)��$�W����r�
�RG'�)L
�?��#�����kpƮ]���\||�]o�Ǳ���� C%nm���B5��_���}�gR��?BXw[`�-AL�-�<�

�/ƇZ����4�����0 ԹI�f�yؒK]KHL�'��Cz�Yt�p���Sn>��%^�Y#g�0k��� ��QYK�A3�͇�.����Ѵh<X��lh� �����G݈}w#�M�j�&'y�Z4�c�2��(����l
5 Ҙ�NF��ϟ��)��fa�%!!����6?�k�2�3��gg������^�0U�z/�C�g'�=ݗr��TPa���ϑ� �������ϒ^�w��os�ܥ��I����/(�Mi8"gHx(�7�<
Y�y2!=�B���VY5�uq?L�KKc���p$jYG��K>��L�<���Q������ ����sU���1��6��>��_�{zz�l�j�����ojZi���ܵO0��n�F���v�^w�r�k˕V�^01���:W��[��N�[*⨧%cf[��D_�ʯ\L>	��OTdj��~�p��
��&$�F������r��@)�|}��z��By�_���d���]� �mK.!>�$��M--ӹF{4
9����λ�Wv��r�x��ͬ��K^e���udwP]�og���: |W�@"�j�x���%�Zs���_d p�=wE@\<������UX�� 9�k�XX�///g;HۜŅO��|%&7o���pȹA�}��a�#��B�J�2��P�FX�����xZ���*)�| ����Π������q����)[]�'9�}A��s?��GYHyxL�������@~8ec�n	�cn����EI*)En
�,7�jfb��5��R`0�g
��6w�-����5��,�]���q������P��Y�8�����V���":&&yW���ui>R���G=EG�� = �}��e�ʁ�����%��o�D��ߵ>*���ŕ٠�M�i�K�	����7�h֔��c�`'sL�Koف؎�bV���?F,�U�8,��	2ZAg��
�˂��9<�b��E���KB�C���\~�}�ד�A�����v�@�.�$�-�(�6�A�\�����|���]h(
�+�n�g�S�\`�s��z9�g~g(b�N���ָ��
@ƒ�m���I�q��8]e�tE�==��?n%feQ-���4iS�f4��n�{��+*B�E���>�Ӵt3s���яFL�\����U�T
���h~y?�Aܟ�.d��\�ejЧ��;)E=���@���o~DJ6�����~��'ަ(?�As�+�r��k0�������Cσ%�w�����4��p5�<���Z��=�����ꮛ�	II�kb���2>��3*|�)���I��� ��p��[�����?\_|���6��_%x)Ȫ�TJ���?PK   ��!Y~��k�6 4 /   images/663b53f5-e86a-4272-a51e-f5b809259b46.png�yTS��6D��U0�*�n�4JTP��� ݠТ�
A	CP�y��j��mQ�L�4�@ ����@E� 4$"B� ���пw}�ߟ�ֻ����^<U�k�g?��u��/������[��O$'nE%���W��o��� ~,=󟟏|F�W>𿿦�t����G�ɩ#��/ׇڸ����;�7:D;s���(��_��b�	�3��G"2G))�)	�-�H��[_Ɨ�e|_Ɨ�e|_Ɨ�e|_Ɨ��H�<�/p�������/���2��/���2��/���2��/����bl�9�Ϸ �?��7��S�9gζ���Mт��řv�����'�6~�t�y뽇N�ugKZ����������E?�G�'���O�0^}b�r/��̪�=9�����g4K�?E�d06:�b՚*������2��/���2��/����6�!7������CSoo�Q�ا>�:��3�"�ܾ�yT�_Ƴ��1\�yk8�v~�V�����g���d)N�.�х�I�3L&�}z��U�B����I����Os���:�O�@�bt����j�A��,��YZ�Qr�p��`���5��^Jt�l��3g��g0�������ҀŌ��~~�hcG����a{	|�K� ZZ��,��%�o17�����2`�`�~r�p�*3�������(�w�2"Ɂ���@�hy��ON�����x�*���/lU��b���].�?W�-�H$+
?����%{�1��x�EF��*�2��K����AZ�� ߸�����4@��_0+��r�� ���g��O���D����N�ʲ��\�C����6t2*�vnȺ_`�",������Y�;����Ui-j����L72{=��H�5����CB�:�F;���k*�3{vaa�q5���[X@���n�2T7Nah���-$NTײ�ڐ�����	]�8�scO�*�XwF��)(7�x��xλ��r�	�F��(��s�����1�QP�Ƞ~���4*��M<7p�'��Q�A�����"�t�A���t���#ڇ����l4}����c�v����b�|bTx��DǑ=���M&BI�$������.�k��>Ը|�B���C��VQ	Z���L:gO�]9����C'�K�Q�x��ߵ?^˫�S��ai6Ǘj��:ٗ�`4|x��Ǐ�_�~��*Z�&c'ո����L.����\쓷RE���a���<�g�$ݽ��̈�r�3'�0J�����:=�3#��a+�^�V��65�Lm4�����Ne��w�7S3�9�70^0�͈����Y��K(��34=A�)WB�ێ����%`	c�y��j^�1��!���Rc�	1�'��p�<�M[`L ~��*3���gϞ�~zi�����'��&�\f�1#��4�j����]IG���C�������<^ֹn̎�1;�CvOm4��bD������:����xY9_"�ğ{t{[!��9�	�9�^��I�s7��'�b<IT��V��1 �y��lb�H
�O��ƞٍ�݄(�S@���<H����$��Q���������*�� jA2�Zf9X_c��i/Gӵ�����={6(���������	�#���Tr{��@y�?~�O>����~c/o����J\��ê�Ȼ��sQ�T�&��`j�11�<�C��,��
NW�M��}�*��<�~UhNHLө�����N/M|z�u�~zԳ@��}�<9����>b�F4����eЈ��Ӎ��֧6��0��D�z���j�4 'O��
TL&^rd��z�s��?�iV�c���4˼��i�����^�� w,>�qt=��c�H�����¦�F�������To�z�b�!~ԅN�m��m���NAn�>13��wSEB���H�zE�^`M��F����W +6fo��I(ƽñ�5�!L�~q�"�qP�ܞ̜��g�A��m��+*��-��f����-t�3�B�u�9��`����5����h������;�s�F�,���Ը���3��G_LY�f6 |G�����#��n#�[K�Dp6�x��}�o�=�{��x=��b��r8�r'6�̉������.�\��]��wz�;Ñ��fG��l������mG��C6�$�'��]���drd��ߘ�F�/�M&&�3�/|N�^���7xօP=\�ۭ�
2�hƩ�VS%�w��>t7�ޓ�lu�;���+Qm�YP�����D7y�s^N+/����{G_�\��F����x�|vv6���	e������?lf�J�����ߧ3���_��- �:�~>�fE�Bp�:�|G7ӬEIĕ�@s�&9��ͼ
Q33҃t�b�\v��=��7f��Q�n�C~��^��ӯ`K����4d|c�3�p���2�����|+3���MhN�+v�՝==D恾_��.6��3p	��w�t��(�EE �B V`��Z������-_8��w4ՓL�VJ��gLSɱ�eq�.E/�v.Ϊӛ`j��������]���	A�u�ݾW�jS}RwCu]7/���E##v##��-���x�'w��}M�������r�E|+��Ң�����A�@Ɋ\�Ew�{��]G�p���̙d�a�t��,m�_Ѵ�����������_w�F/�PW0���Idjw/�/��0_:���}��9)�s�
?t���qt:�SS`U�jh�����]��?�ÀBj:�'��/0�����q�<쌮7'Zs��u/�jF�>�U�,�T�;�O��E�t"�qF���o0s(G�FzQ���jpئ�sY�c��'�A��)fNkK*�}���ݶ���ej�W���p:0�
n�I��,��،`T�QR��W^^�>5�9���=��*��U�쩔��mD� �y��z�E)�lA��i��v07��r�m+������X4�;� ��?�ɖZ��הhiSS��%�%X�C,���:\QΏ�$,���.������?�.*�*~XW'�KVw�1���s��C�J���|ud3���F9��{��̈�EZ��B9�If����O���0�O��K�B�W��6Y/�>��X�[���]X�|a�{����x{ژ��~-��b����@W-��z6��
a׾b7A��=m ��g�26����6�K	�bq�H�	D�	��6�dE��=���f��0��܍�!뺺�ɽ�F�������_��Ved�%��<��陙>��"
0v�:b�(Z� �F�����cG 2T�ysA��0-�Z֙�O�U�Db��L]��,�Ί�֫�����J���+B��&��>�e�Y�X����<��s��y�,����r3T����H��ŵ-�ڋ����y���ڨ�eO�Cql��G�a�/cz�f�l������~�����ݻwS�b��,d��n���0Am�:�R 1���L�".?Ƣ����w�j��橐�]������+d��b/�S��E�JlA&R=F]8M*�.�Y?=�}~W��ѣ3��l�t��[ I:_��,���S�NBG��S���Y���"��o�E/ߙ�eJ&��#�1�% �0�t%C��y�n� �G�Z�="��K���LФ����?���;�`:H���pc(J��)�`��bL��ئ�ZW�c(G��`%驲v��j.ڵ��������B��@>���k���\�7�,�h��յA��{\56P�O@Z�'��!�Ȭ�@r{��H
ڷ�K)�!�L�� �;d�f�i#u�M��y?���A-���,���W!��x ��Y��ߤ"Ux[�'(̌�y��Wi�L�DD�u"##�o�R����N���"��&�����?�ݎF�"��p�U�6�E���"%���u�s{}�C��oѳ�A�����踙�7�C8�VO&B=Ȗk�Ҭ��o2�3Jk)�m�k!(�̒Tn��h=K��L�6a�X��Dn��)参��9}���Hr�2�b#"h#���
���Y�bՁ�G�g�uT"���+��Z��U� ?7rX4y������<�vP����u��$�F�ҙ�.�71��
JH����}9 #6�'�@'�tHc�B��Ħ�>:@��xB@��fjY�?A؁��M�ΉN�aY"6W����1N�����=t�����{�Cn4d'Q^���Rۋ�b����Ug�ꔵ����������[�V~���s�1���Z���⩑�S~���'ZZ��+�TFo��O;�pZK�J�$q��Q����U�j�0Ys�I���D�\*sfpp|Z�p�Q��%5Һ�3n���?�Ŝ��{�����n�1;�T���0,Tl�Į���.��oMd��%Q`���ۉ
��빯Gd�FL���=�O��+D������C�y�`��>���D���M65�&ƠV�3��_&g�2����E����A~q�_��j}ʹ�vR(�ܿFP~f�U7w��G��%ݩ�w���J�2]�z��`���-TN�-^=�葆�R��Ϯ�K�7:5Ǧ�58v2/f������\w[f���vl ժ�?+ ��M��U_a��@�y��TF]P�J}��</�o�d�(b�'��Ю�yi��k����t�RI���<x@�bo�w4R�i�z@���t/L,�l��Ż�E��9��#�P$̔�r�����n��D;}6z�:�aC]��r����^�� �ÿ3��:GA���������0p4�A����/>�=OKcv��'Y��>=G��:'XO�}܅y���k02^�-�>�T:�z����~4RN��蚾=�=�x���\��s�����4����ⲟ�u�\kc��e�X��&L�a�_ �[�sl<M�u�yٓ�,�S\��Y�41ܪpk�	ޖ(j�������"ń��>��xG(S<��]$��s���T�؄���o��?���~sÃ�#��= ��E�@�����Қ��b��Ӝtz!b����t!�N����ǟE�ȟNv��������� ��.���ZW]z" 5Z�~i��co��5�b���ͫ�q�y�[	����R���%F�b.�|	9��k/�&.����������Q
�ѧ?1��g}䝍�&̘(R�-i�s����5��W���'���X<��1x��_��'DNM@��tu�u��#�W��a	��������P�34އ�`�'��R��I��!�ꆔ��쓁��t�jl$���"6_k��xqRV`6���l�p��Ю+ Qe� tW˿yr���!�/���'5��c�ׂ�4J� �S��G��#��7�D͑�>���`]o=�,�t�9��=R&�MC/ӭ÷k�rѓglb�jV�Ps7��t��1��rF����A�%\��9:�}����g.>ygo��E���|����n��ٟ�~�QP�4,`	y��7)b�[Jpq���1>��V��,+��w�^�l[�e��,�U!�4�p��l�쪍y�-^y{�9oP�E�f�o���*����͆���|���^���X$�^�e������`M�K�x|,���s�}�Y�T�Z|�~��_.�)�j�̴bī1�E�
zvG������`�\�t���Fz��s6��0b��5��9���~�_o���	���?�h�K��T���k����կ��śĀ`BZ���Ț"��wQl[x���	gM~�T��&�͗�6��[+�	}��&�Հa����0�K��=PP*��0^z�n?����S(���1So5S�Y��E���˜I	��avS蒶��ܓ�/<D�����#�eޙ��
M6$�m'�c��݋9�gw�e^ڧ�:5ma��o������b~v�C�{�W}}����JK�UY�
�Jc�yccc����<U���E���9YL��Ւ���wA�e����Ë=�E�����*	��XY2P) ��-��t)8aKj����ж�*�vk�dS��XZ�@�x�SSr����D��Z���,�x�M�}*;�0p��iqjʥ��o�y1� ��G$#��N�d�zK�2�}(��?�|�u�V9�'A��1B�nG6���kD��c[ݎ��Ps#i�b� W ��->M�,?�'�!�� j�a�[�`�8� B�8��W�/j6��%�C���b���mܟ�:�B{�����������MaA��Cq	�k�
���&h(%p��a��AXR��~dM&�h��uR�������,sٻE�H:
��GDߛ*g:�	�_��[7�&1l��u]�W�2&�MXo�u [ �p����d�Y�C�d>��w2����@+(��T�2�#�@ �)cF�#,0 �^�K���5�j�D"����;U��� Egȏh��}��B�t%}����G��27"�0�(���I%�:�8wGd�fUUպ?���6�8�Js�
��)���-�@�ʟ�G�ز&�~T�C3��^��suc�4�]�ɖ�Ѥ{�"@|3��Q�&�~^o�l����x��%D#Gag��n'�@P
#���u
����b� ?���(���13�~K������6LH^�o���"�Vh��c��?����#5�QNiڧ�NM��JwJ��Z�#�񿃏�7��𨋙����.� �l�=�")ox­�$s�����4�Q�t�0����c(��dJuT/�tCI�Z�kP����my���E7����zz�kC��߀~3��>t�ҩI�� ĸ����T{�z$~�*�z���4ˡ��?�٩�,�w���h�m��B
�����g��]Cc�YT#,�f�L����"�<\b�h�͟�+�5MihWTG�am���E�i���a�B�O:	�˹��y?�dc�a�"�Ƙ�,�����&���d
�Ks�i�@��v!��6�Pq!9T��3�U�U�Y��j���L��2�o�1�ڊ�[z@��������S������lz怒���y�!����������#�v��)�A7��ߓl��[�;=��Dy�d�`����@�W�|�!��a%�H��+ȉ�m�'t��1��0�	4��E�^���l���#̾�ݖ#���yaA+]�ۿ���O����a˶�㫀�ܹ�Ҕ�P���7�U��U�����P6�#w��'J�kC7�a|�Z��XS��A�	:�'�9�*'^<31,��;�NV��2#� t��;O���QpA��%q�'2��<g@�b��G/˴uu�� �]Z<�������
�=|��`]W���l]|{�E�	�V�d+��Uw�r��x6�-��h�����*uтj�j\O4�ßMrjrFHJXr�xX�F<�A`K�P�x����ȯ����T,_��Xm�N
Z�Dr�o릱����cݘk�%��E ��:�fek���N\$ ��ҋ{+2^(kݘڨ����	j&�\_t�vJ�Q�@ģ�v�z	Q�$�
�}�Oj*C@�pC�`Ț�'�{��k:<��q��&�$����;�����޽�c��S�T.dB�2�`�����o(ZR5�Ӈ��ݮ:�H$���X�y����j�T��wj
����.徙}���kTAY��TU8����WKKK�� ֗�|9.��t�ZR�e���D j䥁�2ѩ���8�{��p��I��kv� g{�`�l�%H� ���NfjѠq�:�s��]�{m����p�3�����N;��*�%�����1��;[4zT\fJ&��re<����^܍�CB�5t?����.]r���BI8H�i�4�P�W�(�|�3�`���N]��� !�v����q��<
�?����QX��k�G)�M����ԖO���c�K�k������I.FU��=�YG_��kD���k��n�����
�ljh��&dHۛ�#
��֎m�rA�Am�`~�a`&/�$����bs�����0��˥��6��l�!�1V�� Oͱ̥��#e�����\w��A�1��҈�ҋ�|�����K���_'�E��sCﷀBQ}�\�����I�?k�&/�v��Bv�M��2[R���~mo����z���sf˨L+4ӎ�
�k1�J�hٺ�=]�!�
�Y�����N�ꦢ���0���6�BG�)ׄ6��Kq�& :s��U�#zĝ�țnD��k���{$���}���y:�>,&fn���$b�3�F�T�f6?�������N8^ָ�$B�5(�d��c��g�C�����߂�V��
3'���g�U���O^gm5���@��x��#����_��Pƿ�u`���_	���������Qua�G�0��x�������	� ��)0������{ī�o)9��n]@ݮ�������ӸX21Pm��
H8V:���a��|�ۀSl�)�a��`�
3%�S���'^+�4nq��
W�T%@�m�;7�$#͗`��N`fa1w�C��3�/���%�����P)�झ���	[�]^ܾ���ۋF����ə���t������@����)߿Mw�(g�f{���z��1�~|�H��?�鬈���@���V�܎p�}�?4�3je���^�^��y��pKl%���HΝD��ô�(������myl��2�Uf�sޠSS�Tn#ޜ���>��w%��T���aq�0�P�kk���s�څ[	�91?k�]��Y^��nV��s���Vtm���js{����8�yF����ů�˃������X�����X��E�#f4�Yp���r���\�|��&��/ �S��Ry�~`�R�q���tJVVV&��O��0Ǭ״HGGk����0%�#��VRr�=����$8�mĉ,aW����)�y������W./�/ȁo�`Q�f��,��`&32�	go"�?p�y��V�L`ַ� _8L�rCP��C����U���V�N0����C��D����w��(o�.�l�"rL{[���B��NI�J���"�q�S]�s��G��=�(�yi��7a���B�N�6d�ks�����a����;��C��oa�\<���O��s�7n9!��qV�����P]X:R�)v�����
jY��?˱�@�Mxq]��mp�J� ��L���f�2p7�1\�ূY����tY�OX�@/{
uKEJ��^itgo�v��X����3� ��""t�N9���.���A�~O�p:ل8���(�e| ��h<9�"8��B��M`������CuP~�_���/�����N�֟�V~�}(�KuS����)M�Ť���Ϡo��@�Qx��7�"Vux
j�Cq��uW��x^'�k��l��u���k�l�?��������S L[z�@��;!�]J��)��"E'w�����0x�]��kCE��r�vAX盛�o�?��O P��5���D�p��	a�O�0�9B�� �T��iM�|���[��Wl��5�ƌӉo�D�@���)�խ�	Mt����9�u�E���yi��Ņ��V'>=0���#��!�T�5sZr���������mE���C\���w^�K��x'l%w�t�SS�u�Xf`�~��1E\f���si6�N�G�>jTNT�6��ۧ�po��jGGGb����Adsj"�$z:��{�B��r��>���a<�e�$����p���x��s5����!�9���0m�5�.2�%�z�� Z���Pu��})J��̙x����˰:���W��᥽~ry�_�aY��zJ�"�;dj�i�g��Lk����Tï��A��&۟V�k��=��mi�	�N���;�w�Z��J�sv��ّj�>~�����Y#���{���|j�>�������a�UNv�������q���+�ԸO^���>{�uC�#	�@����N�n���<L��V������e�,����ss�P(�va��֜��'�H�/ Y,����E�/��+�^�v�C�<�mꉹ@2���+]�"��~�KP�5hs�,�/ZlUev�=�����i+�^%�G��}���pa/���Ga�	H��d7S���^�0���d�졉U�v^Vq�`m叫A骏�Щ����(��9g��ʾLf*���R��TH��I$�(��2[��G��:E;�+E��X�O����ɰg,,�����#D��{K��;��B��,�Y4� ����ҴO���R�Tr��a`A��Z	�Kg'\z�^�4�;�,ςb�n��VB5�Q��f�'�0��������^�ϊ��	½��˲r��i*�Z*�s�;
�������U�X��:N�����J.�	�Jm�ވ��E���cK�78�Uw���s*T�*/4B� �_����?`%�׮,���P��o�\���}���G�`~��2} V.�;֠7��~t/��p��f�"�����;v�\~�ͯ���#ĉ�\��;�\~㑮,V�p<b�6ݏU�
v�:��\̮��Y��u�#���Lv�	t�?�</�8lM��aZ,�9��1j,�l�MƁ��cՒS��U`9�H6���|(IP���;*�5��%$��䍃���.���Jl���0`���E����e���!$&8�z^���	O!Z��C:t�=z�(����Ϙ�8�"�`p�����ea+K#�������כ���T&�T�[���L&�771uRyn����+���	����l�p�n�j@#:7�w.�ڝ�K��-����S��4!J�aKH��������?f�1����cR�J�tz�,|�+��lq �l(�W��[�W*NwLaThkiYTayv��d�e_l|���,�ͯ^��ޢ�@�ZW�H7r'K��t7&�/��.}�؍#T��@P�,�С'�Ń6������R�g�d�����u�}������5���.���m�Ɲ�qb^Z
�{0���B��}E!��]�����'��)#�ʷ�^��a�6d��ϗtvuE����<�q�����U�1#��
[���R�u�]��
A:����sNPpp�]Ҍ�0�w�lMq7h%�)J|������w�ޥco*7@7��ߛbq�f�kXCԱ^J��֨Z�o3!�d�)P},,�ſ����x�yԯ�3ն�]˹����]Hk>1��y���9V�8h������a��L�̨�Y����8l�	��Y��oD�K*��P���}���)֟ڮ9�ȘNB���(�N�^i�����7CL����J��$��맢^�4ɟ�Aʤ�*�?���@o�E��/�͊˞<yR��+�ӿ��~G\���������_cƿ�����j��CR��_�`'�k��G�w�<�W*�Y�
���﫽�]��@��?�n��n�0�4�C����Za�e̪��8{�W`� ���/���(ͩ/n��P�b�[�}��k�|-��C��e�c��6H�!�,��Ĳ�^墢H��X(M�%�����MΈGFFV奕�;���=���X�IX��a���6d���;��w#��1[�V��<k+��M�',��{	�v����?�p��U )�@Juφ�:6�
z���huê��| �*(0pޝ�[��{/�ĿW�p3a�N����0�fjj��p�5J���vg�z����k US�Τ�rI�:���ψ*���D���j���+�1�d@\��=��Z�=v]�b+�}�?�k�H+3[_��`(t��ѹC(�ϼ�X������ٻ�{��L�r>�ty5�c�:��������Pيtc��TT�"(
̖�|�;5�֍��"ƹ�艫�*�ހ�u~|�}zL���7q�g\mgF��ޱ�@�3,R'j��Y`� ��,Gk�-o:oi��m�re������-?�����o�D6�]��tn��/����t��i�b�#,��`��B~�X����4�)J���[�e]��|�f[�4������F�@~�B�ʍB�cV���~�Nw�+B�zwd�!R��0����_�f����/������k#Bd�6�i��#��v��x[Ľ��}����M&��ߢ/&\�!0\�u��
o0s�Ql�� SѴ�26CJ��J-�(�p��wnH�^��[	gg~)ĀN���Q��?o��b�|�v�e��n0����k|E�����o8��י��h�; W-?�kY�]�3���v��|�����N���p/A�%O�0���^�Yi���5T�_�4�W� sY![U�xO����9Ō/�>Ü9@��7Њ9���2`��v� �����E��y�o�7H����?�d���[��`�G��������: ��1xZ�;)I������b8W5�dW����L�#���TE������<iψIg��w�Z�R� ��>?2���!O�o���3��d����+�
�T��� �YX� �k5��Y����eh�%8��e�L��^�8U�[����RΗ඗;�F�,�DK=�K�����SӇu{�(�W=;���;7p�f(��ynk�_��<�����9�+���flHI5��.4�)J�6�4da����u�rww�K��,//�
���]q��U�dQ���Nv�q4c뀱�Э��"��7���w7�S���C��A�f������8���#9̒@�`�mh 魗��-t���E�=�ܜb�7����)���=�'�'��&�_~%t(�����l|4�5�;mm����K��p�E��_eÝs0�:�Ւ��Y�r�䮝�j��������Ty��͗��K�ށ���Sg\i�O��G�s"�E��Xa��Z�e8�u3�n��@G�^�I N����*>��蚷�1Q�FLݝ��%CVs���'&e6����oT���cSb勳� Mg��6y8/�Uf�,���J,K��ݨ�jY�z�%E�Ӟ��;�%A7dv3MfUG�ni*#�
CԚϏڀ�x���b�����	���p��]����m��_�pt�&�j�L'c:9RND�I�L`l;��Ҷ�e���Z%9S8/�?��j��}�Z�H@Yg�*�G�<��?ȗ���b7����-�O.3��JB"b�U�~Sj�����<s�ڸҍ�6]�Rŵ�ɾ{�l�>w_¥��x����P}a�4��WZ�3��TB5$AF��W>�3��l�ݱwi�&~<Z ���EW.'�o;����4��g��d��j�p�����HV"[fff���/�aG�-��ɩ�ʉ�#�Sf�5���O��r-�{���t:T�.]X��R�b���?��΋�nooW���5�̜ P�τ�lT=������~E���*��1�`�ҟP�^7������g�����\�!-�{�o�ӷ�5O��8JZ��e>Zo�Ӫ�ԃ6����te9��B��tj*�B`zr��c�0>��}�ǻ��sL:?8�����u/������d	Ď�z�X�;�������^g>����춾Ɯx�����\5\�)c��7� ��������G�U`�
-��zVR�Oh+).��M�@.L�#�MLLT���*���"@o?@�ܻ�����V�����ϧ2�E��H�I��;��G}D����C�Њ����o�g�y�&�*I�*,rZ�	sI�ύt`�>��Ϟm��[o8YE! �SR	�*�׃��/y� v�2�`[�ƚ��$��(p�7?\�ɾ`���3-֝6y]��Zځ\c�8/������F�zJ��c0�N�,�{�z��2�Q�0�q���Tؓ�G:����Oܜ��k�8�@K����h/��bL�ē�[�me�0��}RJ`���-���sQѹ�Oݺ{*T�t^t5�T|zJRj��ʉ,sb?��T׽_綍(ܛ�j���L�kH���T*;�6S�l���#��[b$ ��I)0��ውR�?9(Kw�
B��T>�L���?�S v���k��I�TlbjF8P�4��v��14�����[v���+��k���8��R����P��_���h4�#i�9���IW�&�N�Ɗ"▛�"�<��HO.M�k�ԉG��I���=,�TD���n�Y�G&~��;񂗳��j�-~s��?���7�'���7��8�Y7P��h�,�K6�%�%��D�C��O`��L!��6��d���V��8����B��8��򪢰�b�i�i�L&N�u�$�a62#�`��N�i���7�G���]� ���؇\&0����_�ϱ�^������������}5kzΙ_g��� ���Wق�}U��f�.܋�p"�w��y��P�~ۦ�g}_g��n�����&�m���~��>L DK3�� m>0!��Gw�%�_sV3��u�P�l�ٟ��ͷ�x�,v�GV:�{"'櫞�T7Z���D���^T�'�Ɨ�V>�,�/��2AD���¬2�{�rPf��e���bn�j���F9Gic!�ɓ��o�ic��,g/KD��E��@�q��� �8ƾ�g�\-�Me��TV(���v�Ut�Cj�c�Q�H��O���'�V�*3#���+��W�:��Y������jX:�[��p}��e����\+L��vL�ǡ���-[c����@A��2؍0@$R{�">AҲ�Z��r�e���"��/b@���`���q3��骹@�e��w��2�����l���.�y2��S������A�,�m��ڗ�S���'e��Axl��C{��kim���~�ʪ帞���3C,v��S ���0��!I����:�����P� ���%1�n�͕D<�-�SZ�"߫f�����GQ[l+p�)|��~O�.���O:��i?�H��fP+���O~���2น�����+��[[#��2��F���'vgpJ�N��"���<|D��Y��(��5W|�6AC���!tSu�5|�+'<�����6H���tϨ������Y��?��:8�d���={e���� ����]H�W曈�! c�J~�mՌ�ԕ]l>�߸�#�	.��]!$��wǂ�"������@�iY��j��c]e�!�<<�u8~��~x�"Z
d�C�,�l��J�6T w��WrҜ �U.W�E�����:�x%E-���z��{��S��G�3�hN|:�g��Tk�:�)�♿w���Z��f	�$�S�N�qhW�v�Ŧ�͡��o��mx�.!Q���������8�
������{���w�Oj��'���T�9�B�����E�:��/�{g�i}�g�/��?m|�	�əŶ�����Gc5��˟7��k��=s��6�.���w�lK���V���C�(H���K~i2�������V�ϯ��zy�'o�jw���<�P�TP"[���u �;8�Z;�::T�G�[~Wyv����9�ف_�p	т�;����W�H��p%�G����Q���EPAZ��o�j�*�B�x��Iw*�z;%X���a���M�b^j ���S�E8��L�d��%ĊD�����sX���k𻀄��1<d�'��=3�A�#�z����j>k��{$)Fh+X3�_Ce��]��AM@z���<B�xKI�Xx�#"Kc��pޠ="���CWr7^f�r�&�\ ��;�z�IX�D�ajn�t��(��E��#z=�����w��Q���KX
���o)n���4˦����ꭻ��y��JV<E4ō���9l�-����TVN����>j�hH���{���A���Q�Ұ�Z�!��Ȑbj\v�ۚD�r�=���.3ŕ>~��Ȇ����+�}���bhc��(�7��Nu����F��yP����%��,��ІDE������D���L���P�U`�6Mc�UW�oZ��̢B/��i3�qX./Mx�Υ�ƶḌ���ڦɝ_T����i���g���$\�_��h|aڧ)�?�g��95��M�8�T����>B�Cj a�;~�)���}�Z��d���Q#�i�FmX�jZ�#@�����츖��R_Pz/�P�T@~�H�Ix�a�?��X$�Kj�Mg���ڵk�:15<a a9a t���w�QՉ�Sjg̏Tn =��֞vmM#�_�����_��`/aLL�\8���Ӄ`��@���9�Ņ����Ye�mO�l*�]x�'oQ��<��-4�ľ��ե���)7@#��/v��⒒z���h<����������k^Y��bM�5=VcE�&�֒o��"��N�`��?���H������m��2C|�n���Ë�\���̳iP��~-/�w9纕��<�f�.��OdP e�=�7���~��KSD[���1×�\c�r��f�;5�Q�V E���w�b�j%/�Q��/?}�O6p��_Ɇ4�gʑM����ƛ��,�ih�^�u���/�T�qP�=�fց�丸����:G~�Ƥ)/�%��e�4TϏKu^!�ѼKW-���<���2m��ψwL�)�������,�����=�V�$�E��΃�m;��Dw53���ܝa�CA��������wj����ȇ���	]QZO �������3#_�N��w��7�a�z]����	�ࠠ��ϟ?����	��)��j���$��U-��AmJ|���m�G��,�p�#kr�����ˁ%ʝ���lA�+$;ʡJ�*�����ǟQ1O�Y��L�؍�5�9^>"�H����0�\t讃miǿ}V��g	!l%-���5-��[@v�������*���g)���,1�(��i�d =�(�{v���DJ,��A��׹���Px�gڨԏ���{�[����h�]�俈��~c�ɩ����="ԟrb�%���QH�����V�z ��c&g���FFF}!@Ӵ�],�w�"�]R�y�L�a�;�p�'�Hq�����Ι��k�����&挱z�S��� n3 0�G�	�0Y��6�DćPb�O˼��N��ߖ��u��	"|����s��O?�	r���<=>~	S
�C� �� �XA��"q�B-�HR��΀��چ���
���}%wOE�ӟ�L�j?�1��[4;��2P�kl�ŀ�HP��G�̙`�DSvPÂ�h�Tא�=�I	Xnj��{y|D�'yflW�8Zs��R�.HA�|�yN+(e6��h*���(��d]c��]j������� �'���S}e5CB��S�� g��eM�w��A�i	cM�_���3wB�5����:D����Y뫕[�KJl/qo_f�[lK��̜�An�|�in�(�Q~�c��f9m������O�+�G�Z	o"c��"�[�tPkY�L�U}f�4	,���:˒�Yb�OXp�<$k���2�;}Q�>@�PjR���}[��~^r��Y~�΃�Nv)��'���~��{���u�3���8�0�h�2�oÚ<2_zؤ�Oi�����SuV޺;��5�;����3��e�+�>�5��3�.:Z�t��%���Dqgg���Ҏ��j9���,~�^ ZDI%�37�|�_��|L ]s��Q}$�}I��U�O�7)�݈��p3�����A�wD$T����`���T*綽gFvF��|�DFKK�Bb툟 �KmA���`�,>+̓�/ׁc-���C��^��w����?M�^���0�Ը!��[P��[����ڹ;�S�yi�I�8��;��� [��CPF�u[��������aP.-S}���4fnz�5��K��]��s�������f���ڐX��u�/Fk�@qBz
�]�`lV�n�m�:�[f(��ù�����\���]0��~^�37"
�@���ן�΀U2�⮫u%@�^ P���'1hEl��o�%�$�6T��YBQ{*�Ea�Y�������{ a���npj�	��넷�/5��)�[�z�$J�}�lQ��L!�}���ߨu��J63ǢZ��g6{�^�i���~'��N�:�]����'���o�U`�{���l�����qcO�>�݀.�e/N}�+�¹B@���6�?J�T7��y�* ��\hY
�Ö~�E�#��1L,������2*� 2�d������@�07Hf-KҜ��Bم��f�T��^�� ��|���i�����l\dkɭ��p�'�Z%@�m"��|�`�?������h@\PAr�@kX'�򧥋��*LrZ��If���8���J��L.���I�S��Y7����#:?�:�ɬ[�4�&/	^9j��S�8�L�`�A<���eI�� T��C��ޔ�����<�}]ϼ�ނ��m+ùw�7��S�X���a�(���b�[a�N���h������i��H��"�� �ςh��
�a��������5�@,Ő��ݥ����Rw#ŏ�1cu�|%��ږ��'|��H>���л`�X������MP��5~ĝ�q���[A�*��	8�6xA:5���������u�����o�:{�K�ڊ�m7�\j�]��!�]%���P2��Kr�M��"�M�vkQ4(M���&]�&+CaL��eH	�眷�����k��s��<���������Ґ��K��M�$��Aw���i{b����`��@-���q$�kq�e!�b���6��4���t�������_�ΗFVg"6S�װ~Ov�hY��?�a/@�|���LFM!$³�#��˿#����332���o� $ j�L�{�!�z��"S3H�T�K_.L�
�vg��;V�Ul�{�\Cgv��!�z$��Xŷ���⮐�v�+V�&�v���u��V�V�N�{r~� �x
hPKR4cC���Ɉz
������Q'�G��J_+4A�\V�e�ҹ��D;w������OY����@jF�~aKw���
�X�R?/T�XH3�5���L$�#�(R�=�.q�?
P�_�&�2�a]Q��(RH�03�~V�{��6����� 矠����I��|�X��Xо��d&/��lc���ެ'LG�%��z�y�����W[�S�rj�{F|�o�W7|��jii�-�;��G�9�@Y^R��yx���Cg�f�#��:O3��kb��H�m�`Ψ����u�1��9���(��npKV�+c`��I�*�\.ٓ'���[����S��D���H��#`:=6?ڕ��d���.6����H�$�4<�m���7�t�,��W-7�����TA�7��i%e���[�6Az�J�V�t|F�	-:��R0�$�(�&S�*�B5p�5��[x� %��|�C�K���z%s�
��0{RZW���Y���k�S��@�y�͠��!�'�%�b���}�m׸���߂k��sZ	�
�~�ȓR���G�TQ�x�/n��,YJ����;�DZ�h}}����:�t�U��ji��_��%xÆ�����hZ�B�mj�]�h�U��r�^䠘��2z��|����Ѫ�����j�d_�n����WK�}�����'a*��E	��9���VVU���}�#(nK��"5�`Ah�U��o���1/�������"�I��}�T��8A�%�ۨ���|e���%��oq6��|l%��+ӆ��ž|�޺�њ'L�F��7���S��[X)GӤ��ܲ;��:���m�L�t?b"l����7MWԉu�0��}���gtRx��ѵ=+Ge���po
Z�D }w5���q����� [:����?��#t�755��:U��->���t���1���dYXm�D����|�� ֢��nk4�@�8��Ldk���N���V��N�����:��H��=NdU
{�A� �Lu�|ŋ��������>�>��Q��.1����;�z�Dښځ��+����+#��y�5��<0߰�H�ڹ�xT���ka�ͧ=�rU-C�1��.���]Ƙ����#��sd� ����<JC)���v��5��c,�f������S�tDai���?dS+��-�'����ԉ�R��r�e�"4*�����G7�� st�o�#4�揦��U�]�wS���(�ܻ� VTGQ�ea��OeБ��?���`�Q��8Zc3�{\��1p�_�U�)�	Y�*���:F��}��)���IB��Y�����ƶ�����@*�Q��W���Z�T�_�xa:���g�)���mu+�%��@�;A�c�͆�;xo���b���c|��96
�(m
la��2ާ���)�@�S�������Ĝ�5-�ãr;�ܟ?8��2����^a@�ru~s��0;���ի��H��L�	�'@����&�FcZ*�詶	].���,Sr�:k�>���s�S�`z';�Wbb":�YA� 2�����ʗ(qgqF�́E�h�N69�ri��P93���[�/��BW�@L:�Zj_�^E��o�X�ʅ���V#�Ɠ�y�+E�A�Z��c��^o�=߰��XA`vbD=��%0�:%�S_���gl�]� \W�ŕ��J]�ڶlҦv���u��C���ZrBT��=w�0����۫]�\H����#,���GO.(1�����C�	iM1�jM���9��9�w_\���a0��Ӗ��Hti�.v4�b������#b�I����>wa�貈��w����[Fi��OO:�wQ(-�����.�*�p[�fϘ�?B�4-�]�-#��a��s^��dGVEch�>�
(���W@�q�L���]!a;x�P捊3Q���x��&sK-�Xl>g>5���p[�ߪ�Ӡ���ʋN���TQַ�0�3\�o^6�Y��YI�#DQQ�#A�ԁ�(3�zmkFq1`,i	 ���%9�F~q[��Őa�����Y �� �y��ǧ�b@Υ�;ܣ������Z�����7�0H��iK�OP�Z�	2Qr�in��~(�w��k���K�09re��f���.9�$d���H��ɱ�'Ն~w�y�V��.H'�Y	�G!�wzݗ?��5���������T��/%W�S��TPi6��'�T'���F��݅���#�	�_Q�ָ�xi��Ps�W��h@�)�{h�whm���zuJ���ܬ�0�]^c��9�o��]?��i�~� %3 ����v�2��I>Ƹgl鷪��g��(VL�Ku�_��Ϯ�M��T�zFa�
Q��hP ����ɗ��g3���mlfڰ��W3�!����c�gT��H���Ooo�x��AȾc���b-��7.H+O.v,���N��㪻h0�ka�Ç�>�����y�FUP���u���В;�!�N�.�
�T:���	����8�u@E��db�¸XWGgj@��N�U����;)e:�u�8��oe�wW,;u���Ө1���
�)��0���7���%�";J��,�,�6���
�x�A&C1�n�I/�0?�mGt�:d�a���V酉���]�[M��Y���y�>�)c����s?��F�+��V49��a���w$V�j�Z���5\�jv�Ü��
i���hٟ��i����<��^�����s���J��]�l����tE���{��)�eG��i����1��`��I��(��Wv���>��Z�v
�HA�Œ�hS��Aȧ���4`e���;_��_Z3S�C�d�Ξ��m������0�.�����#�f(|{M ��T�Z�Q��{�/uȌ��I�!uy)쀬�B�|G^�9�E�r��!�!����N�� =�v��=� k=��f1 ~�*��5ioksKv��GH������|N^ԙ�Ǌ�`X�� Ai�O]d2~t���4$8�%ga��v��i�R	J-�+���q�s���"���u�u2��C��Q~�GC��5J ^�tF�3�W�VF{P
�3.:%�=_p�g�bj�6r�ܬ$�pN��F��B}r�>)��?L�n�Q� ��p|"=�2���E� ��Q6�	ɳ��M��|��o!�*���Ѥk��9���qJ�iK�!����ʼJ�	e�癛��u�$�P<��������
jg�Ƀm�q�hcƨ-�tHS�l�?��5$��\ȱZ����gؼp�"�oԓ�_����(���j-[��°'Q�[h⭡�u���@�҅(�/�̤��$�ѐ�8��j�������Hh�Ը��%��:c�Y��|p]ѳ"4��t�/9�Ȳ�L~U�`l?�§M=ى���=.�nɊ�x�~~S�A�)��	)�L��3���^�i_�ZO��wl����!%�n��=��x��fy쾵K=6�C�J�C���_2�h��p�Tx@.(���G�V�{���9}�m=�!���7vAN��	�"]�4���C/�-��VF-v�]���o���YD����|ބ_P��]��/}�=#���9�:�� Z�h	*�ĕ\�$�Y�zH ��։/8=�H�a#2쾆HV'����u�胶g]���̍�xI�!z��Kڻ�uB�q���h|>��"���<2T����a>-��.�?��=��S��T^�ۇ����]j�w���ť�(�Ԯ�3sD��S�>�x�F�.��h{g��f^r@!\^vgp�'�0U^��și1���j���nI�*�߮�1�к:G�'�3��cB��N\i�`
ŭ=����P��!���pg[ ���N�@�\.��h9DGSn�M,%����D\;�
'&r�/�x���L���^ȕ#��^ˈ�O�kz���\�d�P�_�pT)^[�
Uz��'�D!����Ј����9ROV��ݢ���~��{ٟ��آ*p�xϩ ��c
3�/�4�A*��wAk4�W,=�����<�!��`2J*��!�@�b�
�Ə?/e3�! ��Ͷn3���[WS�<!>�0E�2#�!-XH��~tD�
���mޢ��f��O�v�l��<�d�i#�jM�	e�X�rL�#�X ih-q�;C��6��m9
�S���״T�y�:���βu��%��W�c�����`F"˸���c4z&:vƧ��m/�\������i�Q��o?s�_Q�P���V�9g����eG��/���r���{/揭��w�Y�l�9NM2g��ymǘ�[c#�ё7�oDG�X]�H�"��s�Y�	���T���Dev�q��Ϛ�Ɣ�
2���I H�����X]�`��rp9��?�)[���"u�R������v��R�_�"M K6&|�{]�Q�Ԁ�iP���d3�����
Ъ���G�:ѲL��i���v΀���c\�8@�@�������S흒�-���M��}�h�@�P��Lsǉ��@�Ƨ/�l�M���	�hj�ܹ���:vfW��{A���c���'��T�Q6��*��@x��������=��>Q)jDc9Ʒ�[-���x�c�S\�k]T��>���$.��(Z�q���s4-Ɔ���Y�r���x B�%r��!�S:�?k�
��-0�c�O�&����� ���O����&Hy%.��,:m��J�xCW���x�០}in8ȃ��	��@�$@�՛���[�����:&���;D�?�n��P�� �k{0 �|;Ϭ�q٧�0.0���='��?�w\O~��;�@d��6�Rd���!���lH!�m��9n�Ĕ�%_�qH$2�ᇆ�<�L����m����G�\�(�9m.�Ml<rRMt�˽��{����8�Kjg�4�vB�µ��9��Z��g��w�ƕ-G��)�v�A]WQ<�6R#8B��]=u̓�G@����e=C7�/3� �ė�s����
��9!;�K73sQ�h���f��s���8K�Z��ݻw�8T 7_�6	�ѐAâ���w�!{5��z�	�n��2Ch��.`�0DY�ה����HS�j�-`���8�ܲI ����������xT�J��54,���[���HcI�Sr�A�+_���-�	iXK�ڠ�a?�گͩx�8����m�u�k�g֎���c�w�d�-g�e�w+�	ly������
׼ ��A���A�"IJ��;��>QU��2q��qS���J�u�@�|��D^�F0��f��HuJ����>s���9'Ba~zq�������"�3�b�e;x&!%lk���\��ۏ���YZ'�����7 `��(����w�wG���6�]�#4y����-���_УV�U���p+L��@D�1��d��tWs"���JU�.�l�����h���ϟ:}����-8ܒ:g'�����$ݜ8�興w8S	CW�f�FL�r7z�&����晗OX�sb�o_�ۮRy���� �	�pEEeeT/iMtS�+�q�����c|}�sU��m�����(H�\�[��M�]d�5����b�5�]����+Z.w<�S�M�2�(�*N�1�����h��P'��������M��ȑD��E{
m(�#�o���i^'狎��ks|��h��|hrmC{���o�������I����nx	���ݹ�v%��ճj��{��o���&����3K��x�R��0/��qe:��v�PD��A�|8��{�ft3���lr�щ��!n��J�w)}}}J�nJ��}�R�9��#�@�{p�]n��T��5ϛMB*~�M�|��ZY���u/��߲�_�Z�^sIh��JeC���o� v �pM���5�
�c����z'��~ym�׋�+�@@��/CG�b³U�%b7w0���C���\�)Е�|��&��k�e�*�m-xx�]ځ����3�n����t� �u��K�*����� �}��o� �¾��\Y�yK|	�z+��z����r���=8��j��N m]c����R��V���d���'p�s	2���6��H��9_����Ge%�&1��k����P*T´G ����vn��n�9��;���?@�Z��ܪ���T�Ӯɣ�d�(`9O�J�X��W��9�rǪN=r���Y70�5�+Zx�O/mN[���#��.����8�v��}ϵ)ٷVf�Ǡ�s}�H��f��F��a�@�Id��Ӡ�����G����C���D�U���Є�B�D@!��QX.}�Б�¶Z�m~PK�W���B����d����'�0`��T��w��\"�������&�y#�i2�������c�*�Y8*s�V��㕿�jRl̳$�����D��S�SU�Gk��)�.�ۄJ���`�9����zA��G8��� �G&�$b��9�w#�r�׏ʚI���9zB���:Z��2��~L`�(�D�>�Ԫ��_/K#@^i�"�#��
�&��6��{�	*���H=��I��R�kbЍ�y�)�84򏟻m�⅄�ap꪿�,"�/��M�-��
��O��� �*H���0 J��:�7@�"rr����7�/pOv:�
m`&�&�c�pa�I��mG��x���ԉ�p���
���5_֮��t��9�� I��6��7o>�@p�NM���`�zd<�߶@�T{\Z���XHP�%��u�7�]�9ҟWƝ��Z_�,y�ie�\]�}���m!zPe=�/������m�W�����t�-:a�G^���0{;�5��W��1˂^tޟq_���wlA��{#�F[V�ҹ-N)dGF*Ȩ(L���}^�	�����3���W`bj@+6�^��,�xx�S�x�;��l�:�v�L��@�Z�dǧg�>�T��_�í�tw��?3�GD�*�,p^|\U~^ }��h5���	z�PR����ɳ��d�+�.	3��{��A$�-t)�_;H ��h)����*������ԍ�?G���;hai�0��*O�L��\n�0v��۷�x� ��˹rg�s��/�ޭ��+��A���)����`�t%H�怪�o�oF���G�Ңg�$%%UӨ������U��x�%;�P�}ݱ��'��9�y7�6D�n@U�A��>(��uߤ�/
S�WF2|��?}���l�����Հ�7K72��(��w��Bt�/���8�a�ϴ�W<��Q����n��� ٢�S� z�%�ː*
�������?����6���\r�V5u��A!��� :��PR����G��X)k���tM=�I�$'�c�yИ��]�KB��|�]��5B��m�m��*���5�b�m�|��Æ��+ڍG,h��M���r�O��RY�Zh�M�@��,��G����~'��a�F��Ի������
GB�jEq�#��*-�T��Wo�l�2c)��ro��g��|ǚ����W$�����J��9Bc�E��ָ �X�X�x�Ω����TV�~hM��MN����'�B<�Ğ���I�%��"�d���|A�C{kO@,�T�3PYJ�ڷ'/`0�	�w��M��-�׿#��Pt9i"w|g�����}��H/b�g�i��]E��!��z�W��Ya9�5�{�e�.vqaT��`ٳީ�b��y	�y3���;8�C[�}̩���@�[�vP�]*�)Rf�a���RnM7c�����k`�Gt����e��h�L4�["�z��'��n�; [UlE��q:{AL����>�B彶���Lmk|��ym�ď迊�7���������e�!��=`?1֠�� m��$;��BZ�h�g7�����ĭ�EAe�n���+���
&�y��իj|��(	��b�5��B{�g^�i�n�(���smD�qvno|����KC*�M�gcc�6~�4��I}ڌ���KlP&d�1C��
��;�/����4�-�U�t�t�Kp��:�%��zs�b"�w�`6����_P'}v�w��ڠ=#j(�)N�&�S8�����*�C;���r�پI℣i��'��h��:��.��i��˞�Z�3+����>��==
�R�F��O}���E��ND�*Zڠ}5��-�ͧ@s<�%�U�E&{ OBHѽc|MJ�I�i��m|:=C�<8v^��P2���m�o��n�mv��&�<����,Օ��סʃH�!R���~+F��{�^�Յ�i��
�D2S��N�A�7���xx��;�m^��'��d't�BєqPS��:�3 �s$���1^�j<�Q�	3����E��+�D�bҩ��Ԧ��\;}����M ��'��?���v5U{^�W�`pd��/�ŏ��n4YgŢX�xV��%��h��채2sy��g�>���7�N�S��=�ro_��k��4�v9yO�uvr
������9o�:#3�*IM����9�]�C���C~rwt9�d�'�钠��Y�K7�_f)L~����ۤ���w�Bͮ9Ƕ��Q��	z��c�OU\�yU}{,K��5C�v�������i��ڑW�%;gƮ�H_�q�Gqh5��ؓ��p1'u�C�~�^MLT��!�+?T,o��?v�����5���C�e4�e��=3#?��=��6Xix6/[;g�WH�$R&ZSߏN�D��+^��;�3���u���e�'���`&�m���oB5Qh�D�jr[�����'��W\���&��h��m�5�wzx�c�^��F~MӘqzk�z�9�,~ґg���G�9|_c�[Ԡ��+D+O�D~��[6+�qS��M��FJ��X�؍�C�YrK�#T�UL�
�M�u��΁��hC�Nۈ�����3�@H�������wɜ�,�[���a��M�b<�܀�H��p��o������({�+��B������mbpk}���!��$�GE�2Ԉ�,~��k�E�Sd��W###6x{UQbf~~>��u~1/U#��0 ������r��o2!X
!R�z���	���j��?��C8���*��0s�M]4�;�/�BU�2��ߠ���)e���S�y<���Dj��L�g�Q9�ӟQ��vi�q�*O{W�>�`*r���q�I���u6�Zę*��u��z�ם9/9�4�l�E+�)/<i�{&6����������(g�����-�6� T�5=8j��D ]����{i���f��Gb[�����c��I��	��SOC46�D�i,4*j�Z���^�������Hk��L(��"��ڔ^�	�ƺ;���m�M��������R�q8ףm��N0Ζ����@�L���\�xAV�j��*>�r���/SX	Uo�8�$\��@f�q�oB�t1�K�s":z�J��}�R/K�{�RU6쐈/.iS!�?U��pD�T��XV׻����F�(�R��O�|{�r�����n,i__��jT
_�}�hZ�A�&�Pg3��V�
!x���ՉCFRw����<}��̖\�1�����8�/f���<���)�D.�X�R!2�aɭ-@ޫ�nd�����JT$1t�^�l]�]$�C�
Z�LN`wB;��2;Y�޺� }�P���d��j}$ґs@�{fW��T�N{��S	��� �S_��+i�js�!�M����*��m���޳��dj6$�np�;=,�<���}7�@W9�vĩJ�罄�1�{���7���&x�yԘ�7*꽺�?�4~��W���B��$���7o�,����@��|��[��c�g��~�~CK�v��l�w�j(G�$LWzvr#���)���E��x�MH��n��zC�4���G�iي^ǂd��O��d7�j��"�e���h�f��j�B�m��!�K�U��;#�#a'�j�*�0��ȯ��׳��(I�p��mM����lՂ������0_0�t��PZN�8�a%�_�
r���j�8�7�?緜WKpy���S�"�If���i���S�S�ހx6R*�;<��5U�z��tq������h]�)I��9�Ӱ]8�e�e�M��M��eO�^A��>�:�[=+�d<Zop�p�P������SN��.>�M�������*qA]t{�ɹ�$���:�N@د�`���{K��#ϲ�t�s^�F���%}Gu'{�X@'��c�{dV��'h�cd�&Fٳ�%�I������L��gBKZ�����ai؟�}�+;�?��dz_�Y+�j�[H��M`��\�S�U���vѩ�H�c�)��k�A{��h��S�C��z�Z���hf�T	␭�`u�$�D��ˡ�m�hL����-�����W���[kP^��(�����=�����v{�/Q�����yhM[ܭ2�S�zw�y^x{��vT���ÞR^�TG�3�'}w�a1��>: �N�f��s8S3���NɵlAG�(�f�C���HxZ�2R��ц�����;:H߭�E_9�{X��H���Po�GE.�����#(�"�^���ŶO�z��/��9���u�.�Y��yV0��bj5m�4y�n��&9�����;WT囷�D�7��B1�����s���k�Ӕ�"Ϥ��uʋNU��k� ��1����;3���D<�`:�[�7K������C�E������	��6���W���;j"�1��Jp��
�UT��!4)|��?����_��D��D��ֲ�7�fe>oL�Voϓ����GiJ�=nCv��y��ф���Ԩ��W,=;�������EM
�{s����S� RG�{U�{RU����U�V����I؛��w����N�� '��;�x��3�v-�C6�ɕd>#�s�lL�''`.�]����t���w�q��E���Y���b�m#<��֭R��Y�o�l�q<.�]4�o��w��Cќ�������I Kk�ǃ����qܣDZp����n�ᚭ[�ą��m����n�C_塟�ۑdі.��*��dv�6�r��c�j�rt_�z���W�}�2dꡫ�=Ws�Jp�BWd�Ѥ.��3�ɔ[^ ����h��mnX�K� ����D�
W6��es�:�yz��k]n!�� �q�N�<�0�i��8T�ǘ�'r��@1	q�a������3RhFVS���s��׸��n��=�����2�C�(]����mZ��~�c�A#z�vptt�#*���߇��m4�_�QS&誦� ��-�p*�#�˟��K�kh^i9d���r?B8=*6����$9�յ�z ��&�I����Օ��˱#�<�I��O�k
���rձ��;��Ӟ�)�NY����C����K(����ڠ�Gb�ϑq�U��8|0à=�R�,���=�!�Y�M�XtJ(�h�X���h�^�$ONJϥ�c?�����<��O,�є���`[��?�<��� F�vl�&4E��p�y���Э�-2����%��k�L��"�ſ?�-ɜ�&r�?���M8��M�A�n$���7ԧ�:��z[vS;�\Y����׬^
=P@���,�>��L�X&�_�Z��Tu���W�3��}2Õ="7��]jzX�v�	M�(|o�O,
x>��L���aƔ�H���
�ė�\�;��W9���O�]��Cl�=�5�� ����}l:�+]]]	~� WW�%�3\�AS�"B����݆x4��=�#��0������%}�G4�����C��
���&'������o�OԱ���h���r#�U�@>��h�����(�y��� k�^a� ]�ӟ�~��˰����Q�^!�����0@ލ<��o0v��$���4
f�0���d����fM}��8��n,�)�ŧU���� lt��y�3~�頀7��9i�c?�2����Bȴ�7�H�#eO!��"��"IZѠ�2�_�&W���7o���3��x&4���Hcdu���� ��G�߿OV:u��!R�!�bChd�Oi��|��	lL�#?�XuMP�O؂��|>o���=�s~�%x�+'u)�:�$l�o4{xxT�`����{����24�w8���|�K�2�G?;��	8���nN�������^�|AHӿ|���l"jz�K��"��W��@����O�ɜ"����Y{m9�3J��&9~x�"SD�h���1~1��2��4�����U_H=�$��/���/��3j*�3��*7��4�J�.�|/��K��.��7<���z���~RuU����K�v0ޢbִ'i9�rf��g�.����A������m�8�=�(�!y�!���hᎼ��=fs@�*;��.�U��fS��~y(&�<N�I�ܴՓ8�>�f�Rb�%hn!n�A4�wE�&z lEcĸ��w���@��H��`a��W�n��0�C�$	��5�~��C�'�ji�}�v�xIa
)�'ZvgDՁ�&w��B����æv�x ʝ�٢�c��6�O8vN�b�0��A>���|��3�",��mE+�UO}{�J��Ҥ(���{<��@9rR��L)Z��q�L�H\�����*l�_`�V̵K�+m�f�e���h����ÌM��J�GR�w}��\ׁ4��1��W��C1D�pV>���p��=��:���T��(N�5"�D�}��Xxl3�4��ox��j'{��?��ag�����sT�����n7{����k�M0-J9*���l^Z��_��}�˗�'o�%J�Ю(��cSI���
��6�h� ]��{ܗ�&�~|���:��;ft�9Ry���/�5J�E������VM|�$v���S��@1f'BW���T�k�G��͞���K�P�� �Z$B����ۣ^	��uD�sKT��}����t��DS\��t��8�2�W�&�2&|����9�|�:{�Z\O�LLJ�1G�Q�s�\���G��'�j!n�(Q�,�$�<#�y��E�B�RW�DH���>.;L� �p0+x���\-D¹Â���9��b���6u-�#l�Q;q�����G㶚�Ł`�'2jԶ��
��,H�T�9��/\r�dEL~U,�R��Aѡ�7��%r8��u��D�&�-���ы��#� ��t�3�d�%��{��a�Uh�(��8A.7i��v�)xޫ�7@бԈP�lo����8h)E�%�mW�g�+;��th�x�]-J���Uj9{T����P�q����/t����t3����&vj]7y+_�=0�R�s~	h ?�؛܀KQ���G�Ll��|������/�.�{I�@�ܳy��uاȀ؀�6��}�ҵ�����
H�(n���{�����ע&��j\�j����$�~��|}�=�rp!��@OS�p�@���2̅:�e%���%��B�������nD�k�,=]@���}�i=L��-���� �;�����wH�����Fo�t�736�ʱ/��MLG�.�=��r���s�(�߼qꔑWK�l_�f4cn�#�e���k�����h�ɗ�t�w�5%xFxM����j�����&Z!��AX�tA�`˛�1q���^�X9�/��i��U���Ǎi���3�/$�6Z&�<#+k�Ͳ�ծ���=:�6���+h����;>�v�L�!�S����Κ�(wlr�z����E�G���{�ծ�y+;0A���g��><��&	�(���H/��J�F�$#Q�&cպ�Ca���1�:�2}���>��V��o�n�=u��O�6} ���>>>3�����f�,�`���"�B;�;~^�J��M$-~�~w���=�����9��\����Y�}!����8s�%�h����q}����(�6XM�mMie%�n{����r�M�щX^a�(�6L�n0�/}D�!�)���8e�Gn��#	�l�{\%Ϗ�� s}�j?�m$U�t��c�ܩ_ �^�L��y(�p}l���nz�R�iU����HK��ڋ�C9Ż�0��E�q���Τ�%�h}~���Y�:0֊���X5l.F�G� �s���=1	����91�L������44��D{��'T����Z��^���`<JQ�+a�!��Ρ#�L�`���d�]$��&G�<%	��FMM���Ĩ���l D�75���nBkt�:B��'����0�>�;ohhz�'x��d鯩=F�����]g�K5�x�^�ul�ϣi�9�*Љ���W�Z�ć7���nu(fب����W��X�l�����P���}g��.y�\�Җ�C��zn�T��ccc����2�|T;4���C_��'CB�νV��3T*������|�����=f������jK��B��hZ�n�ki�.�ѡ�mgFބ��T���LӦ��)��_��s��r�n�ЀΡ��C멝zy�=��Ao�����lg��N]F�g������R[�[�:�?-/<��{`��i9�R1��A�<������0I���V\�:i�R��T�"F����g�'x��6�g��o������ڗs3#^{  p��+/�h�8>�h��a֞Pb�.Ȫ3Ҟ�X�q��-~�"{;x�L����[F��kuN�^��Z�M8�fה�OB&�������t��z�:_r���_�����3���S����
Y��;M:EK)����S�Mm�^;�~[���.�nE�0T��0��mO���ݘ�b��.��/�%䦣2���w0b��������?�o��H�K�jy%K�Τ�k�'ԳF��`D`��g"��B)3��ee�34����jMiv��W7����h�(�PZN,�ptd2)�(�+�nv���X����=Z�߱v�
pf&8�qP��o#F��$6�Y]�Z��}��}��I[��+��xn)��hC��9e��kߧ��U�0�t_;��f���h9x\�k\��|Q�>}�Pp�f<rF���.BQP�J�\��d���Ka�]-J% ��T��2يk@�\�,2��Q�_������A1��g��D)�*�yC��/�	i�wV�$��4g��p���ݟր뉶 �𧦕ձ�U;!HR�]L	Y���}m������3-�����wO<��n�i��jW՚����}�
���$kDQ��^�J�<J����K[ƣ��z�u2!�w�q*f��߇��KZ��Q�P�	�ড়P1� OF�L�u�NL�}�����Ʋ�5��Q*�~�dz^�f�q�{F�<�3�[����B ��r�C#r5�o�^	�g����!�dx��-��PL݅�>}4�x z|��M~�X�$Z��� D���b3xHZ<^���ŜߝX�LvP0�ۢ�у����|��v�s] >-�P�Nk�5g�­kK�����~�#}X��q�ͮ��>��[�%g3�4=������{���5Ԙ.���
��������Z�:�,�O@��q�'��ح�y��I�:Ѓ�z�.2�l6�����I��[d�-��&� ��j��Z]1��Sy�p�ƕ�;a�[�q�ѤL������<�5��~ק�GM�8mn���_�l&��-����_H /�����L�����k�)ʘ�߫���z�SyWHT���q�C��X&q�}��uk��J��ϕ�~K�A�PL-��lWd^ý]on��8�T.��~d���1�(�(d�S�&Ɋz��c/��W�<틈aQס7� �-F��m	$�͗R��$>���Ӓz�^��K�xe��W�W9��_S��Y�`��3��|���㹖ȖD�� Gt���QV�: ���R�P���=��:��)
}�<����ѡ�o�_k'&&lJ����i<k=�n%�D�6��l�Y5����+���s�BA2:��z��W���Y���*.�utC_f�?��
�~�)��P%�K���pV����=��"'�EVw�x�v��}j� �Gvy�t�o[c���,���Tn�⢀&U��Z]Q�rސBV��W�,���)ˀ!�c��2���01��'�($�I^�����R)A��@*\َ{CE����7 �+�{�7ܕ�(+~>�jG�υ�'<Xum�f+PE�-���^�΄쟸A�p��3Q/��}�������S^��Ρ���ה��k�Z��0�Ïo�Ү��s
_�����*B��Z�4���3�,.Љ�,��%��o���������sI�̔Bg�*̤��yڷ��U��� >�*Z\a\3k�?����V硿�oE�������M8���K�^��#�¥�]��v�`�:���m��Ya��휣�b�R^�i]wD���Y(-1��h"d�{m����5k�U�������Hw"'��7�`<��z������D�O������~>.����#�ﴞ�_�'�����!���F`۬�]1*�)(WIY-+B��2�rL/� ��c>�N�`��&��e\b!	�����ߥ�6�(�l\�v�tq��/���5���xe�*j��)�����p�^���Hs@L-ߐd��C�����
k�'m��]�[Y�^0VO�e@ *]~ ��5���"�	���)��j���Z-Pve$r��"c��Q��v����ޑg���)c~���p��|z�H��Y>|V�K>>nG�v�t�P��Q�T^�2�۶����
�1�/T C���f,��b�� Ib�Cq�Q�7��^�,�K��Z����if� 竳�FqX��S�*Z�,����c����҆<xSO�p>,grz���w?(܀H�
e�����[��|�["${����!r�Άƀv�be�W �-���������3gu$��/�j1`u��q��?����bE2�P� �f���Id��B):��N ����+�}�
k�6��f����v5>�靁H��@˫�9�P	���(�XB�Z!���[�jXJ<�]��`�Ѡ)�v���l,F��I�)��| ��@W�1j>c~���ys'��i��'�M6�9����?!0�C$�8E���D�(��a]X ;p���"�3�__m��`��3.]zO��£iJ#�^�C����΋��=�[���AyX��?+Zě��74��*���4�:�[G%�s�y���M��|��(�m�j�� aԞ=�4�0���r;�3��<��X�`TZ������L��m��@�{5Z^���Rؗ)�ԏ�l�ދgO�O�t��lE�y=��U2;y)�4���^5.^�%��,�G'&� �ٯ�Y8�s���/{�E(lp, �������F�뽇{
ʱ�s�㹅{�+�S�ˆ$��B(0����]�����|wr��,��~�v�=�'A���y�,���}����0�n�|�u��+�D�u���çQ*g!�Af?"}���)E8!$�W#����e;�T<ic���>�O+�N�uEX��F@��\�Z�E�4�ߌp���!��ЏӦ����9AO����(����8����/ �&������Kjg~�(�Mgo��R&�WҰ^��^m���S`�:�f�{|:ς@�-�{�.�D`�?�� �mF�������aB	z����Y1[��lG%�r�D��Z��0�@��:�[���[���M���:B��\n�7�l�N�i�}4���3�H��!��������߀�tm/�k|��Њv3䡜>/x���|U��A!f#��ku]��jas�F���������0Y�9�xZӁ���-�q_Ѫݑ��適>�ղ���l�#����O᎟d=��O=����i����y��B�>�ĪO��?�������<Uσ;�T	ݻ�+fg����mL4�@4��I���L� �3�d���
���2�#g���?a�Ⱦ_e�9���V�54��Q;yG��/j"�H�ajg+�՗�@�C�k�V�nuZ�f���_0����f7��4S�E��$�1q��e,��#�1�r�n�S]VV������I��`��O�Eu�:j�%�F.<�C}x�Զ���	s�r�5�oA����Q\�%��6Bh���wA-��l��� �8!�g$	�&��d�����X+�+����>S�xd@���\E~�Q������̡�#9R��}��������}�F?�NϞ	_�6�|EtȻG����[*fȸ�Z��J�l�+1�:-	��u��0�gB�hFT�@���kh��1{��Ay�7�(�'��Jz�������ձvLL�`�xTr�#}��|oMħ�zy�3Hu�O[�@SH=n��rq�E��m���Z^�2L�O��i8���zm��~M��Ѧk�D�/\��"���ˊ�A\��'��:��P�l
s�� '�^�n@�\9�>y�=p�+c�����r�cͼ���>b�Cp�mA�?���W��B"�J���>�5�p	����ȿR||��_��5�]�Fs��hÉ���A�!�RY�l����N���7	Mm2.������|��0K^��Ð`>�1.� �.�~�a�Zi�-��2���x{mJn�*�束�O��H_l� ���'A���E�v0���3W@�נ�׃!<t.�垺{b��ub.�W����ne��&�A��K	�9ϐi�$_U�C��c�� |2�\���Q�H�0�g�ΚC�J i5�DW���#�q�xᳲ�� ���zv=>Nh��c��ߕ�����j�4?�������-i-�I����d.�����Tc�dVa�w1~�=�9�:8��1=vM�l���(��x��1kroHA��p�#��mt��F�g���U�w	Ew�Yn�U�!����>j'h��r='롸N��mvlI�����k���:���Qu�å����d���{޶I����s��'�����S{����F?瞅���S�(=�bTV��.]A=I��n����YzV����|���2n�:�ѼQ�Y�&�#{UR*H�S�q������U<���-��@��-{ݬ"���v>y��fX(np��<���W�N�ko�CWK+-�E7F�H�ӂP�����+�[X1Ÿ��kd%�����SΨ��d�#WO~(��EΝ�?Z�oٌp�t�T#8�`3{�0�J�����d`Hq![=�<��r�!�+��W]�)eS-��;z�<��,TҼ,~���Ktg ��ڳ�o�+��J�Y]]��`�v?��*@��pU����ޟ�S�����4h$�Q�J%
E�ШdHi3��%)�$TN���쎐�:Bbۆb2O��Y�Y�:�߿���^�w��~����p߯�u��{����%��K�o��}ς���PͅKKP߇�b�XC�Jh,�J��a'M�S)��k7���J:�|�f&�O[��h����
�Do`E�%�Ⱥr"���y�u�ڮ�i�L���řV\K��H�E�dIC��4�1ִrW�Ps����9aM����{%�Y�]D��ޕMu�jY�[q�Խ ��]�;�m)�F��!�/�
��j#q#ٺ���Q��y�vXta��)���f]&#���É`�8�M__!�.ӌlxB�'o���\�ՖEtdІ5��N��ʝ�'���=�],v�tw���Hl�K*��t�ZD9���t�0�#(ԓ���ͦ�1��H�:� T��t���:���,OgJ�h�#�1��V%ئ�
�]+H!3/�������Gtb�:$t����ŘH�6���gf�4A��٦s�m`���R��:Y�]�ҧ_9gpVk���\-q�?�81����������#���w�%�C8�FS�PA�2Q�ѓ����R�k����&Ժ�LS�B����v��#؃͋�A$���1Ã�:��9_��^�g��k��<?_��I�Θ9x i�.�Y���+�9@g��Ϡ�x�(��3��$�&�v$>y@�I�!�e�fG�ڮV�%��IlN����W��O�C�Ğ'���?`h�Ǔ��z}+v�=�]��i��Zsf����[E�_�����b����3��
�Z�x�X�y��a�-Oi��jc�f�}m�tU�0�2���)��T�X�`1�v�s@Q�(:���XD|��@g/��y�j��"ZF0����/��C����G%��_�?dr~�$v�r1ֺ�a����&@�����`YR��ŏ��%��ʣ�=�6 2 zBm-NΆa#���H�e��,B]���W�g���I
'���.��'�b�Dg�k��e�/(*���ق�����8�Qq�V��ںM��)�,η����\v�����ӳS�.�������'d�X��+DP?ڸ<�jw^�,��S�>�A��c���i4�%�y�F��#��3a��	8�)lSU`m�3.(�,S1X�4���U[}���.�7y�>�̾�_���5��:��j���4dp ���Do5�[d�2F�c�"1�Vq�j�cdb�ٸ��
J�E¿�z���3�׍�3�z�1i0��]p�U2��q��H~S�B�B�w�G�"�
��*�{�?f��h#�������	���m8t
������M��0,xj^�<�e�#Rǯ��R*�qV��4B���]�[��l�:x�ʻ�Y�Q��y{�L�2�}��X�u�v�	���}'P�������@I=ϿɈL���O���Y
�(�<����M��C[�T�z�Lߊ���`��H�����DL�#�FFze�H�
�2���@Q�7���B�Io��!J�X��b��Iڴ��ӹ�Q/iS>Q�_�0��=Bh��i(�Pi��T+��#�i��~~~��*_����cۨ�w� �)9?�G��e(O���Rw�&:���=!���=qd<,�zx�2e�xł�2'O(�^�!׊��Ǔ楞��:� V������j���E��O�Ǒ��H��]�&�T���V������)���X�Q9J��-���ߝ���h'E��Wgo�J%� Ü�����y����%����8#�$��viT����y+!����rG��VA��I�E$��n��n�.�S;�&����Y*�x������ۙ��'���kb']��-t�J�
��~�%���7�˝�;��o4���Ź2՟�W��ؗ�L�����XG�|Mw�^w6oq(wP�K����(h�/_vOs������f����ʇOt<�y��l��t���ӵ�S�/+2ӧp��7+�/w1�z�/lMc�����}Ip���'� Ǫ�wH�5���>J|�蓶���5�Yo��㐡��t3�\��ʽRMK.�ǂ	e�m^�_}�7!�Us!Π�o�ܹ�f�f�P�:�f!����cT=P>��u([C:e����o:�2��;`U,�υ�+�^�ki�2��2���A���]�m�Apr;��>gǊ��+���ΰa؆��7������m�uO��������_HP��c��>�v��R`�o��l�C�����cLdz3Ф6r�8՝��-|.)����KX!ո0]����E�7N��-��=ޝ���P-�Kq�<����;+,�$b����ҁ�錓HE+ksH�������w��fd��$��˕'�?�ܫC�|S,���CNx�y���N�Ng)9��K�Kc���o�瀧���.�?�3լ��'��u����+����JNE�#A�x?##C����=�(�ؗ���w�~S��E�t�K}}=i.�?����c��1�� �GCV�e���_�������@��=E�(�m��/��h
�.�R�JZ6�	9̆�iCgg�OۂC+�B|}ۖ3����V�����X���1t�be�h���R���	%�ju��� ^t����`���ӵ^������9�.�Q����Yfn�&j�݇T��j�H{V���TL,�Q-M=�!s5�C-�����ɔ��<B�c�I�)�g'g$��1���o���k��	J]��<�l(9���C����6\���	�-l�z���>^��9�ӊM�/��%�=��lxD:����ṛ���կ,W�k�P�]�~���ٽ�=n�ߪ8��j���˛�w���\!U���Ef���2̚v�yυV1�[f�drQ����yv��u���̯��?w%�)��+�;����]���]���j�ΣL��Xyl���������i��xC0�\�]�]��&(��F>���x;0����qΏ��狘Umtx��`|�����Vg�@�B��y�)��ܼ�,�L���W�hP�Ӓ�?����s�Sا�� Ã���\�˝oFz�)(W�ǐ�-%�ۮ.'�}ؒ��_lE�$��=��|Y��*��oM�o/�`��+M��\'�'�w�W�@>�qt����ѽ�Qظ]N��a�=[�6���xԼ���>����P�X�0�5曆����v�w%1ӵ�{|�m�h+��o5!�_K��P)Ͱ�9��9�n� ���WY���pִ������YC���R���%ў����o6gM�L!����T�Pp[�����o������k�G#� l��:�j����n'�C����2���� �ڌ������8'f�L�Ȝ�f�r������{<F�r}�L��7�4���x�����9!��� #���BE(�ր�����辅��~ju@�%`�j�풙d|m���d�lS>���#s�m�fΥo���M93\�'ݍ���n�Si�֮/�%�&џ����Hִ����!oB�y���Q�zJxq5DvcP۴C��9ūq��7�t�>J�_����(����8H�ڸ�S�>y��H���������t�b��bF5Ѷf�R{�4v�_�K+��P|$Z�m�;ў>�f�]_8����X�f�1�IK�y2��}�>��*]�«��-�	W��:-`�M�Hv��F!��HS�&b�8%&Q�̪��[�pS�v�o6�l�\��ʜ�v����N�������C���BA��Y��#v��SY��⼇>�}pZqY�Q8�8��j��BKc)S�A��@��^�����]0�O��s��;���]�QNv�ei��)ĈY��ZϚan�꧓|�.՗�J�:wLĲ��	ɢ�?�q
z�"�[0��]��1g¢r�k�/0P ���4�fF��M���I:��WGQ�Yf�{ �mC�𯴡&A�CXE����GCv�.,&R4�<�1e�tљ��e�2������u>FN�	��WG/�a��򇶢����>^�>��y����`M�TmqP̊�n�W�q������?�1��;��v�	,L�~d�.sJ��(E ����5u�EQ�fY���i��:�`}\��T4C�c#���v��w����Œ�J�p�!(�q�c���Y!����Lm��e� "��$I$UXm�d���&$�@	�K�����c�<j��W�>��̌%�5�J��	 ���ӟ"e7��ƒ�;qХ4YԱ�㥯�P�@ˊ��)&�ksϱA�A�r�K��"�������@b��>F �O�����~3�)��9�`���ǗL�9��y�{�A2ω����~> ���k��m�
ʘ �m���BL��;�.šXsoddĂ@w �b����?�:=�ZeV|{�)���]K[.!��_���"܉}S	�B��`��*�G�X6�h%�����G(dv�y��N����9���u2�ξ)���=�6'�_P�	B39�׆��1����<�R����g���'�pS�
�;S^���[�+w���K'm}7��"&l�Ӽ��A�R�N� �v�X;u�l��֧(�#{�^,��5;�Q4��l�-$��x�sw��������]�>^�y����,��$�(O��9�ƿ��=F�K��Y%Sf�C3������$��e�{�W{8��im�}�p	���V/|�KK�ɓi��]qj�L�5���.#�5���|$%&s�=��C�1� ����Z~%�2O��+��$c�Z��i����s;�*�,�	B��rR[������KBii6۸4��8��)It[�(�4�F�;��&�5b�kh#M�3��(���wn�>lZW��?:D,X`�"�H#z:�|\���{S5�Ub����b;�����\]I5͝�װqF;e
�8Zg���X_�@��6;��HEWC�<2�(:������~�ߙ�KO�����yyy��"47�$���������0��[��[��Ry�h���F��
E��;�f�>����@�x�2���S�^�XJ '��`!�d�Sʚ�� ��ϋ6<��uo��)��J����u����6�K�o��-��%�����K>�$��}.�����o��-��%�߿d]Χ��d��8�k�,شtQ�k	�w��'?�9���NP����l��b��/�G���8�E�b��դO]���YS����I3�a������N��l��_��=w�=����_�����Ԅ��<�x�΢G�9�X�x���xYeŻ�p���lʷ��Lr�W���'��+�cC3Uߥu3� ��X��%⋞k�r0m���F����+�
�/o�Qx���H����=�0����Ig��I��Օ(D���u�'����3̓��ȋ�&o��}7uss�����L�n�1���ϒxmК�N�:l��������L�M��͇$Ѓm��.%��1~�;��Ï�S�u/�X9�<��kj'���5�r-�G�q�o�+**X��sx'N\O�u���fr�����|�����!�x���߾~}��X;���e����	�h�Փ��O<w�ɝ���>������!��XK���&�`����yy'���S�=_
�ք�������'��3�6�T�VR���/�?WH}nP���G�w�
�M�7|`ZC���hu����)\+#q��;�sVV[�f�]mt�'�����c��]�����KľL�q����޾w���n5��8�u���())��}l���>�����<��%�t&O���Ŗ��$��Dٽ+��s�c
��z۸F�]+�g	�0�����ݓ5�L�z2w��Sh�ME�*�՗s'����Z���m>��K�~���4U%��d�](E'�<����Ν����Y@��e�zI�K&����`�/x��X%��ܖxhZ�&/#����G���@�}_G�����/gg�E��1�8�v聘�ĜOn�x5U��[kIݲسg���7K���{�ʪ�P�j �h���ۄx��U�yRNJ��|֫�3rK˼���HI��K��+6OP
*��W���}IYY�>�٢;M�:�}�$��1�U��F@�͍����1#���l{�
�]���RZ �=�j�٪��u��a�����x����.��'$$�$���i3�6��"�����ay�w�=�<�#��t��|����P��P��5�p���YƑ/⍿��P�T��L"W��^�H�h��}�����¢d�]�=��t�Ѹr��"u-��K�
���N�
�	�]�FX����z�t:f�0�3yx�Ҽ��ɵ�����������W
��S2k\�򭶬�Mc�QV��t�o�uN�Hԇ�"��5	��ș qCR�����Ż�Yj�l�c֬Ys+�Ħ��� �`9�$�G^�g�2�Y�y}ʑ�	,� Iu8��j�+ٙ�����;�(��}��á�D���,z�֚彽�1�!����ew�0?|�p���=d��5�j�[Z���;1P�rQQ����_��"�R��h>�'�ؓ����g��QZVV������� Y�,�Nۯ��C�����E��x4�^�xx�9Ȅ�܉����x����v)H�7 O���d_y A�	5gq]��V�%T�-n�U v8�i��ݻw
�`�����H?	���e�4������ڊ�F�U�gj;;;���y������,�r�'D�ꙃ	N*�$I�l�䜳�@���TwVXX��E�~g �/�P�=f���C�s��ȓ�ʩ������ɰ��k��ҹ�o5����K��8�@���Y��\>����v�)l.�6ـ� ��l$"a�H�����>8!^�q�"�2���ֹ����꠨�"��و0���6�����[�D��kп�������UZ0e�jEp��Pҫ�4�*�77���;�(�����_o������&3D ���_�x�K��no�N����>H�J���)������V[FH:u�C����g�G^nt�����_�ǲ@Ą(��9�HBy���c�Zw�\i���颦I�y�!)���l�o�o)�eOw O��׸�e�p]�V�U'F�}����`u�h��j#h�8aE��\��I��
9A����~�@4�u��ȠT�AX<�a�?}}}e���5i(�ӭD
�Ҋ�XND��F��g�\q�;��?u�#Ȟ_ӧT�^��F�D�/O,vPШIZ�0$��XG:B��s���ψ���G�������\�Ȭ���Z�S8Jڎ�6
OĔ��p�3���3簦�8�����`_�l�$�����K=��K��Y����zezhl��� ^DP糳�S��?��z|>��
�����+㇓kX��<�Y@���T��c�����	3�F�ӹ�\�����dw?͇��SrEݜ�?)������X��X�|#��8 .H��.z���ϟ>�vR�%t�p�51�c�%�������s0���'���NЯ���Ќ	�Z����_�F[
O�6�a����0o����(i@n��H��Z�o	z9-6+s�/4S�U���l&(9���!�-_JN<���%H�6��
��Z��Ʒ�ՈWx08��Z�=�����	�����ju0����~��[|IFٖ��������|�>b����?%�>e	.�qV���>��V��Rɾ��Pv��̿�P�$� ��{&P<�d2&R��ƙ�!�(h�M7>"�=l��F�;�NG�1�"#�4+O������=_A��Z��KI��F��0z�\r)��V�t�^<ovtt|x�j��ϗ�9c/�:�Iݸ0�&-H\��SI<����j��ӳ�=]]\��IjD߲�]_�(��-�l�PeY�_����3�a-Mf��|(`��� ��<�{b��5
�q�[�)�9���<��]X$��HpǕ��ֺy�~!sI@A���_�&h_bz>D"C\C�za�����P�BfZF��cFF�6�#��8~i%?��}~����BHpH\k���˗焊'B "<�㡥�l2����u=z.��W����B0"W^k�����߲�ju=BGuʈ�|�߬A< �?P<�3���2]P�z+[�����U�m;���o�&:V�	e]�_[	�J���u�\,�E[ֳ2��4S�ѭ�����͑���D�e�SI^y�
Ƒ�e>h%��ڬ�0J�c�Z�٫x���0�[Éߕ�:q8�7��
�: ����ε3@?6-�hu��"�����X��y�p|����=�`��f�sX _�G���sQܐ�3ӎ\��O���5�m�v�@1�����7h��a'lE��`����Y4=h�C���	�$��P���Ȁ�%LTM"{��v�#��R��i�lBO���S���nd����c��pҘ�U��ЎL�M%g�h���� Z��v s~�\ �K�Q�O@ �m����J��@�/�<�qߴ�w�\n�Q�AS���|�o� �@����3}�RG@蜟�t �PCÉR%�A���N��p��Zm����D~P��x��6�0�X����$L����P߉��kyAb��SS����$$?w���E��-m�D ����ƴ8�Լ6�p/mQ9�b;��S� ­�ʪ�<��%��,eS�<���+��\4�301�<���f�!F�Ӏ��|��K;ہ��������G�Y�ś+a̡���'��$�SVvp8�l�� ��fNc?+##Î�7tP�1�pI�M����8��|X�q7��p�f8s��������1ϒ��o ��^^^Q � (ـ�,(���\%��m8z{��K�){{{;gg����b�yN�x��#vt,��U�|�! �K'�}�&�P'Z�PE1p�t*����u-GLjz����ȴz�'���T~��~���Qd ���|T��\N�-�̾Π%>�.k�d���5B�p%�A�b���<Fm�LiZ���\���5'�[�Ò�eAAA{F}x�S��C2�(-�$K�s����x��1	�7������gTy��
�4��F|��Y#��8`�����	�Y �g���sEX�j ����X��USR�K��Z�3��@q�z}P?ꛠ
e����e��_5�����j���L>�&�/P���[s�.�1捞6�w����ETDd"b��H�p[#
��䱱����p[,�@heq��+9g�8�UI�;Q��`pĆ�y���hsf����nNN���C�M��p�7>^�� �Ċ[Ʈ +;���L`Ts��MM�
�\�)��>yG�T�t�)�g�p��_��^K�t޸��y�>�tC�'x���֞#)%�IƝ����?Y9d����@��m��x�u8��V���Y��f6���ڞ�\"XsJ����%XM�f�!BΌ����?`l�Wu���(k5Z���'p�ף�f�&��!dw��[WX�BLG>�_r3���-?:D��!=�PE�e��w��������=���}۷����"�1�_~ �DSq&Y���:VHܴ�8��&t�F�y��g�-~d�%>��ضe��%��P�YXX����1=��?z
�)` ����BjY�tYY���hޣ�,�f�'�I,C� EFH�tΨ]FR�,/�b�D����͓��������3O�bWW/�
N}I�Kh�@q^b�&b)S������\mVP���Q��C���R��,/����]ڰ�����d��k��Czu��@PN2��8<KQ{�k:�O���0gB����|*\�/9��28��1n��MT�G�L�^� QU:�WUH�d@M>m���"͎���/��ֲ�xВ�ɏ8�GQd��gl�l�M���6O�t$7(B$)�?�VX<��_�I*q�'O�o.	+��&�Eo���q���#VA]Э{� 1=*��7���tz[��W-/y�% 吺H��#\�'Z=�<}]�f/R�)ݍᤴ]�.�1MnO%�8�+���9V�a}Z.6�k�__�H8��gh��Юh�#�:(�Qp�[�,��V�At[ �������}�
Tx%���豦��ka ���"V�5�^�SO0�J���9IV(��r���Ff;�<��K6:�&ЋU_�F���t>J
 wW��w�R��y3Pdځ�h5R�ǝqrrzO�l�4b�jM��.��[g�*"�"E�T�֊@��X�j9�N�q��2��Zq�j�	!wb
�c� m������<��K���p[&��j�� �yJ�r_���	����a�c\�P���#w�(#��8!iZ-��8���G���5>�Yپ_t��ĸ��xv�����Pe���Z��ə2�Q&�����[�?����{x�}�4�b��A+��C=h�C��`w(½���c�PW�����eQ���i��k�3�S�1���SS?Q�v�0!��oUD�2��yyy�'��o aXS��܃�e���4���Y�A�o�6���6���Ci'���;�##�j&�BB�c�;::��������^�)�-�ide�_ī�q�����6@��$K (�Q9߿U%eDEE����S'���M����42[���@���W.�����>2`ooo8�D��Z�/Xs�eJu~G�q]'䖖��s���x^~~~&��<����VWWǐ���(��	�[W�e���ͳ��/����8J=ej�/�A Pt%U����a��x�����J��$:��vǓ4�+��(a���S�œy�'z�	&9��� `�#ěڈg�!�Y���8	�!!!7�S@3��pg��	��ё`"@�&�~y��w��PHyrJ6���r��ǜ��B�ĨD�)){(<�6L��R����M-�Pϲ:�:,���b��U/�rw����ꉊ��Kӣ��'�j�~%"<(Z@:#�<L�.��#e�l�"n���h�9��[`,�Yl�ᘱ+C�w�v��c�qU�ZS/�a�I�s�.��?�k�iϞ��h��p�S��p�r�3��3��3><��F7Q���y�����.���!ƭ��_� �>�$w(C�B:�viA��Lv��rd)��������B��&����Ԡ�FQ���Tdd$���@�����X,���*a(�R$_���ܰ*y��4t��	����H>�r�Jf���mkKX^LLL���F��Jj��� ����	a�e8q�L�np�]g�?��`��.�o�}||0�1S�Sj=�t��8*! 	͉ll8�p]��L���|�O�ƃ�\��"������)D�IS�V��Q�>�ycw*΢���l+
��޽k���1#��J&Ҥd�1�'Nl��	B=����b�<�?�`u26>�Y�m�܅�x�:���<�	>�|�\龸p�_.��}vt��_�����/�Y�����}i���+^|8�W���T��{�$2<<gC��8�t�НOt�@�V8d�>�����[�Ŕ��^���?��p�9U
�[ww�a<���ד�Iii��N�H�w�*+QJQ��fy�'T&����f�l��f�A�6KrÆ���ʄh�Ș]L���29���"��f[AE��왭H�����$�u�)�2 6�>��{	6���%ǌ���-��(,$)�P3���144D�*�P��l�'�рqU���fnnNOy�2]K�!(����^�����e�C���'FRa%͖�2��Z��g��@{a`��šq��]���ߠ.Ȓ�T�݋'��ت�����o��}J�N�X�c`$�ܥ���
tk�H@������X�q��o$ZgS7���[F}P�Ћ�n�@�l����
�4�y:�]I	�ܓ���ʪ�	dޥ=�!�yU��u6��POS�hUU��E�%��~w�����v��b��u��l�0)��������Ap�^j[�/x^��<�Adt�X����y�v�eFHH�+����i�e�}� �Y�ٍ���;���*����("� � �
<���@!�.E8ST
g(����h����^YY��`0DvGiwrJ��|<*�s�ܘ���`��*咖���Rge�m���xg-�e=?�^*VR�p-c��ى�X��,���A	��0���̰���qn7J�S(�~Qeq�H ��@L�0����[�B��kEd��������* �����MފA���a8���;
�vy�`�VBBB�Zu�����zks�y
b��
��;)�q]�T���ɭ��t4�P���0�ɭK�:
[��$G���rѓ�[����B
=���(_���s�b��R���&3�(r_��h�A��o�⢿����Le
P&���5VVVw�\�}�H�c~/��u(�|VXX�	�&���@ſr�d��&M�UW#�@���"(	}���5���Ζ�~�/���dan���[�&��$�Y�%���=��f�T{��u}�� �Q�SX�S3NWRp����2Ț��3���G�[�D=i��z����75���T��F ��:��w���85㢂n��g�_h�ۏ��m�4��#��F�u�>J�&�x6d� �-���QY��Y����?��/?�`��|�-�"�iuP\�elMA@#��y�������&���/�ߓ��E�=��<��]���j&�ZB�GB���p^OO�~DO �/%%%ɓs�0;/���M e{SX�cF/b����ւ��B�Y*"**�Is�ޔй)����ၫ�s���6T�3~b�� n��_�G��N],Ėc�9��!іd�V@���>}�l�2u-��S�+���져�|�L!�����)�r�{zJe�x�;�7�<�Ig.�^Sb��␄8���F��q���h�ԭ������k�95� �S�11��Ȃ�@�k����LϿ��z�-]��MK���/�!$��������FAK�A-9eC���N��s�\��x�[j�s��A��{�6�� KB(N�SI̤�^p�'�?DS{{;V/�H*"�@�JC6u�?�6*I�9.��]Z��<kj�2j���͛'�a���F����,��o:f�p���\�
J���&M�uc}�<���R�-)i�8H��AW�A:�:�����Ɍt�*(ෞ����~|�J >:��6��ņ�ed���܉Ȋ�+yu��*C-�/C��?L�j͔��{	����r�^ ��k(7�4��$V=�	�U��ng��x�@qܤc�;���_�*�jkU��*jĐ������&L!�� )]��$+�E�?������p>�_]�p�����d���hˏ�]��㸮`��"u�����It��
���i��y8���f{�={���7$)���� 1Rx;B�6T[E�?Խ����STYY��8��i���kvv��^8��n��0X1��[�註�ɓ��H�ߒ6i.jř|6��5G�ʳ7/�OB��)�vv��ĩ���Y6�Kq������kɝ���p{944�:>>��q
�,Ζ4}�=cF��l���c��2Nx�������)������c%h���J�tj:Xt���^�s���� �3���>cFRYC��EM�hsNk~o=�M��RK�����"꨻:q�Zhd�_D�$vU�vu��
�-����dƜ�9��ܩ`c|g�P����:ܱ�����v݌2��@�(�;�R�[���}E;e���BB�ׯ�lE�!P���H2t���+�f�+��4*��胢�r�AH��������
s\��#,2kٲe-Ǖ����d�C��-	�v��t�רm���(	Md:T���čj����:w��T"��>n�JK-na�T��fM<�X��%,�V� ����iOi!�ˍ
�0����-B	d\�3��LF����1��G�\��eu`%����B�����.�P�M��8KV	]L�t�vnAa~����F��� �(��ʧn#䍠�,�~(R�=���fc��������"&�e��*��䯽T:�|l�+�*}98�h,z��Fc�*��E�;J~$N���[ϑ�-���f$u+,2�c�Us�m������P�Z~&y;�H������>��d	��ɘ��I�,C�QUPQ1DwlS�.S�����W[m��t�����I�f���Ѝ�j4fs�����86�v��딅E���F��`Km>|�ø�ĸ�A��u����d��Ý��;���b H���%]I�~`�)��,newi�Һ�e���~.Vl�NQG��� �R���n�����a'���DP���PE���� �&漁�???�-^T(>�#�uQ����;af�9�F����J��0&�:�!`~](�Ѹ;�Z,�e�>��m4�Z�`@:,3ĉ�j����P���� ���
��0Fe�??�I��j�o�����.��r��-,?����i���Q�n���|��.
rT���u�0�y����$h��ʔ�]��X����`��S�U��pm�S�P�� �hHS� �(�ni>���ゃa!���mSb���8�oKS���V��h�|��g�I-��dS�YJ-�������|F�����W����}q�f��uA`�S �A�������=�+9�2��`���F�F�����}H���H�ڈ���[Z>N���\��X!tQ3����ͱ��/씱
g\�-?�]RR�0�9�f�P���n� /��o�@9�~jRC-���0��F�E��F��<�e)Yp}��3NǺ�x�������f�jx��m��F���N��l֨����@{
JJn�p2�>�AB���#���b\�a���Z�b�Y���N�]�J��j�Lvs�]���W8��')��;-�s�]�~������ҌWb3��7t��y�A���r).��Z�mgt���$@�CЏ��{�pRL���!(555�������
�E��'�_��t���(�ۻwo����_H`��dd���h�q�f4���`��2gv��r`n?�Nof�s�љ�ϫ@G �W��N}�1ണ�cjr2�G\�ǣ��3���J����c�ݨ����JR�JY�7"ԸC?�ΏE)�9.�����\�����G�������e,5G���~*�M��CU� �
_gq^��E:)���w�Jbu�bG������ Nd�}�*��P.��>�4x�d"/��.�A1��F�V����W2~*#�E�E'G}H��<h�f�����d�k���erB��w�z�3e����e�{����}������p3�L���XRJ�WWYT�4w��|/�.����c�GL8t��h';� f//���˾rT���<qpwA�7r�����g��,��۱�����H�rRr��\=��0�1?�@L�����o�g5G����o�z��n͓��P ��W�but�Y9KT"K[<������S��#��������v�������>P,�� �78������s4�eTʍ�_m���,�_9G6t_΃���#��s �wU'z;2Rt��Hڛ��%$��֔3q�3���k��mB�}�l$B����K$���&��� �nnn�x��n�OhM���p�g��+W��%W�b�{r*G�#��S1{���[��w�U�┉���Q�эS�d���	0����?����P���H���G���P�&'�����Y46�?���,���.f��S1�@�����IM�y2T��b���@Y06�}R��ɓm1B��q9F���#�;�er�9�a����w˪݇CӘ
��C��1�l�N<;-�i��U��%���`����^^#sdM� �B Ta�s�����IU߂���<5o55I	�s���/��֠�F|�\��G��w�Śs(u���1%�I�'�F����	�(ऱ���`�J��P�Yvu�;|���	C+u͕5%߾Y��~i�@�!��# �L'�i��=������G��3Ô�jao�U>���S{���s.u��Mʺ�~�3Ф#��
���ohhPp�)-8�8���b���MT���ԥ����@������(��kMv��;枃��� ����a�Z��5�2�Y�zU��޼�Vi��P�37�[#e����9���L[�#�d�ɐ��S�ټ;���Y�c�����n2�"�� |�N����":RJ��p�Z�����_<{�i6k��ʷMv�R��8�8i b瞢Yk�x��
�b������Lf�=����,�_�?� d��k30�t����DmIKo��ĕ@#)����minc�㋠��N��P[H"�')Jk���L�	�bpP嫑p��1�oі�ѭ��wO��ߌ	C����������u�WJ؎���+u偑��Ē,vN�6\o��N5">����T������w6g�D~��Uw�טn�-���l��$Q�BX����.��(��luhv͊�oy
���Lg[a"�@�
�F�eg]�=�������1SH�Dtrtt�̃!�٪�*����-��E�����g6�N����\Y�#�g�:�!�RF����!�lLLLSY����m�;��"/o�u����������6������!PM�����H��<wvvVXF�kn�N�e��#����iH#���
Q���Q�ub2�:�
���3gC��a琒���ɭ��c���n���Q��bo`��m6��7�5Y�2,�N�
*H<��ġ[[��	O5l%6F+��}��U�N\�5�9K
����,��A�Ȯo
5D��x��0����k[�3�5@�q��\A�T���c�;P\}oP8 şξ�2#4%���(b�&�d�^'�P��i�L��
m?ť����-a%�iFH�?�� ��[�1�K��y����<�*,4t�G��N3��X]]]�@�Z�qR\������O�*_��n�ƞ���]��3��
]���ݨ�1�RI]��d��?}�*-)y�␻!0��3�N�U2�c#����Z�s	&9!׮]���	�C����s��ul�*���ɬ*�-��8����u˚��ZXvǾ:(�s����<1q��O��.gZZ�e���7�(~T~�qwԇ�sO�n���p<�>���(���q:�^c���ju�|n�FP�J��/���f<o*J�˶J����8:9�*|��BI�k�-1�p��0�Z�U��"Q#U�wGݠ�Z�ӈ~�m|x��*mL~�LG\��d���01.H��O�F�s[���~��VosW����i��|(���)�^�`��]�I�|x�]���szhx8����vŤ,�|w	mN�P����#p1�ݎ⪟v;�9νh�>|(���S�f�.q���zFF�>��F��H�&�r��O0S�� ���?}Z����۶m�ɰ����Ay�����f+�b��I��t�d)5:�� j���HQ��7� P0r�j��ǳ1Ϗb�׽*?�l��+d=ř2QlNA�:C����IV���qɞ?����)�?G_*�2]��<)�>�T��"�����U8[Ҽr��&�~S�a�w���u*pa�sNYD)���@�N�8�`啼�]��;g�-���^o�o��J rA|��K=P(0�U[���K�ۊ8�(S���'~�8%7\n�}��Y���R�0cU�ћ ǀq���ޭ�o�b=P[Gg�)��z���iiU	(W-���
i*�)��*����肂���U4�riiitC�xdVF�9ɽ��2+>7(�ڟu�c���]:uo6��x�ړ}c��o
6ų�[l�ɼ�|�w#�O7�/N\���xl8�|��ݛ��8������2�w���B�+V�)�M_�h���d/t_�(~������/_�|���;��x�L�;IjLl#���,}���;���MsR�tx:T��cN㥆�4��!>��}9d�c��)4?CΫtp_�n�JK�v��ƪ۶�k�%�U�.l��cF�3���vySs�/������nm�B�ۍ�eѝ�sr�V�}D������P�S�c�;G�ٜ���.o��~}�a$5fJnl:��ľ�z���W��]��۷:����Aj��j�W�����"y�ګg�B��i�9(�G���;����
a|{��!����o�������w�÷���u&����Zf9l��K��:7Z����[k��>�\ڄ1݅��ͷ��ހ�_�y'�}r�s����d��&2��@e�M��99���~5��ֽ}>6��oP��.5�	#��
���>�,�qv��<� ��3�U4��_fd��{[K�q]%�l`|��q��xX2��PoKR��,d�s&FF�I�S��m�@����aٹ��*����v��7�p�4'�=�|*b��cVR���Z���c�߾=	�9�A�@Z�,
�55߽{���uF	��ú_�\{������\{h����Ȉ���䋠ht�)�u�_3z=sTSr�����8���KS�g�svK����t��܀������!f��Qf ���y{_���ŋ��7\R���:�h8�|�ңŤ��<6�)<V�A�j�:e�r�	��~��e�aO�}$q�n��K��e]���#�ء�)�d�>D��D�G����IS �i��v'����a�z�PZ��QIA?�T��Ҡ%��w77�F�� 7�<������J�𲉿�a����`��d.��I&��K-�CG��d�M���N�={6fS����.�?���-If,��b������3��[-Q�$�Ӯ"l�KY�Cv�YY�J �_��j�"/��"��2�c��q	��wa���V��\��2	2L��6^���,&Iu��/������R�,N�O6b�ݦ�(���B�w���@��\l�J��f���Gƞ�.�����F1r���w�ܴx~�ڭޜc��taQQ'
��>��]㿀���@�-��O�Υ�����mD��V��o���S��c�B�̊�CSU�%%�$ �3rK��\�e����ߤ�Q3.�3jk>�60���%����}�;�ī�.DBo;�R�� �]RUq�rµ�ĩ��9��j����A�O]��'��J����0^�����2�2�+MvK@@8)�_�o�+!C�ގ�ᶸ�ޖR�HGo�-}�Tx��27���b/SRT'�rr�a�sw�Y⿛�8�4~Ǣ�oUI���ሓ����9��§�5�2�X �q�@���|FqW���(�yvuu�"{u��؛U��So��!��FJu� ��c�`��ħ�x���%/��0�܍��<x�`5�KC��杕[�Ғ�	{���������u��x�!_~�Ҏ+�4��U�sqI�k�P�$�3�CK ����}A�:��ó\?����գ*�+ �Nɬ�5�4coj{����|����8��CME����y0��A�JI���s�'�d��HI^^��#2wx�&;#A��zkC����2:R��]�I�|�ͨ��
��9}h�=aTϽ�7ⴃ��S�晑T��·1GpHt���1�m�>��[���G9��n�[e�<�� �q[�$�b%�d�޽���G���6�<H⤤8-:Y�m�Ɵ���&����q=�3J�SY�\���^���,�W
������I���
�	��\r�D���j�Ԍ��m�y��%$$�as��3:im�*�� <B2555姰=דz�������}�d�A|$0�c����~���e�ov�b��A�P8��4У~�(��2V-}���U��4�����'��*D�wp	�	 #Z�`�A��J����:�Pj����8ݠ���R�ۥ-d?�n�����nn#�E���a������p�ӄ?��}��m9UI�JJJeX(��X��ء&�ii[�Y��/8WX�ϝn9�W�\\}3��:{(zjrm�/S��ñedd��1�H���H�����TfM'Y�&f2}uu%C�[Fa$ �����N[��K�9�� '�(`6֟#�`�el���k�C$��5����dK��7��<�4@*�nR�v�^�����,�:����sa��j�-	�.��7ߎ���Ɣ�C�ݴ�K�X�!����	{��/�(�2�F�M�';7�S�&���26�7X�'��Jnnn��Ҵ̨�SD�	��訨���(�"i�Y���QE�k�=��ɺ��bbأ����(qY[[�'���d�j�vO&3�4��������b�!�8�b82DI�I�����S�֑���m�NF8�sv:+?m�u�L7z{�����0���D�$��pz�%Tj8!�)��ۓjg�υ���k�Ki))nz�D?����zl]<���M�	�XNS�R���d(�B�_��^wش��L�M�;$�����'r�{�p�ǀ���?cR�'�*��<�K%ۺ��[�(y�@���t��0��<גl����5'�����w�H�_cc#]?$-/{/[Q[[;L�)PwW 7�viW��Y��[i⵭��gT��:�A��/o�O�H�UA����	I?E������P���GZT´Q��V���(��W�Ț]F�'KSI�[�ƒ�����aJ��
�G��ނ~���9�����/�}����<���,�s�����̍���L��p��4�z����v��_�	Q��۫����_���� ;�{�s]J"��[+pwj�@\Q����x��ͷ��x��D���+o�ǿ���[.x��(�yak�1{O����(5־{`��1^���*�w`�ث��B*n��S+�w����$�OَʀΊ�I�-��������OlVB͉'w���ɚ���G/�2�����7G�#b�� ��g7�|N	(o�f#|B�x�dS5�lq�"��l���^"�ߒ}���G׭[���߭�b=y�u?� �4W(�O�nĳ�_ޯE�ree�E3�#k�M��d[��x�/�0��<`�4�^pkkkJZZ�	�BEQ��PR:�M�v�?z�A_W26𗯸�k�XK��O�>���=Y�q���(7�X���9�.�Q�NB�9E轛{"��Ӱ���\Ł>Cu;�㨑d�/��8�n)�0�U�W&Q(�F<�d�nR�$�
nfs��4����M���]]��� 4<��7��0PR+A�D�Q`�P.���Z2n�a�6^^^9����a�#����^�"����ߛs��3l����ب5ۼ�_�!���y�ga� � �~�b��4^��]%f��Ñv�n^�PD��.Ĝ���/J�����rq��c��Q�jR>I��A�+�mn	{z<�b��~d�b���X��]������ؽXzV������z�� d/�]��&�!����5�p�s�zn��U����'6�B�@�|�)h����p���+Zt���aX�nb�lsWD���-"��R���v�qb�V� ��v�?%;(���e�l��rA��Zy^ ���Cw��bܨ2	�f��f�"�~��Ͷ��)��+�I���{�����aL�Pn�O�6�s<(�Kł��kp�f�����v�oOyd[IP;��l�=۵1�M�¶u3��(	3.o=)t�#>��< �S�T�y��k���d�u&S�%�qHd/�n}������0�\�������瑧��*�e�B�.!�b��ح��?{^�5�T�����ͻb�y� }��É�Y؆��7���ěA�O�1��lq#B=��u�u����؅�3�=�Z���PUK4�]{�ڶm�7E�Q�r�XX��]x7`	e��G�5���5~+�e�
)l��^g�g"zI�Ph*�� ȟo�Z&(��p,�y���-h�孕3�psN����W4h������Ӎ.�Q�|�q#�3�>�X����"4=���<#(`D�������I��\��f<Oj�	E}�M��2	�5QUchV�-�VB�2G��ٚ5��~붉���~iI*�������`m�al�bD�-B���)w@f5Z�<�s)re�Xd�����V^�t/Gbב2�CO��7�F��6w���z^��
X8�*CU��CQ�z�A�]��>5!����铃W��F��"�~pJF�r$���ʾ�r�-Z��[v#�	��5=����
�=C��ODZᰤ��T�ķO�V��l��"�d+A_NBOV|��9�1c��{��En�=l�`j�g�A�/�rs���+�x	�^�GL��=x4Y ���/~RD[�эj�;�Q�ȝx&a�s?� ��D^�{%������� j���{L�<<bjU:��N��"{��M��������In`�cUUUx����^[[���H��ߔ�F�}$x%�{d؅˴���pD_��(�y�˯_�ЍS+� -���qy/
C�H�[��63�mnn��k�F��y�D�P_n;jR-�'��
� �ݸ;�yH�c�E#S�L�/<4��o1'��<y�2Q��C@
���M��0A��M6����F*"z|(��0X�p�r;b��8�yب�]�ty���M��
ٌz�G]H:��<>�H�&l�sIlZ�,��J��sm�q�,��7�ܪ�Y~�cj���`�{?�$���iy�,7�+~A!�0*%�e.6O��z��tLsGu��ː���Ti|���>�9}����rS�O.�l6)/����[�+ ��}�8m�]��xIA�K}��]�F�D�������(��h�'ZͫFPs|�"H>�Z�X���q�8Y>uC������C���(h�K�i�㘺��+���l?r;�>�P��$���+����;���]��������E%���]1|�}�T%�)ytd�l���/��C&t�&\.%�WM%�9׽@�ElS`���䖍>l�`��8l.$���ͩg���bc���Ԓ=Ӫ���G��`��-1(��T;:kh�M�� mT�i$�ȶ"�uu���&괪��l�x(co�d`��bȍ�Z�����|��`�?''��S�.c�4�\��1V��o�C��|�;s	e��IQY�x�����{� ��;���*��m�հ�sswI����f�C�[�9���+$�ʮ�V�ݺAA�0�q˘����,ǚt뢓߷"z}��ωcM{2z<*�ܭy����ȃ.��crjMTi���	O�v.�Gl�z��.���Z �w�WB�0�Kt���mgV�A�VF5ц���2	t<l�oA��Fnk:Wz��4[�o��F=D�͋�j.��a�=�ͥ��^W �s=��)z����!Yf�x>K:X>���D܎���P-}V��M�nz�J��eۅ����-AGQ'��Q��;g��o�v�Z ����ڸ�ǈk`�m�eQ��9�8e
w�)���^�F|�
��7s j__.�,�p�w'�����/i1D�I���̴���A(k�:��$�މ�D�Jx�sNl:���l���q�<tw��fQQ��Ρ�HT���=�sY���U�=f1���-���i�^��f���K�zNd�ǎ����62J����w���λ?$��Z[[�U��$#?����bS+H��?��3y� �d��d�qww���5�ޡ�-��2��@���#�5*Y�-~+�&ê(����phc�Ygo�>���B�Y�����5�(6١�
!@���x�Q���6��ˇ��ՉoI�u�w�ō��d�=�*v{$��B��h`� �1G���~Xo�_�˹�J��)���$�з^m6���`�]�ws�U��`�Q��\׍C���+sh��t��W���4Aa	����}�3@Y�~���zJ��4m���z<���)S��^ے}j>�Sa��YA>�s�ώ���R*��`���_�~����#��ΐcT0�"_籐����Hn�*���늖hH_Q��T��>z"�s��-S!!��QZ��4����������]B��Ԥ������3���=�-�������	b���á�
D�	�������@�Y� �5طg�Ac��f�U��x8�n�y��j%hFY�+ƞ�y8>0}kLOa3�P-��LP#S�3�8�;�*UR������)�rP���;� F�w�3���y2"�3��WG\�y3�����@y�P;ޕ��Xt�7&m�������N��"�a�}�C!��s��Bz�V��ړkQ?����1Q���OsA!�d3
_��*�&�ay+�V�@j�q�w9��E�.\�
X��/i�g�\ga~��c!�_�_�[�Ե%��������|�/E��)�[\u�1O�!k|�=�gI�����w�G�V6��555E�YQ�ZW:���qcwH���[_Ծt�v�"D���|�u6���?���N��!�"
����EW���A�}�{э	{���<R��th�� C�g`q0�6�I���&��h$~X(��7xi��}j����uttl���{f�ֲ�j�������$ԧ&��B	�I	�/�֓�>T;�a����ﴥ��jk�98?9Mi���	���{����5�}ſ<���8�m>���gyܲ(X��B�i	{Y/�!f��ϲ5G��wT�j�cE��=�n7Bf���[�94�����%,zt� �u�c����ϟ��v�X�����l�t0���誮��O�IAq��s����DeQҘ/}���h�(1�h��g���\�աR
@�:�DMd�o�@|���ؚ���3s
��\#��j`u�͏�6O~~���dSK�/w�\Ɉ^K����Yk���_�G���n�r��Pֽ��}f:#�<-�kW�(g�呁v�vH� �D���J�H��UE��u�5�M�����$ ��d4���$�c���$T�µ��k��7�t{�',��X>��Bs�A<�nY�������IJO'52C?+�C�i������v�/���t4���n%C��q�	֟K�c�褭<v��$�� ���(�݃���/.��)���zg^18ZQ��=�S#'����Z�4�s���k��$I��{Lq��8�C��z*�h_ߖ<��5�{<��]�*�؅/�sL3��,z��WJ��gc%OZ]א��&��"���\"��w�d1�PF��4�ou��	�������P �ʇx3��i�V�w-B�����.!�U#b��(������6QN�~�¹���Ѡ�V�� [�Ѿ�zw��k!�X�$��b��N�PaL��쉢��;�{Pz�r ��>��;lb�e�v	IC��~sL������OtjN���<�T�7:����浕�NCA~c�~Mь�?{�o�l�ӘAEC
�;��J�<��y�0����V��X;��_��}�2$8�`{��8q2����w���L��7��
Qhc%�]GB�is$��W>\��� ���R����ѫH��-:"<�`��%���+�m��r���C�M6��^�0ٚW��ϔI�F��Y�g%쏨�L���d��وi��5&��v_h����O�]��d|Muu:f�GҪ�א������Ʒo�y�N�"9���|�� �lR��ss`�����K=-Q���Y�:g�_woٽ�Tp�����+
�!����3b	m��:)��~fc`�`��'K���Bm{woQ��W\i�Ȋ���[��ͽ&ʥ:�����6��W�����4��;��e�ꛑ�}>%
A"/��uaL]�\Nm�*߼5����7o,���J�G�S"Y�����Ʌ1��2���z�C�E��\�iڸ�AUB�R�WP��=vS(�O�ݢ�5��� `����R��xr�����+�-g��<�&����c�h�[��Ѿ����g�
��X��p�:�+��v`D����
�S�ACeeecG�\<f�lQ��'�\���	R�{��+��oT��ن+�6�S�_W��w�/	?xv���􈶪�Y*<6�.O}�0��cA�f�R�_�M�J� ��9}�xw�������F���)��M��-@��4ukM�yd�H�w}o��p��[�����r�����w��6���,}=U��j�s;m���00������o1��
��M��aN�(�ns������Evo��^�*`����~++�����G"#�	c^$g�4|�P�^�W����V���!��n{_�c�]|8h8K&A"�T�	�1T&n����Qϊ��ʗI0%���k�RL��G��R������� �Z����nm�,w�a�3Ӌ��*�/���r�9���&�gL����&�tx�ܸ<��e�����<��2i(A�q�Q�D�衙�YײXm�sk>Vǩ�&W����q��Jl]E�o:���;~R�H�IE�Z�B`�6��J,�+���P}:όG�BcZ:�<r-̇(sY{P<DMvN�"E�R5�+��XE�����E����=ܻB?�t�U��0�p�`�h�h+w��.S�OG��ey9�뾚���<߁���~�
�!s,����(D�l"�=��Zg��=���
���G�3p��?@Ku����Rj���=_����^����L�8��k��^��i��/�Hw��(98я�G�t��
�|@�w��X@����s\�s�2/8R!QΨz��r��*	$ް�lM��ޚX����mn�c�Ѥ�O[��n��|ི���L=)p�����Z�-ᝣ7�~�:p��]��:��B����&�W}�;;]��R�Ie�xc�&�"��f*���lח�K"��[�U�C�t��{\��g�MGF�t��I��Z&�¥�|
[K�Ъ��x���K	9><���괟���P�d��y�����7*`
o��!ڷ�z̠P\�'�*�n�(�q���U*d��2���V�$��`c��3;�Wƞ���>f��z�p��n�b�E�j�O~��!��d��y�GW����}�St?-�j���u��_��̑���1�2I>����^ϓ>��*�J���]��d"���[��W�V?Z�Q>v~�Ґ��澚z��aa���>�
�:;��������Z[�k3����T;C'g��GcY�\E���1tsd�{	Ꝕe<�a��4+��e�|��-l�~�c�E����9(/�ۦYSZ��D��TE����X,�&�k,]�%>h��G��e���S�*1U5z���HcX�6P�u�v���T��]aU�q�4�,�-l���|�0��^־�7��~zW��{��ٍ.m��<�>�X>ͣ�j'k�*D���aG+�-u���&>��8�Gs���=�bt{k�4-��խ}����������B�x�c\
��9�iU�4��H�n���@]�=�N�h�5ED�����T��.�B��Nf[B�_^�kFPy��V�G������G�m������X'�Fcxa�}́�"�9�̺�Ci���(������s�Ѿ_���e,K�;�t�	�|% ��c�ij�*�cYn�n��*��\6��Y�k�UOKɤe58Ǘ����pVVV��W-"��#:21�{�v�dk�j���HgK"f�_��	��̶�����Vd��Zt���C�PA��1�|n���cc�49�\�kc!n� �i��K��b_�zf:��%D����iT���,�χ,���LB)��|J��<�pH�r\�	����8,�����x��H��Y�#!����A���g�L0ݩ;�.w�ws%b��6�����Bz<@O�H$	�c��yHp�]���hk��ЧbW�qow!��:�'r#�S�����p7�Myw4�1]ey1����j�鉪�K�i�FM#����i���=��8,i5�%�����kac�ϊ�h� ����ސ*1��_� �s�b���4M�Y��s���9�����ZK-o���P y�C��B	e{$�r����Q�'�E��l%n���8"��X�bUaв��[)�1��#亃��J8��d�P�J�S62w+������6V#��v\3r���ۅA�+R�.Yn/U���飏Wz�¸�o�%� ƹŬ�e^�]&���=��EV�
��i�j�c�$ �t�n�>�+X��ȿ� ׇ��,ӌ�	.Ó�G�0��J��!6t@�o@���A_��P�QOXE$kk�%ƒ��I�>���J.�MoszW�I!����:
d��m�v�r��$�a#6U�^L��y~q��xGEE���;��H�K{�1?{71�Cl���t�3p���T�.0_o��8&/�K?9������Ǉ��Ch�m�R�T���	���f_���lꝖ"���Ȏ�J��l�=�P$��-�����]�^��)��K5Q��8��w|x܄�R(�߸�@NJ�*���.I5��C�����o 5����k�Bs��H�=:2���	�:?���$���l���*F�D�&ʴ`���ÎR�c��<D� �-��[n��o��0��"p�_��1aaa֩�[�G�e��"S���u�
����+v?���}cIv]�V��["��U����ׁ%�d	
��A0m��Ph˾����i	�=m�����'�s�p�~@/b��)}U�� ����K��&K���*'i�q�.ʠ	 %n����������gʺ1B���{��U��L���^ z�ZeWd	�b{��`8�³W�l�Nt���?()C.��c����Jqs��+�}Q(��bbs8`jB��|g��P(��3n�r�A]T�)���$�I��".��"�|ZJ�s��]���E:�O�і�tT�Q�t�gx��.�Î�6��1�i���m�;����q�X�$��sQ�p�`���OGF��s�([�	�:7�ֈ�~] ��ĥ���v�����⟜�[C�Z4���X�/�T�J�+|0�޸[���Įԅ1!���Uօ�A)ѭB��EjXt֩�����-�W�g?�У�Ix��=EW�^u+����c?�%X��xB���IbQ����{�*�fi�fK#���GGG����X��WB�~WA��W�:��&ƜU��
@4����?Do�%���i������ɡ����.ז=�s�NT�
$?�L���n������w>��pOF��J1Ns��nb���9q�PfK�r*�aǋ*ҩV�#ցPt!UX\�SRbt��3���3�M$�L�n��
X10�����Ę���#� ڣ7��q�O��z#��߼R�[���<�T����5~�뚙6ڊ^�	����.h��z�VT�4�6<�e����g��nӿ���/\�rh�C���W��^r�����6��@e� ���B�D6c�z�0��(
Y�
���� pݬf/����Ry�a9�tr5c��>CJ���`o�6�ȐU?v�IL�Y��D�-A�&=WD� M��Q�pU)r�{�{

!��#�;���[7dN���mX��S�A�H��r���}Aľh!����
�;K�4���~2��	9��N7Q�vD>t����g�ea>�!�Έ��E'~"�x�>h��,u�h(1*ڂ3#�x^�r6�u�0�'�U��{�4�)"�Qߝ�tk��H��W_����� ֓�5�U��g��K�+�_4c���_�Ah�(1�V'��]UG��}����&!�gS��N<���@/��І���R���b��S��aJ��"�h�M�[`�6�s�*�{V$Je����tH�Җ	dC2dT��cnj�2���8�H��os���x�$�9GN��Kl��𢡊B���C��R �x��0׃�4F��u�)���mH�~��e��m��|�y��	�*��>YFF+�6>H��-��N�/����~+$ǵ��x��f��Py�ڏi�5ȄBTr�t�.�p@1� l�NY����\�9�'�h��m�22^�u�y�U�^��*D<.�6�\�Q���c�i�<��&x�Ω��gMT��\�p�V# ��;L_AQ��؎�4�C�5j�K}���U����=;�A��H��+���T����v���>�gBm+J����^�d�ᎇ�������.·���`�}��#��m�M(��92�"\,;K逎�!��̙�'�k�I�׻5Fn��bTݲ��D��"�iz���z�L�-�9�rfF����~�
�S�<b����=��Z��<�4�T����[�-���DT�3B(����K��.m����|�\
j����0�\`��t�������C�Aa��>�+�6/��,4^�����*��� ���}��}d;&�����xJ�ء.-�sx�.B��N(�~#U�>���}�a}���x�7g"Bh���+S&��P�Χa�{�\�w#۬A����Xc[����X445'O���>:��j�4h�A�D]J�E�	=%ƅ��t�{D��]m`W<_��K|��-�<�I�u*��.1�C��)x�Ia���Ȝ��Bn^�6`�je�x�N��r;���\����"�	�1��_�⓵�kZ4?!".S��
L��h3D�⓬TcbD)��N�YY�"Q<�D��AwM��A2j���J7eKbX$"ǋ��Ί�>�D��V�v���(=���d�P���o�նP^��ߘ��zd\�⏅���n���^�6����緺if�Y��,�/5M$̭|S�.�V�<�H^ؐKd��c�hր��c��((s� \��S�EWƌGi��7H����FP���]�Z��Hc,J!c���WD�y�nm�X���o*E��6LH� ����]u�qˑN�5=�i��'����Z��w	φ|��
oK8�v�$�[��7�_��C��2�;Q[u�
i�	8<����b���ⲝ���Q��v�n9�6�K(��\>���(���Ǭ������;h�ӡT��00�[<�t.�C�P�s�l�ǀ�(��.;��.�.ׂ�f��P��F�_K,a�W���Z����gx;����3�O-!Rl�ݑ��@X�k��L7���Sj��:^"W<�.��A_oŬM���u�S_���I�E{�vI�IyI�����3�I�C��.�-H��R'��/��誧>猎�J�f�ڌ��X�|�)ڛjb&�"�zJǼ�Tm��8"�$6{��E�g$�a___7h1(� Em~�6Qlh�-\v��ǌ��� �ֹ�!n@0��D����B��Rï�0�Z� 34�+J4q�.��s���GjJ���7��6�`}�Ay�>���	;�����^�ʶ��%��bE��&��p�|����J����r�|�܁�*^)We6�!� W��i�S���������/ ��9���I��:���:E� cu=�}�2�;E7��2��/8��PTB_���r)@[����y/����H�vA�6�u��8GnБ�$�5,=m��� ��P�M|��܋�a>��ȗ�d��`!�
���i+�C����z���!���>������R���Ĉ�e	��e,���Q��@\\\Q
�N, .LI���r5ǒ�?h�N����/?�6�5�������glb��p� pp`��;� ��~Ӓ)��/k՜�I���\4J1+��t�>���->C�6�x��qq�3qy�ձ,�GP�Ğ�/?}F䳔O����赎Od��>P>��p�d�E�-i"��t��W��D��7q3sWL��4�
J����S���H0�Y�����RL�FzĻz��P�9�-Xh��sҷ2�L�a}��r$��(����o@�t$:}vVe��v3��̚$����6wn�Z#�Us�����S��bz9�b��rԉ]H�`^C�������n�I\� ez��
����Es���E��3�Ǐ����I��nb�1(��'�W�:4�Q���2��5��5(W5����}���K�	�gn�"ӡ���gj�f
�rW;���ئXˎ+)����@]{�>I�=a=oh��sà��~���D���k�Q��et�&��'M�����ܷHj��߼Ÿ�7�z
�qLIŜV�8��d��f�F����!/�'�v�x�0�9V:�n�0�(y���(R��N_z��i�:7qziV�Eņ;E�D���F�SP���)g���(y�O��ys���;Ґ�= 3��V�a�����26is�J�11ty�٪�NvNl�S��w�	eV����J4x[[������Q�kj[D���}B��T�^v���Z����f�_i{%:�dj�(���,T��D*c�n�{�Vs ��߀s�q& �ɻS:�*��B��iuy_�!3r���Շ��_�^rqZV$+Ж\����7un��M ��@�����E��G��VhE[��-�q\VQ�=[EE���I���������4�d�i�|
ǯ E�sp"M*LzXn6��l߄l�_4��Li��.0�'��_,;�<��7z�ƚ�{�"�f}rFg��F'�/~��" }w��>-%�Y�慽u�9�A����6<�� k~o$/c�:t�@Y��zеԏ5ۉ˪���R]�ۍ�����[�l<I\t{٨V��{3.n��"8���"�d�Q���������$�4��)����%�)��i��z���Y���ϯb�4���+��I���k�JWĺ/p
�X��m��>���3s�XdY��s�"���xן������/��ײ�b律ⴵ&� ��ZB[��_7[��ˉ�'���Q??��������d/(�u�,{{���R�(BHӽaB^GN.�T�������-X�P����Ai���0��6�D�ӭG�dH~�Lfʇ%J��䛬D����`��`�KVQ�w��;��|y�������L�u��1�9��P��P������䀹i[���-s��S����I��������y���C��e.K�tkϓ#"��.�՜O�x���I����]��KPbӜ���#GrCo��.��@�H�~\cZ�� *)Ɩ,��-����^���:sI؟q�UQ��d
�V/�����c�M�V�tc������jv�}��r_�c��Vp��ag�-C�&%?낌�2ΞQחQ4|BD?F�s��ζY.���K?�x��~�$	�MZ�I˧?�I�Fm��y�����Ͷ-�z����\l/�ԁj�J���7�jS�7��_C�F��4�d��֒!��ۜ]?�������|J�5w��A��Ľ���nH 4��/3������ ���	h?/�X?��q�y[�g1�s���+�b���\��R]� �p�_3S4�����|�`��6Y�/�Vp�K��~d+�]O����'�|�VW�d����=×�DU����>G
Y��d�tYsb�I	�OO�V�I4B1�QJ�"߂����}�)����� ��b!����1�/v��"4�3T����dn�7`��"T��kj��ͧ�6dY�V�N�鿇(h�Z���a��P�#���N{��&�X��lL̝�izw��^���g�т5I]���r)P���j�EJ�{8q���O��{���i�Ґ��Ldg�L�!��z9���3I�S�͡�!�Lm���+�V��C��/�zsǩ��H�n���xr��W�44�Ox!���c���P�4�7w�N0�	բ����l#�?��+�[�]������r�:HVXۮ'q��j��#�:���F�����Q�ݽ��g.���8�~)i�Mԅ���{.Od�	�F��ͮ/�� $�
��Z����Cd����I��v�՘�d�P.Rq�n`�����9y���-b!���L�Q2�𬍫7��z�&XL�lҢ���͛-j-s��TfNaaaZ��?]���\�;��VZ����=\��b@d��[���[��O{6p&�3|DJ�$��'C���o��c�8��E\�*-j�}ٶ^�7�)Z�k:�]��G�"{�bּR�6]�w�%�e�F@�~��ږ#�k={e^{��M佃�]�O��b��ݍ���G���xKP����]e�n?�D�v�J-�G*��H޿���C�'��	��F�&kE�wT���5�Q��ӱ�]�Hjz6�<6�ҁHT[/0;�5'����')�i3�ޛDQ��0���i ���"�p��\R�ս1��=a,#�eVw���+�ߑE�U7)�6�Ns.�1M���y��&g�ScHݟxm^�v"�囧c����1�W_�;q���I7�秤 �e�0�. ��!��̀,Ϩo/()�<��o�@$u5��e�=�L��[������3��"������5��hTD���T���[�#���b��R.�6�}����܇C�d*���y2�S�f�b}��F^��g&�_Ify�\���Ə��b�a/(��͏�m�3X�qN��h��w�9?�z+r��$�T�l�&y��ȘP�`ˎ�#�7�Uo�����^��Z= �3�%�ۥ��ѣ�T�H�;��~�M0���?gL���#I5mK�
�h}�c��+�ε�w/������kg��'��h@����h�VE��jW�B���X*9���6̹�^�E^]�GMH5�k���r�<Sg�BRS����\>V5� =������͊���͙
�%�S��������y��EÚ�����4<îs^�sB�;�O]b�i��#����tΌ$կn�����Z��8�39C��\1QrV�F�&���(�D5�	F�̇�{<�I@luK{��RpD���d�C(m��1@��jD5�zq!��q�
wD�~,]U�+���w~Ո�R{�9jο3�3F^�G��_��S	�׌<�T��_*�9W1ƍK�t�l#.���3�%S���]���äΥϳtJ��+�ڟ�fA�9��.��ƶ=�X��a[��b�0��.��1icZv�=4'U��,�&MΪ�\5�����T$iX��齦�II^~�:��	��?�4����������n�܎�JY狐���E������ ��'�_m�)ɓ_�@�&��!��A�w����Zh�m�TzB)\J'EL�*-k"'��ɽ�������kH���(���j���<�'mZ0\oh���?��lI4�����s��&p�O�K�鄅|aW_~�:$�B��=Yfz��c�W{�z&(�݃\妡���c��v�֘��HA�M�E���݊JI��ʧp��f �C��j�z��GoN0��$y���2e_���w�r_(�:�`M���^~��q��u|u�����.���2�;d�v8���D: ��\| pV�x�=qm���'[[�LC��E�Y�ԓ�����9WI�������|�������1��Qf�}�s�1�M��W�B~��n����y��>O�W��{c�h��f"���"=�$U�J��76=`�ѱ�^^<���7���K�jo��p��N���@j_%��R/a����ݤ:�w��=y�ş��;�-��h�F�0��� ^^=i�W� <��_OZlE����Ɠz�o�ym����ɚ�X�o�o�U�u:�E��*�j����2���[v������h&Y�br;}�K��a�?�.�F��F�<)��ꆚOUj�
�T��F`�G��b�X�'RIqX���䥟w���z������|�ΗG��� Vhc8-vo)Y��R�P�C� �Ԏ�����������Tְ�Z�ɢ��e=!,S|��g��|5%��t��c�fr��(������9�?�*���dpKs�4��_R��F>��z|2�2Պ��ɾV���G�����!��m�:����0�C�򷏯���[��,-�W{��垭IQ��ꬨRM�D�wW��6�i����mq_�o[����\30`rt���.��"G��$��w6xl��&�������?a.�,Rk0���Z���)�r|�ț�H�"���5��C��̀��/?���l�GY�al�u?t�=4s��W���7����?B\��'%�D䔶�,$�Ψ��ۘ%��0�"�f�C�P<��~VG��F7������*��oE@��>M��q��R��mR���E\~�Q\ET���q�����`C���RSW���>S ͹#����<59z��#^�e���ڒ���2�SXJK"�6�9L��|=����hH��3�k��%���\^m�>Q��RF�&ҕդ���~?	!���k�?�H�(���/��x¿�mˋ;������ |o�U**���?>���A����nw�s\a���������f ��u�Tqc�����	0�U��Py��6F���Z���ړ�"��R�%�Q����׃���))� >��:��_����A2����n��u��E��|6�����f�.y�����E�ʿ�-�$=V\cmRJA:�U>x:�bɘ�\��UZ�T
ō��;� ޤ%ݸ�<���i*BR�bJ��-�'q���l]d*��;�5C[�D����$�C�ҁ+�o���&�0�1�M򿙙�b�!��8ȝ�_Sd5���^X���)���8���^K�k6����Yb�;7tU3o���Q��1�G����b�i�@��.Ss�`��*���f�B(����>�mX�8M��-r�����,�c6�}���*��MXwJ����9x��7�� � ��7j"�Ú���st��P*n9�B&6�)s8� ��ǧ��
�\]T�%�16f����S�7=����lT�L��h���m�y��ƩfΔ#��U�%�lip�)�S'���o��9��y�����)�z���0-ȥ�W)��[�ѷ2���9ØB!{��t*�HϺ$M��zu�Cv6��=֨����{��J�`c��f�,�'�u|o��6dFv;�y>�5 8�O�-���6=���؋������=�6Rn[#�R��ߥ��t���Ly���7v����=3�9�g��,]�@u4�d�t
��4�g?��K��
Ƚ����?|�P{�
DnD�� U*���0������!ޑX�֪�-�"�v�o�Sy{��B�p�fE��_��K*)����� hej�l���}t���:��j�]����C7��w ���@ͥ��Y fRf��3Mv�K�;[�M	c��6&O��4zaa-�%-��Ĕ^�B�?��N��<cH3�,���'ͼ �������u�b��pE\�����ƺ�����,���|�v�IGn"-xV+h�&�s�.�&Ś,t�B�������L��v@m���o���'��U�oN����~�*�����$}��@�:��7"#�v�����q4q��0.L!�ܖ���tNZ���YI|�̣�PԒ6�����w�}��ݚy�yC1�w/� mP�ܓ�;)��ܙ���t�ӫ���� <+�@�bm<��^sZ8{l('�,��sڧ�p����1a���Q)�踁�-*��K-��,��R��2��b�,h¬��`rAH	��[�ҙ���3�-8���	@߫
!�Q�uv�T����j����B�-�$l5�]GN�$����A���&=s���VD���)wܥ�8���q�;��X
��E����ωEĥ���@Mo!��m9I��1Y��$t�b�o�����E�M�al;P��C";���� U�C�:��|��pa�HB���0��FM=�l ����jF�u�uZ�,��vi���p�9��0�����%z�����4�3��`O��P��g��zL����Qt&�ET�Ĭ2TN*d�I��Y?��	�b!��ͭCW(�K�0��Z-�����~� ֲdyV�:����V(�|�%�~��V8��If�y����������S,�����`�����?M��~0��d$���a� ��4-�9y&���=4a�}N �(d������Nv�^����b�C���񎬟����������	�\���vkŜ������H�Ǆ�=�����~�9�Sh;�V��J����&j?_a��8�Ø�% E��(��`YP��B}L^�NEg&�nc�V��Q\m�R�ŷT���	���E�?����L�(�>L{���R��΄������+m�6���d��ɦ�<dz����Fؐk��
�^��������s�:�Ҟ�+0���z��d-��n�n�Ie��*e�
�K���u$m����.� �q���^7&�����#Y��I\��Z!L��u�5cL�/��]̝��<� ��wi�H}e
e��n��_��+�%!)��[� ��dٍ�SF��Gɿ�9o.�>��c$|٭!/S��]�F��*vC�JI�	�صk�VQS��*����HܸS�p�|oBߨN�P�M.����p�fj����Z����3DP��0����ʓ�w�U��#��V�����B�%�G��+*���,
οπ�O���G%�A^j�׋vb6�H�/9���k}��jna�њ)�9��./#c�5��&M\Lt���96g�QaJ
L��%�^��!8�龘ZB�g���GB�%�9�{��κ�Hբ���8ti��%A�|9=�<��>s�6�ן� 6M�ⴲD���s`�YQ�����c�^��dOk��v�i���&_�OnZ�.SrbᦹFލ�$']��Al�@!���ǡ���봜������FV�'��������0/�w��"o����ڼyϳW|M��5s8m[��ɾPen諔�(&�K;i4L4��L�,������J~���M6��i�֧����}�Y�3�dV1 o���u����]!q�� �j.Tg=���=��d��p���g���1w���?NhU�l�����ќ�L�H����ڌ4�kϡˁ&��7�B�s8�@O��ّFޯ��:� =�-���:�z�$ɼ\��d��D_���B�Ml��%�r�'{�ԣfL�
�Y���K��NHRc#�2�ˡ���0����xtm朖����H�l~�|���p���IQ�r"S���N"�A~���i���oa�8�qz���p�͌���]fZ��1��.���d��gn���)d��Xa\ߤe��&a�L��"A�փFB �[�sda{�k����uЈ q`eG��VM���FQ�Fu��C�b��Έ�VFZή�bw_����e��M�"��e�;PZ�E��j�}��+�'W�-�J��
b1�[5#oK=�,#��*������+1�jzV�G����}��O��,+�%3���fŞu�����1ov���x�x�8p�������nV>��Q7#��89����]cX?eSw}��F�/��l�er']N�\�m������r�	B�7�F��q:EW��͛�]o���06�*Rb��,��iz��=_ZG�G�ٕ���N�޹�Ĝ�I�^�5�(l�a, rK�ø.����о�FZt��j��;%��p���]�ts�27nt�,����
V����:�m��*����F�@,]7����}u�����j;�]���m׆��Ɉrl�QU�����O����o]T
6�j�49Wd6;�Q�J�?�.{�Ű�+�Sjˠ �/�/��?&j,&��W����6i�E���s�X�ŀ�9sg<����S�Ӂ�����F���/���Qc��v��R���}�����g#�8tk�$����f��8"�r@�>'<��;�u�@pC�@�^�
�K�ls�(����$������M�,T��ϰ�zϲ�ȇ��L���ƀ;b���%�g��Y���f�]��[Q�-��1�U�EQL6��(�թfU���T���\kdb��ͻ���LS(J)5�w���J���n����6M!�=��w�#Y����j����^��?�:J�a7���e0�m�H����{�R�����f��;S*���ef�����?��	���75 s�x_c�ݯ���>�G�;Oy#��|F��j�lf�{�ύ���puˉd\�lSwǋ��I�����"RF�/6�F��ps|��d��#i��H��-���DGq�����Q�JN%�L;�S����ڔ�%ǣ�+,6��:���w	��E������?R`����%�c�uĀ��+N6�4��9�T�������7�V�_5Vo>,"���2�ߘ�N�������"�SQ\��N�MV�LrG��/�Ͳ"WS䂀+���by/�T��=;��Ks��m����t�-6z���7?�e$�����/���>E_�k������5���}j@�������A߉E=�X'����j2442�I��I##����a#�<-<M���l��F���'g&�F Q������O.Pi�^�)Mut�A��޾L(_�kV���ylyF�qi���<=-�O�R�/�U)&F�����$u��x��Ɣ,����0��R�v#��CϘ���`�xJщ.��RO_��N��V 0���2��dY��Vj�ڥ��������+��j���R�ȭPYn�'d*S�.�[�R�&���=���P��ص�cOc��dP_Y����e,��93����?^�s���|>�����<�9g2_W�2CB�l8�o �]��b|�9�zŠZ;�'�hͻj/���3�~��^[ ��N��.B���Y6b��̥|�8�S���&ùd
U\�%��bE�D*�c���M?֏ B�X��)-�0���M�Ȭ��;�ڙT�J�d"7����jޯ��S]�w1�GG:���)?�2]�*��������`I@�лf���+[�<��B)���ܢ����Q�r^+j"�𷠹Xm���(��$!�+bI)������(j�k���46w�_�B��A��r�\d�q��Q?&�s �6��n��D4��Q�Ws)1��X'򤨅�+�
8t�[ӫ�SXb���������@UX'5�w0C�p�G А�ZE*F�������a]� ������^��q��p�.���	����6o��D[B�m�掉Y���k���5�z0uM���9eG��H�a��l���ޥ��j����a���'do�R?_���˾T ��韜{�OV���TM%C�(���x�ݰ6�$Ѓ�Z{��8�(�>�ܨ�Li��jP��[}�r�Pڸ���;/�,]��>Fn��
��?����_"��
H�f��?_�~*Ew�fFa�1����L�U�8���I�R=R�1@k������S�׹�?J
Lj-G�������������Z�:���FB�0� ������2TZ�փ�i���s��.KͿ.%fS��\~ig�\� �[���n�Yx��$�3��m�& ��D&C\M����f��|�)wZ;�a�Y\:/����ї��f�x�X�+�i����B����N�z��1{ �_���w�8��0�ެ�#�A�L��g����.�տ4j�oٔ1�u>��|���ɧ�e�?�kdeK	i��֪Ň���0%礴V��P��Ai�:rQ�?��hX-YC~�
Z4b�����2�)	o+(i��|��a�e0�<]��c}U�8o��\c>Wؼ ��oh�t �|�	���O)Fc3瀫�}+���,C�V���]�6pV�Tc�E2o���a�֭Y�$�t���/�l����'�ᗀ�S��ѶoX5Av�����ǒ᪷���?�\�� �F�j5���3r�!����"�#V<�\c�����X�\�gN]�V� ���s�����tpV��Ӫ�%�\շ��[N���(t쿙A,A�y�h>,֣��*4��1
�?����!$-3����xP�~a~�&΢��#����pb��q��3�N��f�����9}��<��DKA��(��]\j�����!��ak�]BL^�z ����CQ9SCg^���<�7�J�H�=��|4��,��d��� ��7�գ�Μ�y�u�J?1�`L�M��=&_F�2����\TV���Z�\Yˀ��A��j�9��9e�"8[�Y �D�M���f��`�:}Z��Wr|lq�$)���s2�φ@�n,���R�$N,sѓ�@�4e�E�??����*
|r*G_mīڇ���꒙�t��	���M���<�ɪ�f�jf��&��Cq�z,#M�0cMd0��P�%�4i���O�	�A+á���@����O�0�@����gA�}�������Z��s�a�$k�'��vJ~c���rݵ����DK�|�]v����d�� ��@���9[�"�0��S�|=�. ˑZ�pM��(szq�.�F:�\�&2��EZR�-�,���$�?H�SǀS�"�M�\��6��!�)�E��5a�L0���u��t�įP6F�
=bw�� �m0�~�-���ڧZ8���v0��w������@i��~z��se���J=Ȇ������, T_җd���Ϝ�MцCndH��#�Cm�V��)�>��dU`x&��{G���g/��E3�f3�D�$�9xڬ���F�Zm貦.O���	�b}
3�km@`��DG[�$x���#$����y�P�E�[8��Z�_�|��b���-
��`}1ZC���aH<������F3�Y�_W^<��rȚ�JK���m?��6�_%_��6��Q,w`o��l���6b�x�:�y(�G�2�q�U�l��u$����|�:Փ�Ű �(��U��$NS��+���]��N�XNX�k��9�d�a�=}���tvB%6C߰�B��0`�9lr��#-��[�b����x�(#g����=�m����k����s�/!��9 p��t'��d�7-�2�6j�!���
�#{5��ĕe����O�G?��4Aƥ޶pF�߲r�3�9�E_���@A��0c�-����(��=����oQ�ɩwJ�{+y'yAAJ�Z�Yz�~��K@�@���{fЄ=&g���3�~��Ф�\5��uk���h�G©>Y'�Ճ�=?&��)�D���.�(-�{�Y�? �2�`����k�3�q��Dӟ��|vs�gx�)|l�� } ��������-]7��,G��G܇�MY ;r�l��כhEb|;�b�\����)!��jKoZ��O?�u(9`�o���w�J{��_���La���CO�r�g���뫺9m�� ���K ���|d�ˈȴ���}����4�ǋ�vEU�FNj�U}S$9�(����Yf��v�_$Y�&����2c�׭?�/ k���:�{�K�k��S	�H��=	�8�w���B  �h����b���'M�*YK}U�B)����z̆�	4@�#Q�M \}�r�غ�]�W��!-�ӥ?9i�	\Gn���s%�X�M�}RV���6#	�)��0�X��Db�M�eΠ�*��� ��xr�����ksx�id�����K�j��;���Aw�i�=��9����^�7+��ٖț��Ҷ#����P�3��B��?_~��4X�;��k�H��D@�q �� �:�UVN �a�M�23�6IS35����ֆ���W��%���\���
�V�Y� �Z��YN���Y�!�l��쫵��D���[@�-V!��H)�J��YZ۷V-��ؐ3l��̩���V�,4�P������0�C>�Ӿ	��$`#wP=�cy���
�-��۰���澯wҦ�?9�S$����p���%jb�У�K�Z�͋����G�{�r�g#X�d!�7��$0�D���KK��]����7�,�� ��<��O]�>�p�`��.9q~e�L�+)��B��O��z�����>${�ݪ��rĦ�}�:�iZ��X5"fK��2�n�oWz^h�Ð�t�
v+��	��9C�{��Z	��	6�/����7:϶d�BGc1'�p.݄Ο�n�]�[���*?A�dx�����8�LT�@<��i����f��H_������$rIx�1��k��Vh��#�<�@��{�8��}�����(S�qp?�(ѕÒJb��}sף�F�8&��E`B>
�i�^1�K���a����S�?8���t�u2�M��"�z@�_�� j7,n�t����$�t)Rq��9";�2��[;Y#����i``��^�<g�R�2K��	�<�y
K�G�E��u��~� ��i��61u��:�v���ם�r�D��[��/l� ����b���+�'���d�n���}H��1)FTׁ��<�FQ?{��i�����g0����� y��f���pW��<�P_C,(_7�·�SY����\���	�{q�}X�
����!�kabͺ���v s�Ь. \�ՙn+�kJ����
���;1��X�vԎ��\�M�4�`?�El�wW-(:��T�?A"�m�������6�ΐ��.�{�y^��d�$m)<���bV�n�����W�t������#R�
zu����,��,���1ޕu0��l[@d4=�h����z���P�i��e)���;G��at��^[m��cW�kq��mZ^蝄�<b��t����\4�G�y�Z��b������*uy[�Y��?K�DS"���P�eM��>.��oV�Ꙁ+�H��i*��@��ϔ=��B�q��<��I�v֗��:g-��y*���U[k>�.�V��̑�]��U{X�> ϱw�.~��ŗ�2����E�.N��Jv\���(��5mn�T?	��b`�&D P����Ta�Ȕ��^��Z8DՂ����^��ΡT����:3LxG��g���Y�~SB�P
��p1��w�sL���i��5�> ����J��/QM}������Mln�-������o��b��D���������Җۄ���J1�91�&/�S
�Y�·[;���j+����C���t�cz� S���.�����Q�%|�z�@WV��~C�œ��!NC��0�GY!�C^��_K�a�]�� ��*��J�3�R)>=�,>�s��a��6��f��ne��0G��(�^� Xc3��Hb=��Nd?��+��"�Z��Sr2���ć�q,xB�!���38�.�R-I�-(���g��4_*R���S�����Ю[��=K$p���eBa�)7�\(n���o�i���hi^�ILN�)@>��z��~k�2�����U/B�4�@.�'��˖8��$]���� �PIt���V�9���~������NΊ�LU��I[*�SN�K��N�C �j��N h#f�FL�Edi9���ޥ
˨:�@��ҭ�j�fj�S���B.����6��ץul������b��76x��r��P~.zL���A+ٛ���/e�_�U�綱p����\9V�Ҝ���4�m'\�%u����'���!o/j\����ÿoy���^My��G_d8h;�o���-���"ʚ8����'�&T�&�MI��9��`�ޡ�%ʸт�S��>��bE��;�C>����1�d2V�=.|4�-f�\� &�xʕ$��D�N|�����*�zj��?l`�~�Z��EȜi�/�� '^�;H��Eќ��/�UZ���7S�S�����{�ظh���Q�����˫1��}���K\��?�,�:*eM��!-R�%�nW2[�!���������B��T�yl� -��e�-��m��瑚Ѷ�UCh�
�3&�Cv~W�E_���ު񱓸��cp��.É�� �b��r�}�,�V�7�~WYխNei�]��ӣ:�lI&�X�J������ǵmЇ��;A��<�.��Q����Yd�:�
�%3��m@�yCغ7��㧱��2��lCC���R`V�w����BB�9�􀇗χ�`���՞�g=��kxn}᪤|t�Y����dAvI���g�ݮ�*h��
�7�>X$�3ະ8P��vi��(�LK�����ھ���W\F8��p�Np#��AwC��sĴ��j����q�I�E��:z�>����FHb�n�GS��y�E�R�t�J����O���Zb����p�Y ��o�7՟���yr�p 8�)�p�$��3���N�a�~z?����K�-��������x�w��V������񌚼�.����f����PK�X* ��0jwA��b��
M�C�J������3ป�*.�Y0oY@�u�٠�4��$X���G'��Y{(⋢:p��3%�^��Nf�v�z�P��A��"�l'lE�;��Jē��|s)��\��9n���_f^$zs�G,߽d�hR�9$�3��Ch���-���-�����gb�a�K�eee���d��ץd`��[�I;��`� �}O� ��HFx{f��\�\-'���k�佷�x��0^�#�ֆB�vtt\���v�x�4�W���F\���j���k"HST�	���\M$���~��vq�+%w?[a��d��%V9w(m;B��/�Q9D���YfU$yi�eX���hP$è����ג⊊�fX$��V:Û򂮜����<P�
�,G�/`q	|�̟��~X�,�JL��rA��چ������J|b
m��H�e���t ��K���?��6��~�K���3�@+)��f��%��G�C{�A���$sd�]f�%]JJ�R�SOi��q�ȇq�!��qP�i�_���ȼ��h���88���-28��z�6b���+�XB �ўJ��͒>�w1��e����q� 7�wZ�e��)P+STTb�����Ҕ� ��.쬝΢0�߈qUڝ�2r ���Ӏ�]��@	�l��\��~�,��k�M�;7db�kZZZػҟ�.Nld+�3r �Y�_�R��>� ��ޗҳ>i���V��Va�1D�E0�kϭ��a�����EC� 4���DE�A#奂v�J�a�ڤ�U�3����x�К"���rに�srk͈����y�P�aH}k3π��S��
���{E'��t��_C�Q�g]9�\J`��G�ť��lL����r%,�9U�����͏����U�M�]��#�1܆ϓ�8���6�:�FM���@�Ȧ��K���>��7,��?Ö�,�1��[OU+VN�)?�$p.�q,��U������P�����,�9�������:��E)�N[��=�K�|��C��uL#,�����z�f� ]�PФI�0�']�ʹ�e�g��z=;�ٸ��Z QhB/i���<{����������hd��0����9�����*辪�j�ӏ�|1���Ɗ��T��� �k�Mi�z9]K��}πG�RR7�	�㭹����ˮC3��άUY�%� ��)���;ef]b�?���2	�����6A�����>*%+�֍�j|�y��Hܣ>)�3�Pf%��JSo�~T� <�=W���j,`�Q��� "E��(˅8�`bb��3޶w��J�6���c`��^?^�);qV`]�;���M�p"�� ��[��@���ʡ!{~�;	�:�/l�{䇟�[�Z���Es=_���{�=�րᯏ�zP?�SA��d�*�>��"[�7�^��%=�<D���k�������"� �[��%�Ƭb[�,�7��U~s
�P2K9[}V�wƛ���+�6�M���+2�|��M�ڵoƊ��4K����IY��X�P�|���Cc|m\��2��5Rzn<1�/:_�(A�AN����K5�r���z�#e��b���\Ȉ�]�fK����a)ω�iLi�Iݦ�Ȩ����Y����n��4?��U�5d���N�W��UĞ��&'�p�+��D�GC� ��q
i�%F���ٰ�z6�'���B5�Ĺ5��W�3԰�,h�w��e�c~'�����"_1��.�'�����	�
�^к��c��d����OQ)Y��sb"��7�Ŏ7���Sn� $���e�yVh���IÔL�����(8l,w��X�ΗF��u
���q@NG�w!�g����l�z��^O�3�{c�<�N}�e!�U"�nZ� �giK��1Il:o��3K���Ok�=C�آ~¼ҾT�8f�:�M�(z�mL�� ��bJ$�$u�`��M���Q�g�k���2�g[��6�ǥ�2��p��[���%&����w~�B{=�&-��N��f���Y�m��s��$a������x]����(z	_���jϙ�:����BM��-n�I��#�G�`�6�z ��f��؜������(��.��1 ���Ng䅣�3G�D��A���'1��Ǔ�'���
iU�YJO@Z�נ�*��,�X.�MR����=6�f/o]P���8K,;�����H���=87ϓ�48��d3�
�\Z��V�E��<���Ѡ.����5SWF�՛�ڋ���oa6ܨ������ނ�ٮ�M���?E��Oʭ��0{o��:A(�O�*[���7_��,X��DȧB�w`H�K�R7ΰ�����m�f�ΐFjir_h��w��.�����=���TjZ���%�)�)١�����kJ]|=v$�"�t�.�B���(�d6�q�ɦ�0�'_��[�X�����k	��S1��n}W�X�֐���>��ڑ�W6��K!H�x�N��|��̰�jf����q�C�`����w8vSQ1]��+J4����:�^� @B��xX�>�O��8,B
89�nS;i���k8V~���[P�GGG�0��Č��a�E�<b=h�$���>E1$�%[��s�S�v���}q�5��܈�J�R�ܐ���$��e"H�-Ѵ�5�!�~����*}~��F��(9RӔ%���!��.�VT)`��_�V�����/I�7�b��a@�;o�?V���<���������l�Ѥm�1&�~`idd$�*iP&�E�cAJ�����U�<����� �`��tZ���z�U�8�Ջ^����/�=�	<˩x��T3 ��N�k���G�^�_kB{z�h�FD ����~��,���A[̈́s��J죀YX�pa�Z���U���d�N-l½a݆���7$�B��'v$����x�!��Hn�If>���Xgs��%o}��"p� �,2=5��s���s�%�)�#�rW��Q�����z��)�b�Y��>x>Z)��7G�y{F�ft��złA���BP2bޒY���& ����@���$Y��r�	���V|��F�n%��B��t��$@#��#-���0���v�?=��c*q7S��=��qR���O ��n�X��ϮZ
 8/���j�k�`��!���Ub�:�ښ��TOϜ��+���SF�.���.�a��(H���+�~�9M�7�Y�BMRRU3�Dce�>�RRcaշ/��봣����N�r4,���D���><�l#��9�Ÿ�]�4���T˘����
y{��T��>���/Q]���F�-B.B�NSKl�DP��`C� �ч@l��ǳGǹ��}��齾3zL����{��>E�}q�,53��y"���3\=���������x�A�}c��?�k{�s�ob�f����
'�#�%���b��7㑟�^>!��PS�j4|^d���Ic�J�@�x�L�����<�0���j�Q��5��^`H�MQ&��4�!����O���"�ow��4���q�e��m=�aV���W��$z��<�.&�UJ"iOVti�/�����8?�1�2�4�j�jW[��lDr�䀈`�1�/���&9%3IX�
簫�X��i�Y�qx��G����.�y`��g�{S�e�
Jr�5�>�#�җ�NƜ��2���'�
�(�u�;d�~����m�ˌ�b�	]}�!� ��t�ϗ9�9�gv28���Jf�r�����c�O���}u蠗t��!3^KH�os0?��*���Z���H�&=9tUFx��mUxj����j��j����kϮ¬����>�)@����Ƅ�s&+XL]�K��Ģ�\ϒ�F�ӏB
@�bN��Y�#e�pR��I'(��fr	ܛ�K��[yثT����d��}�lِ�O�x����3��;����888(�q���^�5��(*Z{�.Q��L��v�������F��@N؁f���\�%�|*v.���rD}�PɌfPH�{�Z�+��,��і�>���Ȱ�mmmOa�3�ᦑ����IGE,8�B�a��c&�ډՂ�:�\�H.�{F��%l�K\O�+���d��ؓ�Q�T�q���SlI����A�!ۤ�u,�"�˓Wr�;�a�^�,H��M�U(��ݰ��:�����F7>���&��ʿ@��L9
j;vBK����͢�cW�|��	���{�_�y��̜=pc��� �8���8o����%�`�f��{�����a܌�T�P�&�u?{����cb];�	�J,�X�����$��	��iry��.+*)�Sҽ�֠Rŉ���DX�7��pQ�J��$(a�-�r�>Q9�o�K��o�����BAk͵�� ���9��~Mj��R�D�S�4����ˬ����G��R��6)� ���5�����ƛ3����`<�V�u<3i,�ڵ�"خ�.�
��-��>W�ڤ�6ň&G�M	�g�M?�C~�U/I����Gy"웽۔i�;��wן�L���Tg+��A������UMu������f/�dH䣝��~�lE�9����d������I��ڧ�N�*�|�;[=c!J��x���	E'*PG��U�}���C%������k�%���j�)#e�SUS�x���y��Cu��'� . �0��;�fĥt���Z|����oR�mU��C��7"H��
X�exݞئ�J7��H����}G�᳣��a>�h��WD���i�@�����@�ދ�	x����kg2c�n���6�q���
z�������n���5?�wǙ�ҍX���W��V)��z�՘
,
���%�U��:���`fcס�l9a�j�5T`?
�W��+R�%�K �N��(]Wr�*W�]�Ӳ�<7�E�Ԝ������ �)�		eNa?�h����M6G��k}� ��n��pn�u��x:-o��ްc���B�d�Uw/�`�'�>#H��Wb�sJT穽sssE111j]���l���ۤղP�'}��������4`�,��{߬7���+m�<u�1��T��q���VH�?jP�̯�;z@�%E~f �V�+-��G���^�zT8��Drf�O��sF���'�D�Ϡ�߻<�}Ɨ&t5��x�I:Y�/�^綆>2�8�;4�i��ſ{����P͝l�\�(�˅�/%�� �
pA<�����p���&j�x��˫�!��&J�q���.o��.t,]Xdu�?�w�*h��Q�[�����3[�N���a��w�w�sm���ܴH�k���4fc����9��Їq��1�S׀㚺��|� s��\BdK<_I̟��F?��r8u?8@.��]]�3����
ٌf��<���ޘ
�k����,�߼�ؙ�}[�e�G��ӗ���B�h��!ޛ���eH���;~R�9�%#A��|[�&q,j�~yр���w�|J�� ��������2
��bJ�u��;���>��=?�{	�oW����
������^�o���G����08K4}M|���UPo �J�נ!cA��g׺Oչ�h��-��|���B�Qܓ�ځ���i������vx��m��I���*f|��D?1W~�W@5�vdr(jW1�E�=�k��s71�` ���D��D�|E��P��d����Q�$�j)�+ӗ�?ÚN>�:�,��H�<��v�w��.N,�H������Z��V�
yNOѽ�z��S�Ntc��x0@<H�J&%wYsEtf2��ۅ����dK�
)!^W�����	^�PF;�?�׳U=���m؏g��v�5�w�|A�����1d�*R_U����<�c8;�vCl�ގ�\�����o�H,M�`ŭH ��RF����:�N�!8reen����;sd/.���a�J�v%��� �w`,>�e�����y�Z�����@�G����N�H�2��Gy�(�
�!��Eu���e���3��0�.@SR���@������Fg��N*���$���}HO%|��W�NʜQc�� )����Ǐ�V�HZ�#�QO�1I��A�� M�M�O*�Y6��?VH��G�Jb� Z_�(J��'����n��G
[� 3/�j����;+	!�
[��B֟�:�%�}U��
�l3�f�*�(�|x�̋�Ê�y^A���'��P�?!�xy�(߁#}ԅ�2-D��c�X����$�>��r!��~ N�҇O�C@x�C�xͿ�g<ƀ�2K�x>�骽�(Yܹ�>��gb�^Y���0Ot6eWm�gس��u��잛\J��@M�1���
�M��д��*.�Uz�@�;Н��ff��pZw26�g�7���[��1�SR���j|B&������/��p"��*������//�g���x�K�+*sK�b{�y8NI)F����W�7��c�v��� н*�u�����r/`tw��;(2���hVkԩ|m��>�?��>E-��<�> �F�Qi�|�
v@�w���P6%2�B����;Mps���N�h���%Ǭ��r�ĆX<�#����\:�𽦀����='�ۄ��~0>E�Ja.�D�W���7��J8������G޲=@�wZjs���N_E�!bC^p��<�5J�L&S�{ei{@H�	�"�*��٫,�KX����h��Ő��̰_�M�Gu��>��1�)��NQ<PNޠ�c�"��y�xuwbt�UP3�ٔ\ӟ	�u C���0�ί[��i�����Rk���Z{�4������G��J��w�~:�f�����%.N$a����l���B$_�,�	XF��	Y�R`����(�� Wq���_�ʡ�K7!��N!����Sv�O�H�]�%,����`�&�xx�����F�B�(Ȅ4)���~��f�A˿Ïa��5ԷCP�S��2P�2`�Yj� ����G��j"�jR�|�ry)�\�"àEA*�,��
�} �����*S �*o�bO��� ��c����\[�߇!ͰS>�,�J�����W��Id�i��u^GH
^��?���$�m����4�՘�斸��N��k���!�5�m��'��81���Q?>4$��p�`��:��6�*!l}7�Qz��t����R����8��9�Y�P[�o�[Y9&I끯g�F�ID�_�SO w7͘������%�p\��!n�=>)���M�L��%�� >����C�����������Ѡ�������(��_��R@��3��r#;FC�gi�#
��P���o�}�j��"R%ol=�Qi��H!<&0ï������I..�h�CH )�֛��c�r��CJ=�luM.	��D�C�l�OL���,����Qw `P�.�ߧ�\v�5?��j?`����E�@�~���O~�ɲ�v4߽��֜eӆI�c��9,�A�7�G�������ܐ���S�Г8���OcE���ܹ��>� #������FA�� �QT���!g�D/h��Z�%�|6�9��6ZYA����K�����X5^���s�>���E׆�C�ۻ�A5�{�m�M:�W^R<:����8�����hE%dz&�%=��B���v2u3�i�TGa�9t"�;��4�L
��4V^�mA=d��п>�cA9t���N���2)��&�|L���y�.T��il[�����t�G1|�����5,]���s��x��b�!�sӻY�Dg��O�!d��E���!��o�烾vJ؆~��f���6ĝ:w�'�n���!����N��@^iL�&���UYޮ�E�/�*΢�ubo��n��Q���H�fd�t2!�8��������4L�.�V�xR����YEI�B.��8��C~3`�̾����R���RD��0�E�sֳ����y�Ri��Xj�mwOO����J�gC�@�؇��}�������i��_������f�׾~£�a����(����q3	� �z�1�l��J;x՞"{�o?1Qv�w�����	�+��8rs�n��+���5Un���M7!k���!<^���ċ��V�t1���,��YB9t�%>�D<|"OPG��s4Z(�PNC�PZ�;1��k��bib�߾�%�f2�����UI����Z[ZZ�:\� �:��4qK�V�-9RZ ��&,�;wN�|�����{�*�bBi�ӳ�=vt.��Sn�Jn_��F���M3N�1��
쏅=�T�����g�������v��u��Z�J�9%�p���	$�c���\������;|o����F���jY[[��?�^���fjb�pʫ*�{E���o��옷g����Y�'���O�.����}��0� �8�t����ɬ�X17��&��Q�,���R((�ɑ����O��eeKx$?4	�W���E;��{��pM��xm?�\����:��>�we܌�*�x��VVO��T0�	8y���\qbbbe.�o�> >��
��I'�;|�[�$�X0ϩ��k��z\JX(�ap�D���M�[��V��jqtҭ�oC��]K����������j��R��D%�4�À�sp`�א�7��\d�]SWw��j�%+�ؕ�q/Y0O	A�HP������OԷǥ���I�Hz�%��5�h���*~L�=�!�,�A��}�;~U���W�?m�
�����)�@��x_ �?=�-!E����'!6JY^A2�	���dX�R��!$��nD�O����a���}��0����ƃf�@Sj��x0Qk}5�QB��%j3kN1�R^\}�"�I�p`�� �*�@\��'���_��-)ᩘKo��$4` ; @&p���.�z��(��@���{���-�7�j���+:���ÇUٽpڜ�M�֜��`�N�-�j���d�Pj8� ��`�/��a̯�&�������fC"���J(w����������*y-����d�'�}y����@}��������7��ڡB���X��'*jI!80h���9�3�l���*��?@���K��*�q>~��0]�ꓭO�w	��΄7J�7<?���eO;����@��)Vu��m߫�[@����NS��U��;�4���%��.9%nO��)��&O2>����j�_�� ��]>�ܕ�M��T�q1����
�$�V �&�Ŝݞ����_<�;�;�)����jN+���M��7z���.N��V~P��哛Vs� %g�#J\���IpI�2�;�֎t��Z��-v;��}	>s��l�nHopXs�_�#�/�~)�����,or�'����m8鋟Y�i�����������y�ж��{�5��?�Nw�Q����-���h�v�p�_�Q��@�M��c��?��Pt+��\��������c�
�/i)ߍ���٥;�&������SJ/�MR�t	�7�WV����s��:��+pf���K��.�8_������|lg0�m����к�_-�7|�R�&�:�ۖ^+�TmSK=���H~��������\\�n+�Y���ĕ}LL;��S�t���]����L1���&V�hM`y�oʙQ�Wb�>˿�Nr��PcS�) ���]�)��s>�&.D���	�����i�.�Ja�4xݸ�Z�۷��o�O������ŷ��ʦܮG�>��0*�U�^g��a��n�:t�6(xk؁b�*�p��z��%��`�2��B���u-}��ZnzyW���O�5o����~��H*���N�s[��C��	
�ޝ�^�뵁���|��p��R������y��Z��o��w4&:z��䭖4�f�<hʣ�'�ݼW��[Fz�餯I����'�!=uHW��[I�c�g�mBI-����b&�/o�4����r�w%�q���w3����t�[`�⎬n��%�VH��N��J�{Y���O��6VD�(@z\���b�f��ү��o��K����@�F�����y8aSgI������R|��)�`�s��G���8�yr��y�9'��t�6���N�Mu^ʅ��;;�k�TYBm����vu���/V�oQ�D"�V��<�P2��4q����io���/-����þ�9���v��w��yn�̬�T�s4K�s���|]g��j��Э�;'�w�0�<Vz��)H7h���/��35��j�de�ZU�/�v8�o�w{$4b%/��i�;ׂyYd��+G:��y��碯��|#}�%�G`���w�v���<V2N���2����Mccc�U.�HV�W�k߱���{��T}�gaч��Q�kd쳯��K�-�����}�RK1�"����XA�D��q������N����|�tb��ܴW������9
�yTn�X���J�q��
k��@�?�pN����;l�h0�M�V��uv'�hQY�>�?�X��iz��%��?m}Bm���}"iT�����\��Y���2��Ƌ�'X������{1�Ҭ��fh��*�y��%�^XYYI}��G4���AX�랿�k;�Z�5޴ggx텈���r:�g�%�1-�e�r+��ǥ����h]xF*�]�4<�.+''�^�������ź�+�������L�W�K����+ߜ������>K�^+���h]���Ja �rr����<-sAeȁ�r���*m��XX�8���}n��%�F9`��c]�l����9�>�3���d2��VV��m� ����׾�nv���o^�M$�0��ٽ�r�L��Y����� �(�Fɱ9��	�륍�����5�=H%E��$ge�|�k��?�; doǏ�1����{�,��ݹs����>n���l5��󵶳��Sͪ����/�)?��>`y)�2~6�{��/�|V"_$��A�r׎)��P��am�yQ�7ͺjTq�䗄�A�w%���@��f��S��!=�N���B-�om�6n~&��Qf��k�w���;�Vs�� ��k����n���@���ҡ|R��o��{����_��]]������E�M�qi}���cx�]}�q[��� ���t��o��쾛���M �\��v�����`dd��������[䵛{}d�o�w���k��Φ�@��]�\c;�>�(TZu�]�j�O{���B�fE���M��7�#^��>�X�qǍNM9�z��������g�o��J�o,H�< w�색�j�b�B�%��P|Kw�gC���B�����	�RI�a�#�<_n���<���"��I�F���\\!�����5]�!�f�|nTh[���-96�Na��nUUT4�v��I�l���p���L%�l�����o�H�i�R�p;��oGt����F��v��wX �[z��'�_z�����)�G`��P?��i�X�x�j��v�f��U̥ٽ����uY�rRT@����V��\,]�t�]�qO�Y\Z(����n49��x�>/�7��y��0E�z�ݟ�?�-��0�~��]x����)@�q�Ϯ���vT8�]W����,�$�84���㲒�^y�h�6kI�ke�p�;o���#���a�4���k�Q�ht�����eSDˆ.����x��G��&�u��B7�P{��,&�[�B���0xpCCdܠ��B��w���#�ϥ�Hy4ix����Z�<옱��?�ˤj@A��GU�@��mHgxvtekG,�^Z�J����DO���׽��`�^F/�$^�T���A�۷�b�M��P5�ɰ���.������
�'�2~�Q<g�b���j�j��]��mz��|�KL7��0��Iކ�
oo<>7�X rɻ=I���{>��W��M���a����T�x��5����j��c0��ݝh $7z������_�-h~l���$];JU��q���6��"d�߁�;ݸ��}t���ڏ02�����O}Q��/���kl'%�;2�1��.F�w!���)��4�`���{aӞ����~�xg�.����`A��ۧ����:lJU��"����B-Л�k�p8�䉮=��ɋD��+r�x.���o���S�\��=���>G�Z��?���@�T�MP��;��]�m�?h�73H�~|����Ŷ�J���Ax�R����N;���7� ��_����r���c��zdjjb�<���a�X�Z�v���I)��{k��e�A#��3!&�
b�l���(���;R@@�`~����9�R �M���J�wנ�
�2�:���:?�N��%�S_�u��9|����U}�����>JL$v��4}��A��c��j�~}c��Yug�ȁ
0�~͵Ϧ�3��_�
cFGh��d�=<<*F�&����휦|�Q��e�[E��ϴ�Z.�*xʼw�����<�s�״�}V:^�D��s�I��'����`�"h-fp��{��c\��O4P���eL���D]�M�*��NM;����]>p����HOʣ~1��nĉ��W���]�J� �@��~�T��7�&P�?��E��͕)ߘ�y�V���A�c�r��#���U'�\CAѮ�^c������Ai��{����@����*@��_� �m��nRD�î�6IZWIX�yE��s�b�Z[U����@O��T�C`R.� � #�|�F�BDg��c���EGs��� ����������~P�&{{{#1�9�@�x�|wbk�m>iӞa��"ݠ)�r%���I�a���-X���4��;�Oϛ��͸�-�8a��3D����|���Lk��X��R։����\MMM?&��$eBr��$][���3bo����d�_-//�z�f�-��ǻ�{���e��K)���|�"\�H���\���5<��� )7n1>�ip��Ӷ�e�1
0��,�䭥����=���ǺUz����D4�v⻤ݜ�Z�	�B=��ȱ�1ء��i)=���(�0��UC�U��C�3���k�����56�"��*s:��+����m�`���EwF�����Ǘg�+W0t�h���E�=��C)����7�N�5>ǧREs��,;4~I��O�TI1y���tM�~����e���G�����%�T�m��P�H2�
�� T2mlIi24)2�d�2l��D���XGE		�mI�2��L�6Ŧ��?k��������w��:�w=�}�ϻ޵��^-BZR�A�LTD�mS;zyМ&,_�)L )�bHQD��I�;�Z�L�
��I�o�ԓ#��}��d�3�([8Jg|Qa~)���3��S��Ī�L&�vtx�b� ��t�D�/��́P|�G\��J�l:\9��>��߫��BJ򗩊_hƋ�����zf�<�P~�5x9��I&�`�#`W.x��,��8?��l�A����լ�p�;-j����u�6i�&n*��O�lL���m'o�)r�L�� �Mc���t�=�=[�t���M�'� �H�ڻ]�ˉ�������֕��$�h_����Ҩ��e�tF1,xc"�E#wH��B͵���i��3	�$�!w�+� ��
;5����o@�S���7㷼�͆G�w�%}y'��ۻr�@�^|��c�k�`���f>���餜����pP�Vvgs�
F������}�V��~�]�p��Z��X�2��/�e�uZT���q39��l�� #.	�'Źԟ>O��?�����hu��)�d��W��������z:\�nͲ�E�x�I$p�dWy��ŀ7�:���]���ng�B�o���=g��^�|Z������=�+7	Ġ���-���IH�����݌��ȓ���ӫ�e�
h5���I�ze�b�u�t����;�����ga��Y�H�����\�*�I�)��_�J�&}U�U=Z���IA���� ��q)"%��5�t��a5t�z���0�F$C��|8����Sy�-�o��*~�A� Ì���N�0t����E���~�Rė/C"�;�8�m�<�-5�vi��y�}��+U�K��3��a\�FkS>����~uA�`���˗��Xw�t��Uw��/���{Q�C�5\�k��Z�+g���&��O=������e1z!s���/������r��S��S��yk�l~ߌ���d��v�-�l��0���,;4��u�O�r{����h۳q
]Gw�����`F�V#/%�4_��!䜢���E&���dݦ�C;As�]$}wtt\�~��}�լ�:P�oϨ����U�y'���w��&�b ��.�1K	r|mQ��
������|�÷!����޾B$}�D�@k[��Н[̞�K�����*9��l��q�n�N�n�iL9�W��˅D���p���C�6�3�Y�OMg��t���5^�|7\\�AO��ݻW�-��jˉ5��_�.���f������u��,����w�x�*�̷fQ&J&K����J��	1�O��WO{s�pn�g����Iߔ5^��M���y:44������m|��c�u&'��Y:�A_����aV�x���i�����ȏ�#�*�m���wOVF��Fۖ����L���;���y;3�+,:�]�5���a����gO"����R��S�\�K��*^ tv"/7�\TL��J� Z�AR*����?n��D�teGU��ג�@�[�P*#�����5�Զ��ȓK��-yj�C�K�J(��	}�����B�����g&��q�NTWx_���pi[$3/���H�̩]WJ�u��?3��Z7��`�Q��3�EPy�x=s;����l���Ձ]J�Y/٩.���K��a�����]!�F
G}(��X���H��7��ţ�GM�VT�|s��ן?c��@�<#n�'������79��=�[I�LLLnCR�>-Ss.�����M�:p-YqH�Q`��v
�8�b�c�]�JMA�&�쒗��ҮO����p�V{G�b��-[����}��9|b~��#�r22���>p�U����H_�@����MW=�z��,�hZ�kr�+��n\��u�O�8��T*�MV��j?�� �+��)��*vsf����r扬hW����-ggix�s탉B9#�{�i��o|��1���-��LS0d��S� ��|��M���)>>~�g1٨�3�:�E�i>�E?=N�x��?4f�͈��㋓�9lV�G�5�P�~��3���E���_��v����šai���1�1}���P��>ע�-}�4w���R}���L�o��(/�S�����|�~�&����3TS �7Z6�@��()*�m��Oݽrѯ���ԣ�����C&�Ĭ_��*�����/�yzz�N�4C/�7�;b]���^_���l�B>qo��;m���De�w:pv?�Ӣ��[b)�y�oHz?��J���=/�V�W�:ǰıv���5Ԗ�C��a"]���Oވ��Q���{�W����w�fR����xs������b3#I�S˹��r	��F��Y�N��j���h�������gB��eGrֈD722Z,@��~�d�jt*���͑LVB��3�b�Ƃ�;�V��� �;�>���)[�;)�XL��o�Ee힡=��[a�V]�%���|��� /���,(��a���_󅃓�J�S>}�+m/����π��k�G_�e6��:�;}>���F��j��s���G)GYi��N#&6
>��{�<"8Į����15���>Y�WTW�%tQ����﴿oM2�-G}�_�Ʃ)��a:ݯL�%2�k{�7����8�����E����dQXg�K�W05��[c�w���S�^��91z">�/j��}��c}�*�������h\/�����>�i�.C��[f�P٩=��?�Jk
�	z]|r!�^I5.W���Z�k�=xBӱy���Ƃ����'R�������>��\��*piJ=,��1qL�o>͈d\�59�G���/SG��p���E�����RT��-��Ȯ��h�?毠h�<��eA��@f��#�����H��%ޢ&8ufo�ay=���%R� HJ��֧�"1���s�(Z�Ow�m�;�{���c)�>N�EGb�?*M�U����1�������+�sWxcb�&������	sƿ��:�m�V&rؐ(��vi��%G�����*�_���¯��&��Cg�>t5�D�R��;;/Cyeg���|�y��S[I3��}�7�Jک!Q�$�X�d�yi{�-�t�M$���+8�!�8�͎N���9��(&��<�k>��,'/oι��*�������䳝����:~Tj�q���<�cv�(2,QϚ�4�5X��M�wJ$Q���M�ԟ1av	'w0l97�æ��Q�~:S����M�+kn���ʧ�R��.���݀�C������ː݉9���0������B�w�[��c���N�_�I~�G'+�l��\��x�r�Ʋ��q�7��{���v�'<�bD��Au;-d�X�n�����7hv	��|_�DI��!F�*�m���T�g9�Q��/�fH ���\Ԩ�m��?����)�-�RW��(���fF}��%ٮH.�&ek�,rg�Of�Nwб�����m��}xC�gH��CR�i��:Y�f,�#�g�'m9��}�^�^P?�=�y*A0K?�5uys`N��
+����jj�0*~���z�Qޓ/�S5np%�ŋ�wJc���q��΁��:��.�ɭ���ԓ��I��!��n��'��ɯ����e�#�?�hs�M�i	����i|�����7o�ddd����@��u(Kڡ�Evj��Ǻ��m
��v��U���tΑs~h/h!�R�:S:5���;�q(����yn�J)Q������s>D��h��X⏬p~2ğg~�|�Ľ��:��i�||x[GGJ4v��d�|u�'���W�1o��xo���FS��ʬ�,�Ƶ���Ԓؓ7����n~���#���i���R=>�z�q���ki�H�������&��boRu�t�+�Ή�&�Y�{e?�m�*P��e����g�T�-�͛�X�L�G �%�;��4�U��].ڙ��YqyiQUs����ii���R��#AKa�X�m`M�$��럾�1<�l���~�ț��Ҁ�@�侕�G����Bl)�]�����-ڋEńɲMؽ:���n0J������S�7��z�%بp�GO�۵�+�%n�?Lic_t�Y��N�$�'l&72�.WǾ�N��K����zdK98b��7�M����t:A1ث�����'��]���B���#��v�W�p��ˇ���t���5Je's쵼���Uu)�\���!�S�D�i� ;O���$��7^T�j�4g���ϼ_��>C��30�6U7D�˾K[��Ȧ�i���1��*�6^��#���4L-���kl=J%�9�  �4>�Hr�R����_���H����Ew���~��	���O������w!:'��"���L�,���U��ɒ��K �$_W�?A�5A�Y�#W�(����$�S<��M�XT�� *���5�.�8�r,�$�p���(�K^9����WA~++Z2��B���tG�+ڻ�9ө��锫#aW����PS/UZ.�,�h���V������OU���Ay�	�P�m�&D��=%�uuw/E�Wt.[�d;,Z��b��9D�y�������V�=T�m�ŋ�[q0\(iJ*y��D���P�E�f��8_���b�vb#kv�v
�xbfױɭ�j�����B��NY��,�$ߠ�^{�]���	�U}�(���>���C^^ L��x��{M�%��ɑJ3��e%���������x}Z���0�O����d�Sbs�DJ_تʮ<YZJ�@I�ݚ�A���^�L�R�M����E~H�W�
�V4���=�	�I���jI��6�_N�_�=M�'�+��:���̣X	U�����
[ZZ��)���½����� ���
���p��Š�d
��r��u`+�M�-YDGM��[TI��ꢷ�0��{�h	+E�/��3�%&&������Dl�K�4�7�q~��̓%� x��P��4�Ou�b�.�
��R���G�<����cK�=�.\�&�>&@ƴ��e�c�za���U۸��aZ��p�@KFu\�vB���3_�׸�ǹ���^���_"����RN ����·���$Z'yˁ4a�����1޶�C�mBgp9�^������p��҄�p�'��+�/_&�X=I�Eos�t�v�%��
Um*
�𱾾�<N�w�ce�ؙ,�}n:����3꾙���P����>��\�U�-��o/ٽ��[q�a�!��<iQKj���#ݽ�G=XLt9%x��$5�ϭ�e��Mid���B������p�,��Q�2y�.Z���K�;!�傴�s�v�=��t\\�J"L��BVJ��N<6�꧀�ɲ�DP�
OTvqy���U�.�?g����7��fCm	��Y	���O��+S������2xD�w���Ic�=��_�\8,���԰Sk��.N�u`��5�[f��,o��Ud�f�Z��I	� �g�2ݙ��3���]�-�4�gw��u=��]k,f����&���n'�	��� s�K���8u�su�B���#����CCC4r���>0J���c9;=9n$��)X���V���hO��=2�"γ֙�޾Ђ���''��M�C� d��xkb�}�,ࠇ"�P��;��=?m�f 6r��MX�J�DlK��֭[y���{o��'ҰV��vn$�]��B#��(�6 sL�^V9��~�������f_1Ά��H�h�{T�_H���o��� �]�܀z�r�����n!���gJX��Ӛ���o)x3��B�e��E�!m�m��4ՁoC��ˊ�(+���@yE�'��ow��=<e��t����ȵ����t�+\��_<k�M`�x���c0lx4�������	`��=ǿ�����`�y��E�������e*2,|�B)��8��p��a�H�雼>����P�%a��]���J��o���ydX��RW���̍��A�����ν��F1�x7<hL	F�Rz���i�:�p��ҹ�9�pt�x�r�0rq�G�\�#,�,��۫�6��I��n/�z�C�da�;M���-�mSCF�5�N�M
���ےdj>�(/M����c�m��D2�@{�!���[��n����;��2P��T����?;��	�|�ˏ-�U�/�4q�t�S�c�ɧ9��-H��u��Ҽ���Gg�u�ۼB�đGU�<�GV���%����Q�n�By��+�,�,��
Q=���>ӕ��y@����s��^����OU��na�V�~�E�Uʖ}�T�UTL��<�Fn�`6��;hοG�|�à��.���1'`حr�~��߄X�Hĩ��n�M��z:+�7/T��6��q�a�{��#)��DU�AP6 u�.qJ0δf?f=��{EQ�2,v�un�,����������x<ӿd��!��c?&F�7�z�*,U�n`W����vѯ�}��"g7���y��,�����~�MbqQ�����F^�;m� ��������VC�F1�����xE��U{A�D�mh�t]�����V�������0�@TΡÙEX}�mY�J�cX�XA��(f�<$���{�gBdIKޠ%³Xȸ��e`����q�N#��ڎN�PWaV'�c��j�Dӯ
�3�;U�W��66@Ex������z��`��*������`H��%���uV��Ug,�:���~���!B$���e��E7��NN�F�� KX�O5��mG70�j[��4��d��A��F*�t�~�h��޳׉��|t�tl�m���^|�XL��:,fZ��\������6c
J�(�ՙ�x����d�B�ϴ��/9}��DAц�aJiQ?�㭞\�A��{�z(R��<E�ր���"���H>��u||<�����@���D�@w���ė���;:�`��DrQ>����_�����ax�"{X��t��!OW�>�%$���/�+7� ��u�sh�����2LQ ;Q.��o�th!�\�$��yE_ۍ���M'tx+���rh�z���)�M��F1�D@���6�k�f]bIAA�r:)�iT*��7P�����X�wߩ��-�|��P3T�r);u^��~SnQ8[Z�����]lq[H��<����<I��%����*Y��^AUxҗ�'�F��R҈���8��&���7�ܼ��7�%�]�:`�����b~DЅ����E�� Pp1z�[�].7�g��#�����l`���i���.)�l��<MJ���ćXg��������[�C��Y*AA����[����}�,i�Z���{�y��ԗ$L����,��h �6	�(�=|iȥ�F Ф�	�HA�~Ɍ�q��eґ�*u��~�����G���'��UB�>�;�Y	��B߄7��a�wSL����ms@�	<�<�<��-%�a����|J��(�5S��X�����hC�U���+e�z�&�=�*�8�PJ��=#EA7Ja�E�~Z�F�0	��x�����7�,�)���N�� n�<��w!���s���W��uuum�+��JΙ&sn��,b�n}I57�_�w4T[�.���C�,|���_�D�+wz�*��Ȝ��R�4:����W�X�� �/�oP����,�i3j��U�;�Uړ	/�=�+W�Jڱs?N�5Ɩ�Z�W�!��I���mD�Y%��,��f�PGL=%�P�oO$(x���m��ᑜ*���9��:��	su��)m�ſ\��i��L��5���� �,�@ �jO�xiq�+�5�;Ɛ�^�(u� ����-	�������(jh�M�C�!7�V<��I"\�r�������I}��z�v�������}d��cVA���|�(��^jb|��H���T�%D�VqeQt·4�|N_2--�N�d�-�'�$y�pF�ʞ��q�nEI)44�@�3�}�4��6|��ڟ�(�T��D橻�m,�4t�w\W��@�!(���b�\Bݣ�t�6��#�Ԕ�W�a��+�0�wa���\�1~Ok^-�}i������ݡ�O)����bE3�>����=��Tʷ�������l���#�[Щ���r�x���{���"*��+dF�}#b@�Q�'���9)GUBLtb���Γw��c�8�JP�$F%�|���PҞ^'4�;̓F�������~\��T���
����R:�?�ڤ���%>#O2,�殍�v���+O��5?�υyh	/��w�_�[�⡛����Ax���(j�@��lP�[X�;=Ĕ.J�n��P!��v9X�u��W���1dh:Ἔ�g�3�[a�u�	`]��_���4)L��3���l#��/��A�m.ɂٸ�P�ɋ��h$�m|�i�v� �Α_�8���0ZQØz��N�9��1������?�1�TX����g�B<ǌ9�Pͤy%�d:`d���C��g4F֖�]3��/;��|n4��z�׽Y~N�]�/�(9��N9a��ԪƁd\���'����kV���J��z���/�$߶�4��"�m��@w�Kt�C�5����Mt$�=�	�Q�edd,_�������6��Ww��T��y�4�� �%޺�k��ш�m�f3q�b5����0��� KЖ�ہ��=С2��GI�,�l���A�w�igl�����}�#�s�D��N��"�M��.�`=��7��x�
|'��S�^	��VF�(���L-�*��}���r$��dJ%�vz=�����b�LZR5�p.�
���E���$�}�����-��O�a�Y���i�,���gf/{.�{2��<J���������R��Q
m�o6����+rؠ���(R�a-����������|�D��nD!��4��j�|!�\y����$P4�ps�p7Z��)�weee؛Pȅ��N�>f�h��M)�vp��Xi>{?���K�^�X����>�]����'�*�o�n�\�AE���K�9�R9f��~�pbG��gj�ccc�}222;�S��R��7h�pv�W�l�`�z ��=�B��(a�:��u�����͵7	�Sk
37��&�!��0��H��۷�Y�t1J{�W!�����ڨ�D�LU_{;	�z.dv.7�ibB�hZ�͛7!����LE�:���E�J���4�[J��w�����5�pvw���4ɐ~�4�b�k���N0�jJHK�e�j�0O}���e��4t�-)���(�d�m���![���s�e��P�uj�Nk��f��A�\{fwO�����T��Ƙ� ?6�c��G<,?	�2���CA��>����]�QMG����"^��
笠n'��������s�v�kz�j�fbb�s��H}$6�h���]�w^|e*ԙF_&�x�W�?�m~R�x�e���!���)������Wmb�F+���b��a3R��=������썞���L�d�$a��M�5�H�pq�v��LvjB$���Z��+��vTVU�>ݝ��>*�f�F����G�),zZ�ѷy.����AkX)�������|�~1�]���ߜE�#�w�,El�i ��<UX�zr:c��M��=i��2�7��!�顫��6m�������3�vF�m��U��5�
������w�X�>�,��&9��t�z�Ӵ3rg����vBfM0!-��i���&����J;�ƆJ�ƅ��;`VЋ���?	ݙ��6��}G�s�F܏�U\94��Z?K}a:#W+��Pu��b�٧����F���A�	s;����XI"�J�,`+�q�PT�d#42��³�&ub¯�?O)]�a�{�Z.�C��T�{��pl�����4� ��z��/M
���~��
���|�ֻ��� �l�)��]�._�Ltwu�NTr�tr���?+a��o��KVR��bҼ�?�z)eO6���V��Z����൫���� ��&i�If��.��C����f\Ϊv�	-��,X��J��XrD��6_@�:�M4�D�/\J2=�����K�u��s����X�6
�����������@=݄�B+0P:�z�R5�pu��c)�s����ˉ��G�m��~f�Ni�v��#S��T�$�zL�6�� �U�7�dfMMM㚫����T�9��Wz�x2�)��]�����V@��%֢K� �ǀB�
���՝�K�ma�b%�}
&��s�0M朡n��| ��>}�777��V�Aq���&��Ǐ~�Y]�n�6�.����BQM��Ho�N��}	]l�@Y�]]��xY��5`N*�-�����e#�� u��A���`K����4v�K���F��*�����D��˂��g}���x��m��@ꈻ���E:�"�'a��S����$�y�8n���Bk�u��1�դg�?̫��%U�}r*��X�ø��Bu��F1!0*���3~c8c��A��=��>::����/qu��X��y:ő��O���? 09.�����<t�����gyB��G��>u����N��,�*�N���KT�g�3T-�g��������W��L&���=4D�}�.����S���0*�A�O����|Y�W��f�Y�C/s��AVEV]Q޺���-̜>)�J{�#��_'�:�uv�nnI��;�hc�����s�'����� M_Q��6G�����2�-"��S�oa�ܽ�'�xP��[]��@��9��W{��LI���&����b��3	���wї�O���۹O��ߝ�{U�R����:�sϰ �7~m�_��n�X���i&�}Qi��R����XD?���y] �g`q$������8�(�>�u��aŬ��F��+�}R��`̍�0Ѕ6O�����իG��*_T2P�S[0�� ��m����vM��g�N�ڗ�����5K�4���r�k�t���6�z ��_�JY���i�)pM���Bۑ�nV�y��e,O�������,�n#z��Dk,�.*��io��̓�'T ��Z�F\�Α�Y��}A���?��5�g�����G���>&?�/y��{I�nC_K�C���m� ��wyys�����@oqIl%Y��'�I,H�w�9V�∪�O�^����\�}���G���t�0��)(�6`o�Em��Y�f����Nx�����4D���
�!�|��F{/*�[A`��+�#
}&��o8�?Ν��܆v;�ura����j C(�1�K�$�$�UzF�7���HF�0�(5�-�%فn4fz�mR��v����C!A��m����`��+�Ϟp'�Jt��
�d�ީ��?�����6
��l��Qj~�'�'�u�>�9��i7��O~-[X|�:b���Lz����7Bm}�J[uu�#�vB�0`��ގm."<A�����E��^��S=N�ߜ�I�fY�$�h�Vb|������j�q�|D������W�&��7��C���U�xX �m���Z�R�q���ŋs���F �o��@g������͍�>\�D|̳�r�v I���/ҷ��h�V�D&��'�B��:>!��G�|��͓�<Y������$'����5p8_�<�Rˁ*Y�lr���©N����^�wd���(�^NoQ�F�$PR"�ϡ_fwk�D>���{������K2G�D�IT/��sh���4D��H9��+/�JH�����"?��Qz��K�fD�1�u��2�����ӸCLN?��{��l�-\� �UʧqvϞ���# �觷���{R�+��_*x{�D9���DnyL ��Y	�\�Л���ԁI,e"�<}�D�����3�����}�=;ru|az`2.)ieapp�=���V蔿=W7��#}��r��h��&�������m����x!���d�&i��&���L��+-��A�O�-�\d�P�-):_x�J��͗�yw,ŕ111���,��d��]/�_���l�#dfe��(���/\�7w�B�=��8(*�I�5�4v-�F�%���#�w�z�ҿ���C�SP�����Ϧ�U���hsb�az��@%��H��Q��Ѷ�"�Zn*r�-��3���n�L�?-v�
��˟��5ꩃrBF����T�����Ν���ݥ�&�w�z#���^�`��2I �n{����ϧ��3�j��Ͱċ�A��K�ɿ��"wZW���!�>�vӌ��p�힁���������뎔�9Ӗ��n��?
*"�.���Ǐ�f�<�����Sq��8X#|K۔)V|47IK�����"�������ù��I���ߊ���<��5b����}��]O�^��QefɊ�ܦ7��,��=b�.�X}�������ɅYi�٫^�r#��H���	�8�jS�!��+!��`m�ddP�mQ��v���{���%'#��ΌI�b�qJy�����׆�}�D?G��n�hf.qu+�W�3���O�<㪢���aޗI ��ɛAk��Uk�a�n��F�x�r��M����? ��,��Lꫣ �b�}rOL��5Ð�aX\oO�G߂N��"��>Y�/�P ��=޴��CZ���xkp1�D,8U=�FR_��������
k�ۯy���¶ˢ�m,^��R������b�>���cy>�얤�=�\Ǯ�r^u���!�I��<]㟐��A�^���;\B�1���rz_SS�ι�%mܾ�	t{[P���gL.�M9��{_dK9g?K��VZ�`w��T�'�,��Va3�' `���龳�Ȉ������y������2rAW��氉H�ݗ6�L�y�>�|�KDF\삤9�nZά��r�roc3� ⋳�aaa7�a�M���"���ߘ9��,��"�;�)����%-O�hmm-IK�@�~VD���$��R8��d�d���3���勝o���"������dB
 �2w�n�6�]�*��@i���_�~9�>}^B��$on�i� Ž�xqVr��+���s����a����!����W���1V/�R��P��)o��s�\IC:��΄\��9�<@���:)4㱕Q�]��i}}R��.wff��"�,8ωv\>4������,�E�i�R�_�,���f~�a@2@�!jsW�VM��C��b	Zr�ut�A���FJ���C�<��B��
�.����ǫi7�۾y9 o��� Tzc��H���Оu*�_������$f�ȩK� ���?@7��>98�Y�6"|�4���
��zn���2�}��YȰ� �f.d�Οkՠ��vy+�>�+�]l#o�F	�
axh��C�Vs�q<��S�F́�.���杌qF+:v�A�jb��4�A����-Dٴ�i$ͧ�P[�D���������g�ك�7�}���J�W��D���jލ���-vsy!9���B��mSoN�!��|�,�~l��ɋ�XEH���ȇ�牙��Q�ǋpmZr0'''����&�+U2��99����O*����m��� K�۝�o7�x;r �����6��ɽB�/8����C���-\J��S&h��(�4uww����(A�y���t�ģ	����)����u���(�"�5�����2�0�zrкw��ŒL�_(C��x�FB�PK�ܹ�Z�����5Q<���T!!!&ox���T��ȃ���s�{�Gq��l,
S���M(�m���%j�ح���Z�oC�Ȣ��'+[�q��L$T�|D� �§�f?��+�)�S�y��Oz���P��rA��g0k����#����g�t���;@�	r��p����ae�I�*��r���
F[*��\G��Oޑ�(2��~ �~?nY��X�AQՓ�����ŴJ�Ae3��\Csss?xhߐ�2Kz�Ei���H��翧������m� �7�X�n�Þ��YK ?*���#�/��.���$*1��Dn�a�	���!�Y�2Ɨ�hJ���(EZ��夰9ҹd0@���c8� �=�Ʉ_�������L ���<99� � �1�m���S3o [�ڈ��y
)w�i4�;A�����y���E���7hIjc4�����B�����u�>��4��a�7�0�Rے_ul2��
����Ͻr��O0�tv~C]��iL�9�p��d��=� |ҎCn�z����ʯ�Ku{	����3ݗ� ݟ/�XU�B�'���n��� U�p��*�]A{�@ݦ��Β�1ǏW��7,`vl1��m�a���S��������f�<�9]}}"H�KLӟ��%�AD<@��҂�e�S����/��w2�?�>q�l�hmm�U?xpV�`�lA�-�
�>��A�}[��ks��-�%�f^�"[����}|����,�d��db��5���Q�"���9�qh�h>'�����7�l��0�yW�M�8=�ʀ����%��q�prDW�%�c�"GV��n�az^�S>c$$$�c-�V4�??E�����ʊ
����J���c �����!}�⹕O�e��=��J�������P�����Ǚe=��_�~��®M�L��~�������`�}�g�!�2G��5�����{�w@�y9:RLѓ�g1�xaD̛@���M�KHH������4������;�|��ۡ|�vd�y�d\h������.�Ԫk��R<� ��A���([�+�f��0餴����w�n0}���K}��<)����)��ME�����{u~%�0�ߴߡ'�=!��e��U���N@o�A��ӷ�Y��
@z �5�M�� Pe|C7��I���D��YB�gqi��{����?K���_ ��C����?��a���0��`�sD�6���I<��F�d�"�ws�����G��>�X����0:���1�芆��6�j��;"��sc��pG�W]��:I��$����<߼LB�m6S` R 
�yϦu����N~]+��J�C4�bv�]�ߎ
��`4x_���%J�4��r��=�����z�Vj�J��"��ʕ��j7 ��=�!��R�}�'����U��y�pqӨ����4���w�0������+�� 1(en(ʙ[�� L�N����z�u1D���w2��n{��*��C�.��a� #����NrH�i,��>�`�2�P���|5�z����K��ECt%�"���9^а�Q̡�������� �"C�����`5�0�9��I��X=$H�yD뚑h�K�M����X���0@%luu����5��C�$��N��=�ʛYWEs��.<�� f3 r�h%�:"��0d�yu~���̪�_@sh��_*�B�������I�!�ܞ�ۃ�<�V����.�C�#ȗ/]Z���}���蝍�"œ3��I��!�쉾ïE�����m�0�P@1��g���<rd�=��c�p���{��+4��K�ݶ*m�'it� 7P�$z�!����L��x����Ƚ�_ׇD���Wٰ*� aZ�O�VeC��˪&0���Z!9��[J�i]]�\`V`V��iG�z�U�ly'S��>�G��I�(��L~Q�^BQ��K.�r�:���B�����M."k�XzK�'-}�b<5t�{��vUt��d~r[�V#mo�_uQV�AJ�bs� �n� ����9HEY�����m�>7��I��.�X��~r��b�������C�9q=g�Tx�n�[�������W瘚!�$Bڜ=���o�B�R�`!� t��s!��Ͻ �΀��2�'�h	�F�Ɓ�MK�âEi��>ri�i�i��3�J.�y��t,M---E2��8�/ �'����xe�Q�z~�.<�
3J��b��P�4l7��jʊ���_��g�o�v��\}kNT\
�JeT{�rM���/m*�TY�o��s� ��@C�P����bt�5��|LXE�
s�e��o90�&��!�H�.�/�\Ho!Ĝ���J��d�rP�467g�;%W���&�Z�X�b�2߼�{g�^�N8��激��[~�NLL6�;�~��Om�'��0�}�^X1˾�p{CQ�Un����m�D����/��?����}}=������6E�Z�@���*@����8�u����TQE!SȈ�O��Ulz*��͍Oo�ܽi]?>@]��]3RD_��pォ)�=V�����pߗ���)W��gmh�Ԩ]u�1wU{�.��T�J�"�P��N�"�Ko)#��(�.~l`��� � %(F$��j�(���h��ס���������9����d�O*�8�D��O��Q	�c�{�����lyPܨ�oU��[�^�Ԭ,27��,��<�w��.Y�dRhb��(u��"6ɻ�%�\��@���K3 �Z��R��SN��q�+�{$'�.k�
�\^�{y����	���:޷�	H�e�rL;��D��3z���N�����x�6�< ß>�6,n�p�ܞ���3288H�%���;Y���I1��r9d�Cz��}�:p~�\Ԓ�5,��
�Ld�	�0%�R��a���9����R_PN{��_0F��U�U�	�jܗ�&|��z�pܳ8��P/u��_��� <Odj�����'%$�5� ���kU�șq{�&���ͱ)��7\�}�p��I� �h���k���P���? �0�U�����}�re�Fa�[�����Ew��Ukp��y�:��0ԯ=3����	�*c;PY@��&d/b�P�/�*/Z@{�?m�Gϟi�;p^ ����0�7����_���-r�k>��Y�u�Kj�Փ��+@�~����C��WZZV�1٘)���G���谂�b<FCbՋ�fEI���C�:�� JM��	�'���w��ע	oG7�K8 &R��*-Q/������1��A�dNI��A`n�o�I����"�.�G��Q���b&�l�=NM?��������>7�:�Z�����l���.rB�[��Cb�P#���#�؎�w�$Ԑ]�J&y��B�ʔo[�u���2�_�+	�W�����~�CcH"��}
/[F�����3ZW̲hT���c��!	L������Χ�8����R�����t�ӎ;v��1�RD?� �r�Sl�����8��x�9�����tP�M�>B���� ����I̒��5���8�[F��`Β�S ;�ZUy�������r�D�ߩ����:)�NxE]�8�ɃB��ݟD����-�����<f��
�ʚ
�#��&�e�8��#�?=q����&���4H�'m4�)Ed�O�gNG	�>%��ٿ@D����Iּ����Q��d<����v�c���E�c���i���ifY?f�C���9XE6�o�R2�Ѩn�M;��s����Y��� )0���=#��9�ʓ�pcS�h-<HgY_o�FU/�A�4�u��i ��w�O�@�5Q<I�vy��0C�2�H���<�g�XL���ܚ<��p��$��m��t�d��u�6��3(&�]�̑	w����Y����b&_��Peؗ�=�Jo��)--�y�����H�Ul�vh�3;��:`��N�|�g�r*g��T��
Ӿ���L* �8'J�O�8[�B�E��
0�� ���N�P!m����
���W"?��D�0�H5)2���@��f�q��О|�nG�D��������$>ޗa��C�\�b�ъ)��0����~�_dmd���D{��cR��^=�D����#�&�����p�[��Ź�� ?�B�`П�����lϣ����]h3@p# ,�sss�����jS��*p
��v�H�ʂ�S�{J������$�Bg�	��1'g�I�3Ψ�%�78�˖�����f."���A8Zan~�z��z��z��Ja0��m�X��џ��^#���}�%�3�Dw���6	���+��m�=Q�q!�(#�S1�}����>>��d��7��l.}>�諸�њ�&�d6V_!�;�P(Scِ��mݐT�4S3�������t��d�B�܈�#�c~�f瀀 "����@���>3���/-*�z���w�_��۳�c:��mr ��)!�lV�����W���F_%$Y��D-��/���t�gE(������{�7�j���ї��������x����)&�U�����1L?|���Q�Q#�2}��ɞ�UvcO��	���{���Ԃ�{Ԣ�����(]���O9Z��=�ɻ ���W�?�ȉ������6�v�ax>i��Z)xQ���0�,없u��G���|J#�:ט�c:�|�ͦ"Uc���ۨ��}���ڙaSy;m�K"3��|@�0/S�.Ϯ��Y������<�V�뗻�f��	L�0�M������L'OG���I\�B!�VFB��a��@ʛ�f㯎�'�߿_�6��x�x�5�&/OX_ut�?�yXSW�6�>�ѶZ1N`E�`�8�d��`�BFdF� �<���jD�(ATh�Id�bEP�� �2
bd����ɉ�~���w��{�?��pv�^ý���>�lQ�i��$��~�a�H�H�r�j�N��$�9,$�D���ɾř����w׬F+o��G�����[3���4{��{�:v`s�Q$z�������f��#m3��I���Źs(J��KJvμ5��;:�����{�!�
�=�I����M�՚���x��Q����m��h��hkp���a���n �peP?�Z���sYYY�.m;?��T��q��b�����;7�����ώ���vF[�8�����:��$���U�
r�9dM����EF�������{�J��/�r�}s:&6��ь��qX�3r��uK_�h�������5=9Z>L8��Ȭ�cT�Dw2����h��������ӗ�]��ëK������;�����6�L}���mY���v������S�no���ǟ�M2L�An�&
���D��dXv�Pk��б��.-��uK�;���ۓ��[6�Q�qͿ��59��a�"xpNN~zT8	~�)�i��U��>CCL'!��G']'���>F�H������/b��}�	��e�͞�7n,M�i�!���j�	(���:��>X.Y<3��a�Q$��R衼������5:�h�ɥ�w�����9��]{�z"���CC��?�ŋ�#e���n��_� �I��X''��߲*ͷ��M�4�����������zFڡbt��-��ԸH���vf�?r��DRg�_O�k�g�#K��	�5Z��_�6�VuY��]n��w�{]��Gl�EEER)���xzg����5q<`�U�SN��4�dt�;����ӟ��6]+7�
��w�\[� �<�xxF��ٻu�ɓ'��#I��L	щ���!~ꭂ�\;/95T�����O~���37�X�"��4吴�����������"���m�K�������OY�����{/�Ժ�^g?*v��p�xy{��Mpy��7gd#����]�hv.,k(�gӹ��Ш�wlP�������'b�R�A���z,�-mw�1�A�{tt��q��=vd��JIh����X^����Hc��c&�T>�5��tS�鳛�|�'�Z� �����\�G�%4لϤ�!���@�{�����8��;�Ҭ�bC�R�$�����-���m�Z(Zy�<^�% 83~�AG���˹�Qf���_|?��l5^a�� }�oJ,��M�$r �7Z}�;9m9��7]�mX6R���9�b&s�a�o�%PQh5y�[�g�H�UG�&�%�C�k|@Q�P��}�j�������};/o��\���^��rG�g��z���(�9"#�V���Z�Mo�y��<���J�m��I��+��2h�h.��f'<�O�>o/�\J�m�D�I�?W�?Z�R��ۺ��U�!�A�./�K{%B�9��æ��(��BÊ� ��_��c&��v>�-��S�jQ�~z��uѕg�`��7`�������Ѳ%�D�� ]�t5�<��L �Ti�2̵ٍ32[��<�#������$�oqm�'�ϫ�Ҫ�P��bmH͕k8�R�S������]�頻��hY�h���ݔ�h�4��"E��q���Z���4/M��`ck� �ޅ���+w��-���L�9���Pv����?��"��뫆jk�e�k�~�GHww��//6D�%Llv*��ah���T	R��� �2%�������!���Y��[e.��^��|
nG9ѿ�H�_�B��N�-B����JhKS���gF�"�ۗH���ۺ5��z�����(�N=����l�x���䌄,hBY��c�":����j���ڮR�d��u�Qc�?�Єb����c?i]���ѹ�����s�g\���Pդ���9 8WS�9��'T���EE)x�?M��z(w�8�edݒ�HT_��4�A��b�n�����,�Ԗ�R���2 ?�+6$X�!`�C���@Q�:���!���w�(��� ���bQE��S�Uo�����.��u�w�A�/��;�F��62ԼLLb�UI�=j>��>Jrrȝ*�F(��j떟�b�y�4Լ��uQ��1o��5J2x��=��Z���J�-Gx1����L7k��k�������D!R]*�9���T�}��C�^�z�<��5ڻC!mbr��PT+��&���\�j��W��n�dZ�v���ˢ��~�(�E�n/)��yad�*���O.i��GC�TԆ��4�Ri�66wՅZ�,���u��=��ak�6Q���@�//��x�Sߜ���*v+��l���ބ�U�W�r�y2>�����/؂ |�?R��a�O6T*�^{VZ�c@s}����j�,�e�)�SPL��������y�L���E
豐�L ޑ\��[e���l�s(uV��=�Ǯ�,]�D�_��PTO�O�����Fw�B��(�
J���Bd�&����P�B9[[ۛ���A�N' 8X�İJՕU�[G����1�r��6��� ��JPX�j�VDC���@�B�9DX�I&''"w�6K�;wN�Mk���2RT�K�p ���䴹��^ͯE��/_�loȰ41v}��A.�&��$-A��:�읃��ӊw��6M���qAY_6P�O���$l��[#���ޕ���,���}|r����uW�=�yEɶ'ߥNl�8�w��Z�w�3��4=o�_����d�o2ɾ5"�e�a��j�g'�&�wn�l~2�>d΍م#=��#,���l$�ܚ�V�Ҡ�U�� c=�N[�p�Q;;���_`�H�:�MQ|��FG;��+�����L���쌹zu1BO�Ug���m�L�:�3H��Ϡ`��_~izzzl���0�:N]R6x��W^Z�U�����2��<�����Qs�w�����Q�|P�q�{�lJJ��P�l����ڊే��;+���w�����؄�| �=��,|�4A�mv8��~��{4��~�j�R���nn?�>s&a]���7��^��D2D����_0���"����7�L��H��B�s�Zą��9P��'���:���J ej=�q���ڳ+U�8'�������㯡ms��,h>�=6#/oEee����t�t��� ��;Y�����	�)����ޘ����ϟ߮;xJ��H���ciAAAFF5ǩ9���J��g����ʃ�"s�Mq�*pt�CCCȈ�N��W�7b2��+�0����X�9E(G��Oc���X&Ky ���� 7��ۗ�0���A��P�����/P� ���5���D�yc���p櫰j��y�P�)@�]�����A)���T
%�.��447�CU^�b��_�j�-��a=��Z&��
����a�4��sؖ�=0�
i�~Nc�m�
33��:c�GP��s_�j�	1$���������ROf���L�vV\V��3��,ok���b,|�~�h0ǅ����ٖ��j�=�H#*:���w��TKZ��>CU*6"�m��2 #��WSm���jpj�k��� ��&�m����^�EO��˄�1�o�y�ˏeeeG]\�Bo��3L�x�@�����PM���:8;���U�˹�G�BQgQV�lls�ȏ"w͝�񿔶:���}}e	�����B�Ag'v��.4e�%A��V%An�/�� �'&%������B
_q=w���>t�6'On;+�=��wGf����?�t��`����|��/�����f��c���3Щ���w�?�JQ�����oٲ�����Q���~MY-g�p�
�S4;�P2`�S���������>/���%%��Q|���n�"�svV��
��
ԅ�#7 �S�Y5zcc���_<��h��!���d.;s挫��"��B�+#����XQc~��֊p��������h�u�sԽ7��}l�ԍp�546�C��
Z�E�LmEQ\��.������R&��i�� ��+W�B�K��C轍��4
��eF�g\=O�w�ȅ��)��^�q(M��CyCP67���!,��{�"˜�U�6�=�G��]�_�����@X�:4��!6`��Wv���54���'��d�fdli���>�|�9�1#'G266�j�����q�q�"����z�C�r�޾+o蜤bY{�Q��k���i����=������#(���Z&!���|��ڈ�2�J ��xj�ʕ+�����]S�TJ������.\� %-��x%i�v 0����G5gfFK���Eb�ő<0�����I
$�/G�� ^[vɒ%[���P�<S�����ii���$CD	(��e�z
>������i�p����88l<}��Qk�c)SrPWI�Z���2�2����i����K�Z�9��ޖ�u�9%ӎh�*�]x4 @ыe��IT���ǐѡÕ��уy��wzM%���99��2x�5x����"��e�%��*��+��F�x+pY�`�%A���������ֶ��ు#���{F&�	�&��I�?}�P,_�rM]vժpD�P��Q P2.�}�d�UH<�DoDDԍz	�Y�cЮ�x{�v�0��-	��NP���B1���%3��I���nY4/D��[�PB�c`@	K���C��P��"N�-~H1.�+Fz&+͋Ԗ/_�ޔ玲���<�s��i���)���wRS'��ii�tx_�b�����s,c��*�j��x���[�n]���Q����ɧ#���{	�Z��`�rd"�Rh�j���u����|����!Zr����_=��s�2��			��R�ԉ����@4LfѢ�`�%�^*�X�W�J�[����yn?����om���)'��bhz�
Z�1��O�b+O�I��j�h��I�i�B*A�EC#`1��D������zFn�v�4k��g��x8�<���x����zFo�Q���uy������ݻ�'N���׷9~|`�S����Le�0�PD N��X*�A��-��1�Wo �@��E/w��M"���K���

������	���~E�|�_}AQ���!�kc1n�(vxG���d�[W�jkˢ�J�٭����<Ӕ�&�uz�nގ>f�����`���_�A@N���e��**o��P��\K�$mG@f��Z�������1m�O����ً��j�]�^�&��q[��K�-�Qύ�=��Fb���&��ޫ@���+{�����F��1әj���rI!��ޔ�1�������-}�wo�B�=iZ��Wz>?i��]u���T{p��cG(��,SD��z�� zN�`���%p�P�B����a�Yש1�x��o�*c���dZh;C����MN�l�ܹ��nZ.�Mٸw��3c� �y��}���f��+��q`2G�ׅ�$�����>����p����
�������!V�_�xQ�_Z2#��>���1��eY-}4O���YV��u��8�*�n��3��b�^6;�,��XҸ�}u�����L���$����3�OK�q������Z�	SN�Kj��͌:X!�]?���r�-�B��,�<w3fS��{+o�;&�z���P�K��d�;kr��S-�̭�{h�\�K�vKz�Wʡɒ�kb-�nh-�ܹs��ڛT���x�%�D ����k�\��bQ�Eu��ES���:f�৫�����n����#�[��M`��m3���Q��VP#��ɼ����f����8�\ӑH�����@���n��!`b���������4���ETg�R�x�<�{��F�v�?�2�h�U�۸{]���t�����/�t<��,�^3�Y�7�0^���x�k�FV)u'���}ҳE��mv� ���{@Z�t���:��4%�X����Co�@/��B�{,z3f�{���L�NF���>�&��m��]�Zp�������AE�c�����$�x�4�����<�kXE��·C̺}�^�RhnԩK�'uܕ�����l���3��?��(Ċ	�f��u5�	��)��]�:�b������
�&hU���,٘��<�Ӆ~'���b��xF�&���"�fb"�ewo�i���on��'k-[��?.Z.��1�>�:�����q`i�!;v�N}�!����k �86����~{����̺��r*����Afݎ�u���EW�\)Ki!�l|���!J�˜�q���~�;$Kzf2Ug˧��\7׈>�:��^S*����M��j�w��JX��� Y���ؘ��ð?����+�$(���v(��g�+B��z�����_.~���○_.~���○�]�l��<�p_.~�����&ǂ?�ƿ
�W��X!�|xQ�W�/��|���˧/��|���˧/��|���˧/��|���˧/��|���SHCސB�`����ݹz��&��w>^��|�-��Wت��N�Ν�=j�V��),�n)��9�t����[�Q�ϩ]_��8,����_5^��=f�M·֡?�^�ݓ�7�v^��r{���oߢ�?Gӄ�����(�{��z�T���/���R�������������I��'� � U�`ݶ�������~�杰�q3���Ʒ�j��g.�Ő���l[��қ�|��!��C]]y�=<F��7�B����B��/�吪*-��"�������$� %i��6������|��-�I��4G��-=�Iڈ�
wʙ{����.O�r:h��9>M� R,�v7Au!���?�e�#𦯵�翺yY�u����?ۺ˫@Qd�σ3tBΘ�>�����_��i{9�&�9�r�5�\^�Q;Z�h��[��:�">��*��C�^R&!+�f@}�E�9B��ϒ����I4�������?��������:�
݁�E����'Hy]Z�uNQ"HqK�O��W����"%�u�h.k>y�Mj�x���;����3;�7���M��`��{��k�T��!��- ��uujτ/!�C�XdZ�<~�vH�=kw	|��E[|��/��Z<�R����b�H�tCbӝ}��1SwA^?���g�l�ӄ�gE���t�]K���N��ލ�ݻW{�*4�_�������~�������^x5��a��b���K�#��FdL3j����N|�w�p��0���z沃������m��y�{M��~b��9�*El]�g v�	|�׊����\O~�.1��S�ߩ	��|��*M�b�M�ޞ]�0#���g1���?44$q۶���z�q�֭[�%`Q��V��
���G���bQ�
�ñg����1RNJJJZ-ŏp�K����!c�I�8%�ڮ��������Еb�|!��^'ш���>48�c����9$���v�Fm����J��w@S|��������鯲����	FEPq1�3(��7e�`M_�6���}�����}�}���>�z�����LjP��hA����2��{Q`��SRS���K7p���job%^Y*��Ou��Q;����o��W/�W�z���c���G�R��Əa�6]A
]��@���+��Ж'� �d6_b�B��8��%��8v옾���(D���]�Y�`36�M��MॶLd��+��wy=+@֖��������sZ%�.��Q���Y�����?�< kS&�!A1sI��7?����mXPI�~&�N�6���_"�'���W��%d�$b�Ow�2�ד�َV�q�*=��p48*������~s� B�["8Z[LL�X�P�����T�kE�I�XZ��K�]��v,P�i�Xd���jv�M_�M._.)��X�^�2#�4h�#.9��z�*�e�_��0��/��E��i}�T���^#�:�ho�X��o��Q|�l�+,�z�C2�WQ����h�~T�q���®��~�:���]��,�M�{/���e;��,�w>|�LصClW��`�0�"96��S_UD�� N�ӂ������Z!�j8 #d��-��8���?�ˏ?ϼ2w�+Ne�֡��TH��h�`�Ka�cc�5�� ^�6y���嫒�nv�B���<wx��Ŭ��\�������-v�;�z���d�.YH6璂a�&�E$�+��w����rW�q�L��ܷ����h�u��2,,��F�Ɠ�s"���k���֑f�M�Y�#1�~�Yݿ�aI�y��n��z����Qm���7�8��p�ޝ
���!z�$�˖&t8!ҡ�v�BJȷَ�g	�m�F{X�
�������m$���ߞw��7~JJ�$�����V2�uw8C��lֻ8&��b���"��CNt���.fu��YU[{�<��������s{웝F��x�ʑAud:�]�(�:�����s9�S�A��%�1x+��ա�x���'�O��u���Ѻ�+:��.\�c�Ĉ�����K�E�:���"���M�w8	�K����L����#�1BH^FC�`��fvcoK.��3B�ޣ"�$���C��������I�C��t���zp�������zSzvI������!GHQ��*����ڔͰlV��%r��*Q����j̠�#�L�r�e*�1O�1OԢ�5�a�U{d���D�\pNd��C��H�+N��9�Yw����"u��	CJ�ur�ѫ�n��B���.{�'����l�(�V���G�p8J��L����c��dait�v]��?ڧ��� >Ml?y��l����v���-�و>�	�NK���Q3f�>b�C�r�`)м6��1=���	��;����K	o���n#}��ź�:m:m��v8;4z�kK�����%}��>��e':6/�������`�DO�B����-L�R8H��k�86D6�jұQK���<)�� ��n�e��M��^�J�������O~�z�c�Q%h܀��W�S�=C�*ۻ��߈>�	�:�&Կ�Ʀ����w�L����V(�L���̞w'bR�%����]0�ӧO7E[x�J�i�.��}ߜ��[��!�߂c���D�s�%���7u��i����(i�ouy��x�X.(����ˣ5�/;�J&���ry���l�qn"��`���5�'�㝰#��Jƻu~s���{_��z�Y�e�LD9Si����Lv�
���W�%��aH֐$�_\}NCz���߰&������հF���N�@��YE��ty$�ꋲK��
�_Z�����nXD�8���M�t S�}��F/5���i<t���*��Y�?L&�6:F)�|�� ؼ��(�� .�t�K 9剚���Oq&��#��"i0�cD�B	,�%*�~s(^6�����6A�)��m��s�<��	Y�����:���)����q�����v �x:m$��$����6�1��<�A'�_�|��ZK~��i�v��R�\UB4�kI������ۍ	��{Ж��9���gn�sA]��-Mٽ�7	����No^�-0�qƏI�KZ�F��
�ۇ�ޢ��Ĳ۳/O��;�&͝i}��S��3駺k��/�*(�<4���P�Zɹy3L��+���0�޺mυ��9����|��,Nյ��3���i�0����4�Y����w�%M�u�1*R�0�0��Ǣ�޽{���!�$Ϝ��@-��nt��I��؊�FJB<¿�h4�ƭC�5N�k.H������	�������b%��ܸrc&�&�q24��� �
s!9fC�s��*��j;4��i��@�����ʊ\���9*�Y
qt��F��%	CJ���N-]���,YB�S��r&��5���ڗ/_jeܿ?����}2���i��I0��������$���4B�yA[��w��p���':ke�\�޼~�>��.��MB��� ű��w3��R+"j�/�{31���{@ӓ��
\3y%��	}�w��j��h'W��+��PN>z�H�`�-"~���?q�]�����w�z��j�"�d��znTpc�8Z��;��L��+�$;cL��ǯAk���H,I6lG�i�C"&�PW�����]	ۯAF��_wx'�q� ���d��j�B�)�eA�h�tZ�d38��Qq#۱�n���4�i���N2�]�Z�}��'�y<A��C8�0=�.�嫞�Ç���Kn�p��F�Q�6?A������Jr����v�~���@��l%n�TE��Ũ�G$�=(�v�CMM�/� |k�E�}|wӻz�L�gR�S�EV${��1�Nл��r~��K�����_ze��ݗi�,dƍ��l�k�	�ȝ����)��i�?@h��4Ӹ��'y�v��MM��ٙ��S�d	h����c���i]���j�ˉ�������A^NɢԘmD���(���D��EZ����>�����X��8�*�ᑀ��ޕ�[i��\v,���`~�~���.����/Bͅ�cmE�QK��Zl��`r�[��5��g?61*��Ba�Yl� 2��<6�ei_g����V˸~d��H���}drz�;�e���G;��&!�<R�{P�y��<��.ȼ��p���N��{Z�d��R�D�(��z�ѻ�f;��poL��G�+���Aiw��Uvo D�R��2&��!L�S[ѓ��p���J*��ǜyZ����urZ]�n!Z̏�d~!�}3�ۊ6���P�-nVb�H��^�`P���FR������ׯW���!�$"��Y+Jۮ��z�����Bi?�=�3}hk٨c��UG;�1�7�2����C��i,�K�» !��!Ӹ�l��&�V�&���T�"����nU�֊rɾ8'�/���9�p�I�yML�삤�tٍ����X\��]y���C� .//��[8���3�Z �4F�DY�29�˨@��R���~�/�v��B$r�Fj％�c{�]{�5���!��0�ג��Mh�&�D���3SLk� ���F�7�3��P�W������8y;O�������n''m62��Ԟh��=�)�Iu�cED���꯳�
��c	��IS������,�U����f|�v�l�;�XG'r>���F�VT-��Y�Cm�J+`����x�G���Zx��x�Q�AsFz�@���H�}��˞,�Xkd6��D���y�E���*�ԑ�'j���J����&��hn�BJX�.�	0RO��M*���uE�i��P�g�:le=r�u�#�ni'g(�1;ژ�Y�~f	bE×�V455=a����N:�Xi���Y�=��pʐPft0333s,���v")�v��iUU�>�r��.[=~amz��tAἁ��Fe��3
Q�F����Y}�t��3�qsP|���k߲֝����c9��}�iWd�qW܋��>ZDV�g�쪯e�k~B;�+�c���d^V	����G;�ʙY��		_��W���Y`d��M��T��T�����*KX�Q��w�3=m�;���.�޼iS�$��Q��mȝg����p�B���r�8��t�A�I�.[(�1��.�GFp�1�3F�o�o��y�����WL[_<V��ڳ�CJu'ù�8-��"�I���p**&�PP�[@Z݈�d�� ��o�?N�z����{�ky�w\����'jV���L.�xد�=�32S�/d���!�#�]�챀�~�ظߡ��"��!#$���%��g�<������hoIl���������+�&�;tZ`aj�&�*}9��N�N��	Z����	Ov�1�I��7^�k�
�Wډ�h�z�wb���n'�˝��^�tZ\�-�^_%����+��r�$����%�����(����v��/�Z��!X����	�r�Q'�*����ۈ,K��_b���d�]����F����lR?R����1e��7]Y��:4�ot��co%|s����<
C��$��܂ſm��������|������B�8����,徖:�煝����������ӃA�p������D�S|�;�D|eψdapSk��I�ȝ:���:M���c��]qP�����	A(�⸲i�@(��s��L�;���ߦ#2D�zڻD'��M��ˮ�y`��{c�Wճ��z�
���(2%S��Jl{g�kE��O��E�+:<��aKC��U��0�l0y�`��y��p�Dfuͽ���s$O�Z��)}�Ԟ:择�\���i�KǇo��0�hTDB}ϴ��9V�������IE��AD�!K�g�j�@�£�r��$�!����cI�|�#NP.�����~��,^)W���̠%r[�[ᔾyx&x�\�Fx-Ӌ�g"�B�ĊZg��v��/<5O��RT����
g��)؋���N��V��0m3L�?����9��:�k����J��~�t��r3w!@w~%�e��x�]1*H<��bv��9��~�o�����q�1N�] �2ΐ�^p�ҟ%����Uuj(�B�DCI:���wF�=��}ѽ�V�*�;_+������?~��-�D~_��_r��޶�♈ C����ُ�5k/��&#�����C��a3vװ(���އ�^�Ȳ���D����)$�y�N=�c��"��cG\k8k�X�\�&�B��K��Ђg�-��c���r��~�K��J<S�g���:Q��Rsz9C�W��SO�#�N-&`y����OD��X��U����e��C��.�)ii��u��Q�^`��<����a��dB���뙰r(�e�C��h.++C�ύ$��4K�u�L�]��vE�!�4gtr:M��]<�mC���bj�%R�s�����8Y�Z����!6����O��q.6޳<�gb:��l�V�2�Lf?�U�<+�����V�q��w碚Nʐ�6j�Xc�x�� -����;LLG�D�{U89�&g�����c�N4�VTT<$"�Rd땐˼uK{��i�s�����a,�yJ��N(��Qv��2-Ea���j�i"�2r{��T�r�RĢRf��z*�:�1�y�!2d֡)@����U�ȼ;M����\�/�
��R�F��0w�[��U<ގ��33�������*�.��bټ�5?��x}��d�!~��=����ZȐUnР�J@����CD�+6G���n�͗N9V��ޗ�1�$�Y�`�U�8�x����gW�Yb����B��QI��.��F ^7i,3�}�t�!��<-с�}[��J��S��#VM��K��2��a�ݑ#o�ހ
�'�����8��]s�ξ�76�gg���N�|��S��K�O ��o�=W�\魼H�U@���y��~y`���F]�L:l%�2V{�$K}��u���P��N�A���+-�����������i������֒�&v��tP	�@�p�M������ڣ��\v���w�<-�/G�$mO�|(u���>�ܟ��3�6�S����w7"���d��i(���/݋������kll,��ZԊ��U�S��p���T�4EU�?j�� J��ѦNv����֦��Y����WeO�i�k;����k�����(�jPI'>�v� i�gh/��w#z	��=x�,]àaH�V�]���_�������T!δ.GI��"���Lt�!�ۡ��y�9��PBKT�I�xZ�6�Ȋ�k�@���`�`���N��%�cl�����C�VrE�����Q�&9��ۼ�	v�Il���{%��q�nk%G�u�ʪu	����#Tc�\K]�h4&��_I~��/�W�ASAN��v('�����oe��~�
1뢭��e��A�H0�=�z���l.\^�� �t�%����@��� ���[2O֧��y�f���t=9�Ξ��h�RgD�1�i\�p��XȌB6�S�.)��x�tK������GԄ�sO=�/6�-��}�+K�"�ڇ��?p��k���̍ı�����?�̑2��~찑�\OUi����d|����c�S��U5�u�]0Wq��|r�,�7�~b�Lò�E�❮��港G4�TE�n���,���/4��~�Z��sӴ=�?S��V|�i�Y �?8C-($k7r��FFFVJH�\!��� �P"�Ÿ^���ר1�I��j��A'��Y�Q ����Ij��?C3���)m�F|�&q���sO%E�間���W�2���b�s��%5�UCS���1�*����}5�&����D�+�Fw(?�^"=���gտ��4F��5���ҽ�N�9��I��m�|II��2%�O�ٍ�;�޽-�Qi��Oΐ���OU��u�p����=����o�!ghH^kL�r��R�%IXp��<�����!�O�+�X�i��Z70`n��Y�66�&Z�	.B�Y�3����*h��0F������ϱ�7�|�[��6�n�4v�y��b�t����Dʡuy�2l�l�K�a�܇����`��>�G�z��k��3 *��-����wN�($�|L�y0�v|�]S����K��X|dH�a~s�j��kbX�Ӫ����C1abĸ�"�o9��_���V`W�:J,I�>�M�$���ơ,m���Lï4N$���z?L��\�X�gv������� �I�SG��H�|���(�쀪ТV9���X'�Ơ�����5挲��Au�Zr�ZR���yv�Y���[�T\v%�	��&�>�e"��ZQ����XY�(������fS��*n�.�"�Eh^*����(=MWptphҒ^���Z�y�7��^���X��CY�X��0��F�C�dp�j�@
��1�=�%�ɒ����gN9���W�c�cIL洛��	rJ���f���U��4��8|�gA�q";uR��M�}���M���{OU.��%�C����uu�q��=%��t�w	��*ӮZxf�|�V;w)5Mj�\m��s�q�d�~i��7�3��[ڊ�~u�����&�v U�E k��9b�@�}��h�����=*g�'e�=�6�4��@�����2�944�oab��Ig���I��i��z�2�b���L�SNkν{�c0����.e@s�5��$(rr�zL��h_LD���z�%�f(M�Eӝw/�c5	���ށ��ÁTW;P�;j,?��VM"o=ȭ��ق:�s�qTbELH���7y�32S��l�3eC��#J���TG�o��CC\����f��#X���m� ��%%��S{Ʊ��Ȧ�Ä�Ɇ$�����W������t�~�z��xW��%J���(�r�8��*h������ͽ�Dy�nN�t?u�q�T�&�Nk�"�P�����!�1377W��a��������}v]]]9f��H�0��G��VV��:M`����u����#4�8���)��3ќ!o�RY��m2��iP#�ac����N�u;��Y%��krVR�����9Tr��;�n�\#�vYd	�X�&�����d��-�H��p(�!�6	|�k��M�4��-���``���D�(۽�"A(�wi����ɳ��<�J=�����	���Y'S�lo��*������;��-]���Yo���Z2��M�+��Kk{FR�ъx�V�H�JN�ݻ��⭜����)�gD�|�@����"����Q�?�+��뷹\n��~����*�`d�`<����&�kG�\P��
�`#"<��yB���sqm�OE4����2�����2TY�r�Ni�B�w��o�J�?�5OFI<��s�˷�O��.���O�eT��"X�ho"��D�:��"�"f�e���L?�\�����䴨��'!qįh�|�?D[������yvc7Q��O)e��)�%�Kշ���g^�q�)A��%�$(3M���-����y�U/�yZZJJs	��XBcf���T$1Je�{d��ܘ���~6j�#(��]����������qq�°jBdI�6!�k�����qI��X�|�$�j����x���555�׎����R���=ȰV�Iy���N�_t���f�s�\���ڟ��l�7<��貖��Vԏ�	ԣw���c�6�F!W$�m����p��]�&�Wj�C���J�tel��DKօd@-q�����C���"����C���$l�b��r��[���L#X%��r9��U`�}�D����`t���(&��[ԥX2�z�CdA���	��W���)��{3�v[ٝoτ�ƃ���3D�ǜ��[����8"d��Qo_�ײ�ں���~�e_���p��8�p|����z=��[��o��}$f�pU�����Qm\��E�6`�ȠK��:�b�u�P�\��K�1G�\GnFĜ���_M(<}A*ݱ
����U��?������&օ.�By�Du����F���:o���֯�����cx�8�O� �[��P�l��C�z'�^�=QJF�D�넢 ��/���0�1�r*�S��S�����>�и������DF�-V�:F}eY�Xx�{�A���-�6:���j�j�p=��Cw�����(�5�<g�&��~�w��V��#ԟ,��n���$�K�Qȥ���{��z '%�+��zZh�d���m��h��n�Ih`��\mHp�#� ��5�O���K��ވ���,��{����r��E��	���
�!A]�H���FZ�<�o�Y�ΘQ[����y�|.��R_���t4!�Y��y��b}���ȑ7#�V��k.��[�"��r��#��%��)�kG���#bioo���^�.�:OM�7�J��DQ@�!�-j�s��%An�(1RjB��7�����$�mK�����eH�͡��lv��O��j�vF)_6˧���>TF��o�y�5�~����ˠN�;;v,���9"����[N������J�t��Ut�v��`|����N�.	�yė�B	i�'�R����̴��t���D�zW>�~�x�P(lՔZ���%!�]RF S��g�щ�ΐ�<	������H�����'��G1;]�!T���')(v��יh�*�tQ���&_��X�O{����過Y�֕2�?�;��r�djC7P5�5�(ʵ��q��?85O� �-Y��M���)�^���xH13�Ǖ�=��������؆�4nS��b8+g�o9�9�)fh#���%�[���_<��gЍ	)@�9g���)Ą� �õ��YE�갅_��Ox^ I(:
�"H�����=�ë�r퇴[��oJÏLf
�{^�^�r������<�!��Ƙ����j�JR��\1�%�~��gup7�A,b�I��K����s/V��#~�~�&p��E�#��;�i�Ԅ���#��~� �.�>��x�׽�@�y B�ie�I�����T��V��<��z9���A8�w�(6�{�ՄSOY��w%��v�=��ۼ�U�g�n��@[�?Zrܾ�"���`֩C-^+w�g�(��8�_?Frn��	�<v�tK��X:a$X=�k+&�"�����LN���Q0~Vk�/�21����5���w�ʵ+�	�7Cb�Df�Lie���'�!�Rpْ��cפ /L�5�Ί�6}��Q�u�%r���NN��萷�8¿>li9�������"�z�憦��z2��g�(kK�]�*��Y��>���H_��'�uے��#��{��S�jB��*,������c.��j��A���P�7�U��c34�_��j�Dp�u�C����@�\Ǵ���~�"THّ]�K�	G�{�����!*����)��ܽjj,�`oo�	 Zǽ��(ĨR-��»y���"�9��������i��n"�%8e�%��"%%%�qJ�o�_������P̢�~b)�9���"ەl��ty<�_i��va�[hÚ�r����~�U��������z6��y욡�˗�n�1��$� �ju� ���֒�\�.���<Ra#n�#Y#D(�I�_�N�Ԑ�N<��X�M��Rt* �ҕjVۡ�<�N���(�qC�k?K��rqee�5fG�Tr*۝��W���h ��tP�zt��x��)���32L/AA��a�[}��ک�P��@n�Q���X�8�s(y��:� ��B��goQ�đ̪d�N+�	��X����l���x�]�܏��5���@F���')>�=�����y���5�"@0�r�A� X@��i:�]�3������(��0��$�!�A�����J�3���[��~�)(&�&�6
'I�r9��<�evM��Q�����e�/_>���K����.�m��ur�U�K�S�����9�__�?\�5!�,�]�r�X�g6P���Vm�߈S�xo-��t�Vvיڍ��^�����D��jFzZ5���j8�uM
���䜈��@�1
ـQ��2��]:S�I�ѱ��ԓf��j��o"*d�\ ~r��q����j�:�s[1iH�x
>�+Q�/��ȿ��G�{(IM� �*�B6\ܻ9������V�vLN�7�������-��M�=~6�}ͳۄ�E��@����.k�*oB	�Y�,,��>�/�	�쯾3A�h� A���Dm�E'�b/g�Sܙ&=$��z�Y�,�>.j�Fn=��Ҥ\e��"�W�kį$�1��:�����)X��"tN� F��f���ꖢ ��:O��>���Z���X�r����/��^s��]��P��\�#��=�{8�i��{�$�~<�λ��7~��<d��۫O�&����e�O�G�{Q��=�u��v���U�{-��7���3��U(�9N9�v����1�"ף��	*�w��|�w�������0k�..�Y끅�!��n%��n, J"%5UKNN�ƽ4��(3'߽�ʸ����u?�u���~H�/X>���	v��N�ՒPns�'�x�;�@�AM�)�ދ 1&S��(-���,�Ă��A��k?���,��i��hg�RL�SV&�_���r��h��"v����F�y���(��i���:���rDkk`�wtoH�8����Ī���&����l�n&��~h���XD����PUy�	������ce�g��:���I��K�@�(����%�a,E̺�G-������ߠ���g��Lf���F9-Slv����yE����A��3����'�̲9Q�����Ch�_e&qZ��V�z�5��/1�����%Z�����ה�.ҍ;��>��Ri��Ҍ?ˮ1���a����>��z�@�I��T�S�+��zk�v�<yc%��3�������Q}_�mv�Rd�w�[t����5Ǩ��(��J ia�Ĭ�2�J-^�:~Q& N��i����8ik�_�֙u'�.�����5a��w��V�1�aw!{�5Hk�]1s���	�S执��?~����g4�`�L�offf�	�C�q�\�bC	�]K]n&�R\����گ�6�&IJiyw~�oyĪHCZ�M�q���:`��w�O��R<w�U�ps����V�9�������b��ݓ�ĠW�������í7.c/!$g��g�C�4���g��w�m�Lz�5W;w�;9̺D>N*$��׫u����j�X:mz,j��ɗ�a�g���Z�_v��IN�v֦\� ��_�����;��v@ʿϮ��O�d$�NNo�ѯ�B�:�s��ū�.�r�ϻGK�&�f��=(6vin{�C���f��ࣜ��M���{�7��g����������i[_�Z6(����!�5�"�E�@D�@�~�}ĉ#��3XQ@�(q4,Q�FQ��o̍>�R�7��{��{���~,���2�Ӕ����w5�j�
}��D��=�!��H��eR�R==�H�Q�/ef�?���nD����|��_Q���<��!���O����u�Ɖ"��~��:v��Α(v�U���&=��j��,\qL��)�4-qJ���`q�:z�␈��� E�
�Q	a[�l;����*\���A2�ˎ�X��N(���u6m���8��bVֈ;xZw���׏����^���θd���p7,s+�5��'%��8�U%b�8�fr33��!+�Q���[&���1���!D��K����#Ʌ�\�o��a+@[�˵�e�da�.Y	���X�ҟ�`ہ'oWh�-T���*ZNNNk��J��9����,\�Dת�(�>U�Y/r��p��4MF�=�?�|-vlԏ�U��J��!'w�J�w�Ĕc+�%��/)»8ΐ{�J  ^ 
�>F��_l;���O��:@�BZU��w��ۋ�Jm*���Օ6Μ<�t-��LƭǞɻ6�YB����X�
�c5�	>�K)�Tff��8��:��4��z���٣��@�o�lNff�K���k�\|�~���Ɓ�V4{R�MI�߸q��''����0���au�K���@�%*f��C���$��������t1�({����3����>����?�Fg#d	9��F_M2������5{y�o� o^� �ݭ{Fă�'df����V��H��Zs�\���ɠs�XK᛿x�~�w�]�C"�N]�G��-��eӣc�7�r�Y�jH�,�^�?�N�͜����!�`M��~��u����~�����Č�Bg5�3_���݇����W �����๳|w<�qi?���Gw��n&���?K�ea��ZW�L��f�k �O���+�Kܔ���sY��wtc��#�1O R�@�[G0�o��A?(��V�g���.I]t�#���[��E���L��v�&��1pk�k�z��	4��Ix�����O��V//�ALL9�
W��q�;_��U^�+M�������l������[���7�KJ�&��+|ޏ�� ���>��AV��ݹ���CD��_��v����"{ֽ�i��j�b�.z��E,��,?��
J�/���.�u�yw�\�?X��!nT�2���{�8ՃD�������D-ӐW����n��AF*�i)��lȝ�ַ�9����<<�$V:�v�JP�x�-��y���?Rec����u�_�RH�dK.Z����7�!I�H�v�����[����l[�N���]�����>���t���\�="׳�J�mҷ�޽یΠq��v�ƃ�6��c�ݤI{���Y���+�H_�u��g7��3)-���mA�J[Jcq��$Դ�k�g�����}Tԍ��Is�Q�E�^��F�e�>?בF==g9��Az2��p;�m	K�Ŗ��糥�7 �lG!���?�2��3<��`���t~����D9������l���|+��X��+�O��)`M<d��<^,�i][��	�RZ �FOP�̟|||�YWH���n�D�5JT��[!Wc��s�&v�%���gpLS__�J�]
������NG�$� �A�S�b�����u����nz�+j����Z��!�~Q(�|-�`�f�6�7�����~xH-�[Q䠦��چ]q��85[$*�I*@<d7��9#����(1����v�$0��DY��[�f6�p�b!��1��� G�M?/{�RÌ�I�Q�)���H��2���N:R���|��e�&q��n���?y�~}Bqa�Ǐn����z^~8G7B���.h��R�uFo;���f0�;"%�}H��:���E�*�����,f$F��U��7��
�u��@����%�N��O�+:21o2M;��7E�����n��n�g�u��r����v����y8��k���4������C��ʬ�&:�[�"��� y:��>� {�b"��n�]nۑ?3.$O�L�~Ȕ�O��xU^Y�c�G9��ƭ$��6���[�-�7���p��9x �U���
�������]���� "�&w�o�<$�`ڜ�����y�Ђh������
��Syi�K
&R'���Č��G+��L�m&c�-+�|�6���̧�F.=���1`���JP��¦�>I�V�av����&�����o	�U�ڎ�R��_�~��<=�@E4&C��i��p��a�j�u�y/����|>��v����iW� �𫦙�d]]4g1�k�Q�ێ���x���4���t,�~�Dq�F�t#�g���%5l�F�-��ִɊ��;T
�����Eާv^��7�x�+4r�P˔��h݅ǑCX�Dt�i$ܘ�Y�����;��j���;�<���J��1ߙ�25�7��hX�����Q�ω,�c��5��|>���G�:��{Ď�Es!�cSe�O�(�d<�]q��{䄋����.���%K�78>n7�61��qW������u���B��3 :��Ш!o�k^�ΦBfے��q�.d�3�M�M�!���ˤ!��I�L�ސ�~XM[�m2W�2�ʳ�	�O�>�F���I��b#`�
H�W����i�*�ã`��8��3].���M�9���MͰ���
��^��a���{x���.:E�;��%�P3�\l���0�I��m�1z��v��jժA�kw�r>C`p�'Y��d�|I<�������D�L��
�ƀ`0�Fz�Zm�I�+v�)����F�O`��YO�2����t5F>j�F=�P�2���(|��?Ě���6\ugG�ye�i���ш��=��"$�a6����� ��5���oY����#`�|޻p�,�oH�0J�VyG�C��sS{<x��(|�P�]:�;��b[[}6o~v%a��IW�q����O���������酹i!M�bz��L�������۰�g8m���]����
�5z�B��%��H�0����A6B���A �Y��k��r�,^=����Si��◔��q�#c1_joAmU3�'������33[V�ܾc$����)���lm�S��[�m�2g1�Qc'Ǽ��44���D���uq[R�c����Sxu�X��b�e���m@u,�m�����t�a�:�DY2�'p}��Qt.�`��J�l$5����� �;<ǅ���L�&<E�p���).���]1����FF��l��E�Y��v�4���f{���GqNGtR'·Z�`yH�-�s?r�X5�h+o*�	
���5xֺ����&���&3i��?Rv���/�����f*J�Tr$�p�E<$���au�v�t�^D�9�3�q�� �e��[�ϔ[uE~�<��(%����3&f�2�}�mSp�v��w�ܙ���9�ʁ�~E<���kܓe"���^$������^[Ϧ"g+9!�_�Z���e�12��`���z��`����6��Tf��0��A�`��P�1S����mY�z�]�$ FNsS��UHa���f�X�:���j����r4���utԫ1s`_���n5l+X|�j/q��߄���2uȣL�͚�F��0����l������q�]�a�b���&P�'~��E[�wq��	�T`��uUl���ׯ��%���R�D@�ϵ��ۖ�Ӏ�1�7&������F�m�
xS��� 8��V���y�zL$��S�0<��I�Fb�33��Uj��1Te4�(�vj�"���+3��c?�J6��W��Axq��H�Wf��Ԅ��]�.ŝ[��_�-��= ���\M%�kyE�Ak�K�������.���������&��:؝�?Lh)i�;U.�}��Y�����'�n�[�D�rO¤��6���.q��vu2.�-(��H��(��=�g�ʹ@��l���� ��L�tt�6f�'�,�~�p}5b��JJ�����tTB�[=g����Ss���Xﺉ�F�b1�`-	�uu�3���2�Z���|6b��� �=��b^�*&�N��B��<�ሒ7#˵���?�%V��ӳ<��T>l�Z|� Hј�e���kF��(em��8v5/�k͎����(y6
�3#v��D
��^͎�#j�yYYY��P�䐑R��s��
S�Ջ�U�7��[М#YmhO��gΌ�c��e� ���:�NDyY��˦MÅ�ù�\\���m��- 7mA�H�4����Yr�y���K������s
D-f��K��6	C1(5��׮�KblFn�n01�|��(%9je�6�������^%!5����X���D�+�����,ᾤ?���`>K�0�m,�s]T�K8'f��\�tZ�H���Bz�%��[�ʶA�n�c"r�< ��D�%6B��`��S��؂5��E����n�^��~�SQ�5(����ŦBC�?#��s��G�����Tnʗ�J���pu����#[�(4��Ex�]��j�D8�>³�lL�+���"�h�D����|�B�������D�X��P�������9a���n|We�F�da��+��AXm������@��_J���=1��]�[?�g��^���� �}�����.�5��=��y�n���"5ݲ/S!��}��m��kD ��}���DL�D���CeuU���kK���;����19ݥ8�@�-�˒�,�aFM�lCi�s^J��Ơ�{xk������O��<�������~4���.�DY(`s���s�Cm;1ziE{��en  v�-WZ�TZcrB�1-��`\9'��hJ������OR<�ƚ9窐����*Y�pb�E�^�z{�J�궉�u�B�9�,�_��\�}^�q�m#eo�$z�>	6PԷN�@ّ�괤��H��j�:�e�J�$X�)h�E0�8ÒF��u��Q��qZKs�xQ壝��5�WC(/OO�4F66��?{�v���N�nlf�a���1�p�4�X��ȇx����$��ppuՌ�z��H0bl�>�Q�),J���ˏ���'�Ho5Y��Bf���`[���z�mG:��D|�َRݏ0��c� �P�>�*�CL�
㊅�$]^a���t�����()��i?�iN�-��c����?~r�.E�K��� `� �$�ϟE��vA!r�2�l������j��e���^�N�M�kE��ҕ��T�YIW78�'��s]����?�-�;mؐ���E�8O[��>�b��7!�o�ݾV��յps4�cmŞ��H�ZQ5��� |!��[�;
��![�c��6PU~�8��u
�U��S��3�Wc�����x9ZZa���k��������e�����8�ۈ9�o��9��h�Y؇��uA��ӯ\�rvس�Ѹ;㳒�Z������~��ne�"f���þa/�œ�*Fg���N�e��:���;G+�����vV��ʟ~�G&8�=���z+Ȟjh�
�m`P�&ƫ��ܧZ\�{B����X�H���s��I��A2��qS�_�ό>Y�'@;S�ѝ�Gh<0�����T�8a�'ħ^�6J,�c�wx���v��n_'h���K�(�O}���aQ����;��ow@��B�D�b�q�+��P�G�޽����E��UbZ������4�z�  �^ 73�3�#�ع�7|x����F�i�`�zM3ng�eБQ�w9�CbdZ�q����~���~I��PΓ��m1��u9g�5���	��R�B�<ؑ�����H�h7��u�w~E�<�� !���$Ƌ����4���l!��jo��GSccT,{x���)O�PV�$����q��}�p�o��nᎧ�!Ğuqv����Z�����s������+�g��f��ƺ�k3w�R�� .5F�������{�"��nK��d�C���5��ëن��Twf�AᑶQ���X�Wz�Z��w�T��`*o������!�#�p`�q@��7B|����ŋ����X��6��T�Ǉ�ʅ�==�/��I�����	R]d5�~�s�S��*G�,մt��Ml,���]��Rn�i���x޻� �@��(xO�$��xC��?�
��+N>����d�F����lݹ�i,fz5�\���_���DBD�f�]����L��|)''�	�JyS	���C�B�
��|a���O&�4�a$�}��^�IQ'����J��͑�b`��GR�>�
wU����wt��p�X���4v��e5Ht��*?II��7�̶?Pz]���ll"�
h
�1oY lTg�"���95ƹ�<`�@�^;kv��^W�M\��A�3n2z�Q$�?�O�*Z�SF��7��4�֕�Sl�8���_�mt�MCv�~��{m��G4?�}�e�O��opPݤ�C�O�e顇��#�Wv��?��昋��	�_�1QD祪��?���dD�fj��t�~8����|��n��q�>���u��ٔ
L!���AGky�QY�ME�e �����砞�k}��0W{�-��XJ>�n:�<�=�p���O�QB � P��d�\��q ��F�J#[�E��P�y���%ާldz1B�.v,�_T鈎�^ɫ�������ZЋd/!�-%D�����T���;+w��&�Ֆ5�D���έ��Q���0��>�v�Þ楩$ܔ0۞�"N�֜(1E �1�ˇ}}}�A>����0T�,�!�@�v�?6��.�N��%*$�2�
���{�2�@V�;�&|�tP�h5�/k�����Բ,�D��N�z3&��������Y�������B���]$�Ի8�@8�\Z�6Q�>.��ZʴH9����Z醡�� 3z����Ӳ�aT�n��ea�..�,���=d�x�߇�_6�#��y�N�����%�5�`4�����1�j��K�=��;7�B6>^�7U����y]q�8��܆�BP��ۻC��3�!�_-@}2�$�ڥ3���&�ɖwJ5WV����7�c=��K}F�j���o�}[�D�w��7� [�r�n��/B���F���d��f���p8�����= 3�σ�o@�	d�#��Y�%�3���7\��O���u�Oָ���^mn�h���YVh/�_�
T122��ɷ��A�f��{�ғ~��m?Y�����Z��+�I,�U=K$��ϴ@c7h�B6}2�&�q;���>��w�קԓ�XZA�f�ɪ��U�ވ�#�"y%8���ぎ���l;���켼<�j��&1�`�2�oh˫��^�k\�Gf	��0h���#o��vY�u�l��3h����U�����V-`��<�_�~��e/�n7g�[�A�\��í�?�]����Y�A���i�?(q����a�d���֭�Gy�4��ڞW%�"�;D��]!�;�Ʈ؎s[E�s���婜e�Rͱe��QdJ<�����ib�f�L6��P"@����b�a���]�3'OP�� ��G�h�c�t���Q�����q&$�R��`ڌ^;�^���&ʕ�@���S<��u!��?���|5��<���5p)�?K&IT���Av�$����o�H�4%�f<�S�[��9ΚU���@����7{�K�^�Q���}��LZ���^���r$��|v�����i�j���4�s��s~��4<�[��^�7��L�>o�(CUC���9:������0\/%;��Ejj� ���0X����>>>swf�!����կxx/�3�;���P2�zHi��Z^�܌f������˗��ə�A�gO�xդ�m�~L�� gr�4�t;x\K[֠X�s�2 �:900���; 37��v�$�9���S�6�վh��+����� ���ՠ7�������2u�-�ϴ�8��a������\�ja���0�_ET��s�%Kzy���<r����R�UM�{�Ǧ�9U\�Z���D(=��q��w��/��I��!y��#�)������Wo���Uq���٢_9��?PK   ��!Y�1.:�  )  /   images/8d2526ea-6e7a-4b7c-a99b-0902daeefaab.png�yeO�-�Bq����.Z(�����-,V(��Rdqw�Xq�w�E�J��H����yor��͝��I�L2�|��d��5U�	100��0%����?t���	��h�#7��'S��s�A_�?��K��K���������ח��孧���-���}�4��-p%}��c�4s�����ݹ��'N�"Ł�`my�׊��Da_����sY��]��`�~!�6F��	q�8�1"&��^��.=U��>������6�^�>1Z���� �Uw���I��1�vd�6ǐm�O�w�#T�7�<Bħ�O�Y�5��/l�8��)��*�ǥ����K���f�G�Dn,*��:��֘�ݜ���oN�`���쪰� �<)UjJ+��-ݞ=�T嬞o����B����0��p�W�	RC��r��",�¦��e��7���P�A�H�1��y�P,�F(�1}O���6ez�>�uby~���I��ڷ3��j��$<�洀H��%��;ϖ�o�V���$�=�+6��� �0����@s�	h'/?4�M�ίC݌ҕSp�u�~���-���x��귾3kF�&�>9�ڭa#|gTLw�ܟl�5�aI_z�߆f�~[%tQ5 ��:5���FjH��������fQU���Sז���_�8�w�:+ ��/ʦ+n�q��n��<�"��Ԑ~|���:�4�1=�ݡ�/'��^�E��8�t�f�x;;|*��ǌL����������4��?Ż)*�9�/��W���/.}�i�d͜���Ss72�6`I��3�������h������پ��I0�R��)#dg2�w �BP�p�N��	�
2�6�R�h���[��[�@�X��(��
O� ��A�޸�������A�m�	�Pn�*E�'��CC*c۱~1Қ"Y���k
�臨�RyL"W�x�E^��x\o�<>�|�z3 Is��$�[�I����*e�m�ȓX �рH)4oD��d
�X��/"d����h��q��}_W. �4H�$�H��E��k!+�k��~��x*{���Ģ��-���( ��h��(�|��7X]D��L��oۜ"I;ZCo
w���;��-kv�5���ID�Z�'䃨#z��[_IY .����S<_����cO[��u��^D����T�yc'�n��N��Y�C�h�ؓ��T��Ҳ���6-~�|j�������\����4�L��%-Q��ٔ�VZz�6��U�N��%Ď"j��\��!����u��I�l_�Q���w|{V��Ⱥ>��Š�����n3|x|��w��r2,p����m�W��s�I)�C��;���T���p��P�g8=�G�렶d��(��|�T����-��iķ�\�d�/w?Q����6��#O�?���ˈZ����c�\֍P�}0��G��۶Yhol���TC��F�%r'��l֮��o�x_���_����GP{0/�Z��Ӭ|F�L@a�.��s���|�3;�٦9���u�%z2=�9���wD�Z~"u�Nk��1y���5wϠE K�<�zzzB*������+��SR~����	G� �yw<QiG莆�������ʭ4�K�{��u���j��Ѩ�ft����q��42>V��CVo�!n�B�����=��!���_ʕ�c��'6��~��f%�k���&@��R��a�5�e��XDo�{n�̀}�wǐ0d����̓ �P�:������jӊͮ�!�Uu�7�Ќ�^o�S����܀��eI�s��|7%r�TK�������K�du1\a;ֳO!�Fz`E�����ބ-�����Uv�����TƳ.��]ܮؖ��.v�bA��.jM�Ǯ���������.��<���2��{r��""��Y���&1Z����׍���u#��G������o��UE�;�~ʰT^���]2*-�J������h8~�����s��:��~�l�h7�Wg�%�`�	_��U��:A��!3:iZ�^T�)��ʴ8Kw4\-�/��~;��e+��1Z�9\�ap�pb��leaE�]7�@s}t����X���� �Cf献/�[��u��kF��[���i�e�`��aS	mH���F�;ўH,�Q}C>�{��gذ|,��Ŗ�`
9�Ӫ
:P6���%� �84�H4G�b�},V���h�Bg�\[��"���0� �o�פ;*��Qv������p��3w�����J�#�G'Xq�i����"����Y��7]���T��'+8�9�$_V�TN��&�|�g���5�a$3����ܷx�fo`��܉?O�j���n����S��+�^rA�n1�b^��U�"(X�$���5��q1SH�J���Ʉ��$K�Qq/���NG�O0�h:�}y�[�.&j� �+�ma��yr���5��З�(����WF�&x&�4��[@9�ɪ�tmF�	����9�E��~�L��$*���\d�o����齬��߶��9�V��@�V�����'yG'X�R��M;�ˆ���%>/�$�� cv���T>��~�I_��~Z�Pv�޳_g�d�
U�/e�p͇����3�s�c�*Mi�!R�ث�8Y�	�N��YSud���d��y[�l����/XJ�v�)��������ٔϾ�fs��a��$�g��5R�����?V��-p�b����3��z'*�~wWe��F���9����W�B�_ZL A�,R�B��,zֲ]y��^ԺR���Y�z���D�J0I�"CA�����0u�]lC��j�� �Kr^!�������Tڸ�8���ϰ $,S����W�k�ì$*�3��,�0檋�K������j��/��s{�É� �	*̓�[|����nM;����3�+��V��G����<�0��4Z0�:G��Ps�Na�:�`U�z��������,đr@(6cV����N�ئP��l��;SE�6}��F���}[UC���v��Y�?6�j��\8�jabU�3�AD�?/��s#���7N���B�Cr�C)=^� 3.�_����1�c�1�t�I�9�t.�`4��
���M&q5�ޞ^J�Z+��1t��8ii(os#�6�(�g�=ϲ^:��Zc�����O��q
S�����!C�*�]]&mQ���%?"_* C�E��#�
��J!�F�]#�L�-s� A��c�t1s�[vn��qۢ6�.�cڶ���7��~jJ��:z�6�A�?B)�լ��c���n�U��ceII-�t���Y#*������Kuv�:�x�<�S�h/\�C@�Ο��˝��9Z_ز"�o�� �Z��].�9�ɵ�/�W����"jQ-�0�+UOQw��8%�ERV�.EbM�J���b��[�AA�&�Xw���5�C����B{�"����R7���$c�R�13���?.�T hS��e٬H�e���̱�*��Ҥ0�D7��(TC_�K��&b�	����zX����>}C��}$c-Ag�H=gwٰz����4V��MRp��ޞ��B�������lyyb6d�`��I��E�d�K�q]p�d��$��U�H�L���D��� �MY���Z�����*��CN���J�[��5KK&�����Q.4���������Kk��U�t,m^}hg�p���^ϻ���Y�6-�ݓ2:N�i��{QK1�@C=�0z�Az�=�PL!´��G.~�:	@��*�{��r�d��%^)�����������/���Ո|�b�_�n�d�'%�%�|��_m��zKW�#�Cͨ��9����I8d�봍��rS9�ʚ<gX��a��z��+�Q��|�l�,+�����U���ƉP�B�Ix����uX��с桨�y�q)>M6[�d� _q02}����IV1��Z�YzVw�|*������\E9L�%|��&���OI^/���P��'�q�M)y���(o�F�����A�3�^(~n��3��¢�Mbt�Q�0��[{�	��@�8���Յ�^�e��5�>j���^�@iI����w�w͜jG�RB���,���qK�qK��_q3�c�	!=uoGi�,���EA4�kk��=ҢB�}R�e�\�ቀ�]��[b�������)�j���#�&�4.�uu-�!�-�T�2��i&ig��p����������	ҙ?VA�Y��^NcU(x��J��ѱ͏p��ص�sf:��3^~#�=2ܲI?���嬸d��xN,��ΤL@���rl��z� *�Pmq#����__7 ��H�B<j'r���I��m�H�3��\�hxi�[�q�ӗ@[,������%����b]�pvR��Q{��̜�޵뤗_2�)y��ѝ,km�R;D����2]�L��R������n�h�9|X�q��a|i�
�W"|6^p�[�Wȳ�븅�`<kN�Ә���?G5�^l��2O�V��]7	��0��m�:���PY���&�%	'j"��,3cj_Ns���+`qA0


M�z�ax�(�)Ƀ<g�5$�0,�t�<�1ֽ���lj(�`/#�g��}���	,�}���8F�&�b
UQ��!;�b�#b'���dV����@f�(���\���S����#h��O�:ݼ��a�XVR}i�һ\`��\`��D�m�K=���}�ITw5!��	���
~�n`()xz=s�3�.B�f�X�i�k�%P=�Ԋ)�jcɶ@��q>t�M}�K�/xW��Iuk�[90��o�A��dy0*�I
0�Ά���}3�?�O�V�m����|4(�e�OӖ.��-Ɨ�����<��ϱ�#E��x���i`C+�D��+൐��T�������1r �^NI�i&c�u	_����xi~��j�o�t�>�d�S��,%��Xd�z�7i���C�_�{���⢫tA@z�.�S�}4%Ь*,�{�4����Dȩ��L�I���%K��g�%q���w�y�_�c�{qʺ�L0n"/�����zt�/0nGt��d��G�=�x�%;9����=�б����&�}�+�m��s_�l�bV��S��;�r�9�.W�i�����F-;6uoN��I�l��i��~C�"�p8�C�� ��؎�הݮ���%���l���ܕ��1k�:�g����=���{������G͈ne���$�(���^�������q���[�N
���D�h*��(�#Oht�aq�|*�t4E9��mK��(T���]a����8���f'��)��z��������\�t)���'�����`05�t>���Mt�=8mx�U��&��@F�<�)�^|�8� ��w5�j'�=�M�w[�� ���&�⸥��n��Ǧn�!��~a����y�
/����'��ڑ�9dW�����2¾5��.�#�쪩͋�@Um���ZlK`v,�]�#�>�7�1�a�d'�#��F\1�c󱢙�5��i]) ^�8PHN�=�"�D1��ǥ����аf��_3I
�G�$"8�0%����������������[�!���8r�kB/��S5c@B�ND��|�X�2��v,����\�)a�]���d:0N�s����o��\��ʈ��Ҥ�!Iu؆Vs��*X�tq�֗}Ȩ\��a��n�ћ>�Vt�ye����w4�F�)����n��oW��y���V��D�e�(/N�#]`z'�`P��ec�����H�Ħt�����O�]��B:�S����I�a@)5�J�z�@�%��9���Y���\�+���)��M���
J
G��y\�Z1'�Xߌ;���T����yS8����:j�!0-a�H<8���f�$��i+ç�t���!>�A-��\���ϵ�� ;��3��4o�u�Iw9f���f�4"�h�m�$H!{�O�g�c��C�C�)��ঢ�S��"5<���3�o�9���fK�!.�������f�^M�Y���T&۴Js����n�"��B�|�o�[�9l`���2ˏ��WC5���-�Z�C���c�zo���=^t$�[&ˑ䨤}�JzgM집D珦=o�M�[N��p��2�u�kx���ڌ�Ȱ��y�+��.�T2-�SJt�-�k��]��.��0zX�h
��ڒs�%�E��>�e��;��ã�/fMۅ�]j$8� LA����F�TM	��{|��EWՅӀ��"�õ���y$6 N��jC�^�&^k�DL�Л鴯SD�i�yr�,?PC�b�^����N�y�P�tm���� w�~�/q㵏���&����Uq�б%@������� �U;��?oT�-�S��4�j����JX�/���yH��v��Iĥڰd}f�kه[�[eo~i6�y+[�2�Pw�2Md��7"a	L�I!$����GNqZ�m�8qI{���;Y��l]�u���������Yʖ+��_��y
�.�h��f7z�\U���}�S"�y,�fP�Q9���5XeYL��?�.�������]���+�Z��9�j���,�S��~���:�=��������t��P����E����@tuX{V8z?Ѕr���k����7����+9�����뢓oC��f,�QM����E�-��M}��r��$����:�v˝�G�4�]Bp)���q��-�o>�����*֏���ץ�R��-�rc\'���F<�"������\t �$m��@p$���]-8�	Ǜ�&����u56CӐ�Q�� o��j�}||}Lk�ů�H˓��W緽 �.z���l�p��drB�1-E�� �G���v#q�߆�[��׿_A����h@f {,��ӤB�0�B�+9@���ȉ����2%]<�Ǜ�9����ɤ�޻��
"+�s5��I���N�t�{+HI�~���Vr��� �D��v<;�n��S<�x�4�at(�B!�n�#��J;�������>�Z˔z���L���:s�	����8���8<4 /���q���>�5���^�P�1�C0˓��2o�y�����o�Q�,VfϞ�իwCR�{�ϐʃo��*�� N�Z�+'M.��mݏr�)����(u`�{�e�M��9|����/GD=/���BJ9��.���{�f���������(��5a�vx�&�V��<䒛4���I��6�K��e�/j�k�Z�s�2+u^�����Xf˻��{k���s��ZY|u�F z}R#��O�:�S_�E�����ho�lW�;�T:��z�K��і.� ����mjr�b��lT:�˒�:T����Q?�y_��_C���]�3�^�I��.�$t��@��K|>��+�%�;&`�1�έ��9�s�@�TN�_&C~ͪp�Z����
HwTS��L�Pq�0;m�i�4�w{,X��+�� ��$�uԡ��ۧ�~{�Y>	#E;�D�YUq�.%�[��E��S�V���R��n
��O��:t�m�D�6TѪh���lF�J�ُڇ��Ev󧟿�
���/�������\N��#�_ J�Za���/�J�κ��Ȕ��w�QI��dˢ������j�%a�dP&���GW��W5v����n$h'Z�r��Q����R�.W?�MW� �Y󜖱���A��S�_��%=x *;��f�eA��y��#&�}�>`�k<+�z&�x���AC2٩���}ŽQ}ָ`��{�T���+�:�Q���}+e��T?P���L�"t��	����-T���hf�[KzGd��Rʦ��7�Ü?��	dX`M�-V]z�#��k�����5�>C-C�PK   ��!Yu��|  w  /   images/907fdf8d-ea69-4713-a731-45c9eedceef3.pngw��PNG

   IHDR   d   !   /w�   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  IDATx��[w|TU�?o�M��$��J*(ME��O,�*��#,�ڐ�YvY���������]WD�JBI!e�&����ι���˄��o���03�w�-����ᡗ���-��֔Z>l��91E� =�������'^����O�[����6��-�7��iy�r���;��{�?dK�~��h�9��P0 �Gw@0��S� �/KC�z1��y,� �U<������|�@ P���^q���[�Z[L&-�k΀-9��qr��z�J�C8�)�	I�P�Aj|�R�ibz���Զ����u���{+������<8�1諼��E�ڲ���d��}����y(�Gá p*�p��).%%Rl)l\4a�<u��Lf���`�e�Є�8����T*��ׁ?�~y�������N(,(d�e����-v(B\��D���N�;[��
@�Ӊ8.�.W��ղ��<����_P�U󛚛6z<�u�V�q-�����]��k�����Ld�p:�u�\]��z�iPzV����4�V����A��ʶ��ۜ���s���^~���S������KHa��STy�פe��$aGV[�[�Z��1X~&j�I�j~�	�T��!����۠>z��g<�����P�9&�ZZD�0�ސ������l�����px���z`��M��q��j�9"�Sq^wT�1{����hR��]_1b̍�Z�)ZbbN���>����=s+
�=����hjl�J���F6����M��k冔����U�1�V(=��@�V"��S���
�b��HOg�B�x�����J<�j����8���"�o��H+���{�$Ԣ�"-�dԶɟnyo'~_�����Du�+))�o���5�v{��&������h��W�^��+��f��_[���l� 33sK��3g�Ogk������Ewt�5;�֑�����M[�,ɖ�z� �ʳg�b���St���F��	��+��v�2qUv��G[{�!&��)r��t �HKM���uv:Oe�ɸ��Ŷ�!q^����/�)JIIeZ*�@So����	c���=��T�
h=��a��~¡P'6,,\0��J`�̧�~:p�ۣW(5#�̚��Qa��[��eV��N�(�(��h���A�"я�����i��l�Yyd�-3���n��w�3F����	~���@�]]��p0�x�����ْ#&���y�o!��D�L�ߏ���B��	����h$������)L�j���+�|@�}�ʗ����I��k�T�!��ن��Y1�l�m.��N~�`s����ьu�
"�"��dQ��Ғ����.d���D�-/7�G�E�f�g@FZzD2NJNJ�8z���������I�|Py��B�O��f3�c���1lxU�Af��O�.����W��PW�+��»g/~>95+'Zd'��j	A�1u�*$O��'E?ؗ bF���Q��b�R6�8է�]�	��j4181���<�ЕER1#C�^qj'��S���5ZV5l���ZS}��G�KK�5l|����C$�ed@S��Б�;y�.��ay��Xl�}�v��|I� Р3u��� 2u�/3\AЁ7���1�=~��2 +33�4�����}�s�֒��f�#��!���YP�?R����vtt@ـ�L肄�/jhl`81Y����T�:s��CfH�;8�c�_R
f�9�w�\Pu�ʏQ��8���g��ׇ��5b$lڲg�G��Q���<'�����$7�I��P�Q� ������|0,[�δ����V�ڤS�:�G���F���W1���<A���r��h0�D/Tr��1?����nVF&=!�,��E	����,Y0``�/
��t)�P��H[�S�E�,$7b��/�3Q2���Q6���_Rr�r������.�]E��"��l���G��R5���UA=��E}�h��l�:C��xX��Z6��V�p0A�H��N47`f�B 8�Y�3�d���eWWg��{���X��t�d��A��#8��V��͎�SN&�oii��!k���ڪ�9��F�l�1R<��;h�j~u����Q�ZHc������}�?�c�!,�S)|�t�6˫�~��j+��d��7~*+��:�&Z��I���3p�����\>l֪�3T8�X ��9D���������wN�^Y���Z�{\_��X�<&b$F�xj�
}�c�=�k}�j+r!�d���~ic��<�T`n�>��w�փ0q��A�bL��r�Dlk�q�O$�s����G1�w���)�#f!��t�ԏKN�����;���a>���<�m��	�
�u���)(�7dD(�,���|~Nc{�Z�v�CDӓ�3��n}K�FiAAl0�f+-Q+?~���~�	B���`�額C����׽[g�3�Y'f��7���	�B*d���{��B{��溑Y'[��Rk�}�JG_'�'$JQf��������n�}}�]�͇;����p0�(
�9:�_=qFUq�^~e)<�x���Z��{�h~=ht�j20�@G�Q��fC�pV%@���'��L��5	,�zB�8;)�ɢ����[�O��ô�π�P��6~f��dY�*���w����j���44���n&�3��!�qT�s����:�"M1��@�](���t��`�%��/��VDf��XHC��F��W�F��|�Ø	sL+d�M>B}��r�`���!�f���d���^��0�K�����,�ȡ��B-<�[(aS���ه'Uw�Q8�Rw� ��Z({Թ`�yh�br��������rss!��f�)�v�A�^eK��8v�p�u�\:�.��!%�=��V��]��0�0�0�KC����Ē=��L �s�+�E�F�����A�p������W�i^Bb��};�\Z��q���o~�ƍ���Y��Y��!Fu�`(yʠsI����&;46z��.��=`/�zh�zDL�:�Bmp�a{���"��l�����:wv�cIL(4r�[//�q�]�+��?� �>�+.���F�z!2ّ
=��!^��m	^�&�X�]����H2��(��.F"�l��`'u��6����l��`KI�vW��Oa8��匛���[kNV̛���=���t�}��.}�݋J�L}I��y!�9���]C4g�/
B�Ҏ�Zq��w)�wbcZp���`3�ym��{����J+��n{�Y������"r%�e_b�Xw�����SgG�'<���
�/��E/�Uc���h8����Sz>�p����3}��X]�à��Ҙ��J�gGb�d�*����Y���!���2�H���vu8K�̛����0;@3��\�#�c0!+����v����V�@��B�3a/�Y�@�`V#�R×�	���Q�䷊
�4��$����k�!����1n7|���Zy<@N)�|Ή{xϳT��\��6Ims� q-���1H�(L�Ổ*\+�w�%�΀oBڌ���7��Im���HB�+~����d�@������`�����y�Fge�!���(�d�z���v{3\3�:����s�D�R����3	j�>� 	��V�KH_�0�ʸ�m����=��PT&�`��e\�Ug ݉�RҦ,m�/EڊT��h�7� "&K8	v�1��Dm�Q(;��Im�v��^�C�x�<�����0Ԃ���Ǫ��_}����J�F>����
Nu�\]|���]?|����¼3�`/f+����Ӽk��r��ڦxL������-s�B�H�ь)W��H�t)�ב��$Z�	�S�
�;	?�h�w	�i��~ҀA2g���5 �3NG�o��O'��5;��.�5�����f=��@jf^��8�w6������s���ѻ=ڂ�xv-�ϙ:�1�NWn*:&�1��x8MRq͑�E=/Q�ڡU�'��6eS�� ��������@\D���E�C�Nb�3�s�A��r|p�_���PR6��J���ԝ9�5%=gzte��n��%��6bf��1���G�46s��ɧ��
ǩB�lO8��}�s%Ҳ��d�	�I�I�%i��
�-$�q�'C~�Pm�\f#-B"��B�iN�p~�gHc�#Bln��n���.	��#�7����#A�R' �9TI������_|͘&��N��w���מ<����_���U����=�h��p���×edPŽ$��U��gX���rO�V���q�xb+�"���$T��ʨ��H~�C�W -G:�����hj�Y�~��I��?ܷ@!`MJ�ᦏf^z夵��˯����	�.��:1_7몷�����'��HG����b�317���ӕN�%!��5������6���L�<{ET�yE��Ԭ���fB����s��]�m���}�w��H��H�W!='A<�[v^���� n���Y -�����G��.�b��=c<�Ο�g]4ꚙ�K��^(���[�}tҝ����C	d[K<�`q��|i	��^���)�W��dҿ~ܱ6��|�F���3���衄���e����-Q͐/xMb��.���+�0:�Β>#�D��4���%�߀t/�} �}	"�� �o�q2M�tџ TK�^��� ��R}��H�cI�e�¥�<��`��͖��`p��R4����U��]2�w��!�����m}.�q������d�������PZ�
��L�Z�G�T����P-Ze��t�	��T�4�9�B+67N���@JԢvh�<��4
�P���M.��r#5F$�˂�F*�-�`��.�u_��ȟWC���f���Z��ՠ�꠪b�y��͙�0��� ���2�;��G?����̜�'tzc�t�]��p���tM3�hG
���A͕>��_�ObNt����[��o!��V�@t�$��q�n�ɮ���AsA�F�%����A\���<    IEND�B`�PK   ��!Y�Ƚ׌  �  /   images/9185dcb2-65ea-4de0-8d42-42cedb1b5634.png�x��PNG

   IHDR   d   -   X���   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  IDATx��\�o��ݙ�����uڗ��!Q�Bp�D"��h(U�$B�F_���?�C�JM�!-�А�J�(�U(I��E�|�^$k�w��u{�ݝ���?���gM|}?~3���眹3'֎_�A`$�M!p�8	Q����~��Ql18���gv`��ű�K�Vr���x�p�z�3���rW�y�4�0Ɲ��t��=�r�Ҙ�xq�!4q]&��:׸:/s����Թn�?V̕%�p���:�+3xg�X�@?��Ⱥ�qO�W�t�G�����X�ѳo���Ij��;m�I�Ae�ŰĠaä���	.���'�eV�	C	��h�*��2�z�=.�q�k��I�%WZ�A�KD����rB����'H)��8�{?J����>�9���v�4�'���~��.��7�'`��9F+ o	�'�!p��/e��!i{?�CP����Ij�Ҹ<즺aj;C}��Ǘsݥ��N\₱�ߧ�$ސK�\��G��	y��s���׸��s��%\�I��,� ^�cg���CT���;s���/��e����2f�f�}x;����Q���r�����2	��b�\͘�#���-��pb�w��u6�S��;92���&�}�5L|�,�a��ʚ�K��D1p�eM�H��ugDq�ߣ�[5.W�z�D
!����	q��MB\s%��Zs9ߦ{�/�$��b	ӓ9����M%wk|ao��3�=�)㭱�I��4Me����K�_�%?�q�<��5'��-����Ү_���W��:�of?�˸S@�w�ۻ��~Ϋ�1\��K�
�^=e4��"������W]�r�\�ո�k��書��հÛ�����$����ǰS6�}�������>��ذ�)���Ty�"��])����ZMtXT^��s�V>�q�<C%C�u�2�~󘫕���M5�;s���R^����D����}�s_!�.I��VH����k!�){a���2��0ڔ[���̵��`@��XxL�zp�f�S�7B��"s���q�<σ���ҿ�P��J��h��Ȝ���g.����U�^}Qx��t:��C�Z%�d)�jдЛ�s�1�J!�H F����R�����Ӓ뺈q��U!�M�#���c��"(�Bt��]R*��V }�����H'��t��Q!���xUH~&a�����!١;غ5 CG�4�O4䏱z��אi4)D�Ζ)�L�8:$�U�vQ������:�Gx��x�.��~���n#���q�EA/W�W�H��s��������/�]]T<���}t��.��j�G�E��WX�_�|BE�
���Y�0��/-S���F�]̓����@�1����n���~k��j�ل�C�ޠهđ��CW�c�+��+���\�B��T����8���u<6:.��aYC[q��Z]C�r��X	�z�Z�Z!�Fcr=�/��Ut���q�@�\Ѱ���\�d�\���r�r>jp������!�=w��B��B����`t{c��	��겻�GA��lZ��v}�m��_�Z��v�qb����/�^�B(JKO���'a��iw4���������~zHي+ڮ���E�S>��W󉞻�S*;e�d��vr�-�+�hVXG���f䫊u�S�#�J��Uj�pc��mw|}���l� i�!�x_~=����oܺ*�5��S������q�8N��\����MW;t}c844��'G5���!����}yB����a9F{(?"�_�$9�c�3TC!���
)|�B�O����ؗ��0�W&�RxT�R����s%v�iѥ)��	^�U��=+���0-zJ(���/����R	o|�6��}� �3n�����=zw�G�X�ξ���z0;���<w����4^y� Ο��R�¬����i�C�8��y,U�0��UI�c��W�1��u�Q��\�����p�{`�OO�0Br��V�u�0���\�=�r�9=�Va2^��ͅ	!�sZ4+���w�n������ة�jep��!b�~?�7�՟�{PiѤ ��?�(�*��    IEND�B`�PK   ��!Y�� �f  y�  /   images/96fabd4d-0b16-452b-94e2-688cfcbce531.png�	TSW�6~q�i�2*VA �Z*((�'A�0I�PQڊ"��"2�A@D �A���9�s����������f-���s��g�g?���^��ݕ˄�A����F�<�-Y�X�����_>~K��/u��A�����������t;�d��y�����)k�h�>s������mĀ�0m�j�;��k�w27���$[&f���tt��,�ｦ���ݒ�_n�1�`�=��k-]|�!so�O�~oy����B?I��l���K=�w4��؉#�[^����c�}}҂#n%�@�'�M}S�L�d;vg�|\������zƺ�WOڪ��g����VW	@*<�6++KK.��6��{��4紧���;�쇿V=漘5��L������9/U�c��r��;]�[�Ťk)�zj�]i�19I��DU �ƻ�{
!�w(;\Q4�_v��ͪ6��![�V���1���|�;����0�j�t߮9=X0�B.���L�0�C
�17��p�d��ۉ�� �n�=]>�����A�oVtɻ����1�Nj���v�.&F�3T�gČ�iL��S\\|����7=5��SK�����,�2���؟=���/ʖ��k�޻c�ׯX�p�@|TozƬ�N�Q�TcIx��z��j��xd5���:ﭛ�_��cz����5��V���D�Va	-$���E!����Z�����n�\6�^{�-��0~��ߺ*y�MJ��_����s�r���0�Y&Q�wNउLL��V8���@�%]�A�?���z"᫇�\|G�*�ς]��q�����"�"&"/��M>&n{T�=���j;��{#�-���~~~�ѕ��Fd�UD_��a7�rQ�2�ۇ��.M�H��-��y29�H�Wwg!�
��YW� �ѕ�=�QV$_?�l�m��7s���H/ds{W�z���]��Z�w H'z�S%\���4����_$����Lz켣���y����a����vD��WU���u���#0�O�qb�П9���!�������@!����^�}�{�1�sN<rĂbH���Y\n_��e}�NM�*l�1׀w95�����k�;ga�<T#�B_��zu��X���|MPb�[{��O�%ot������$�u�B������)ڛ:�F.P�9����3�4���s���,�D��Y�!I����I���0\��4�����2ښF0�K=83�jLӐ�OV{�;T&���{6��mr���n�9��2�fq'.�ZҜ=�l䣪��5��9/���ԙ�6���y*�w��,+%UF�lr�M2�]y��]4Y�)ˬ�ޅJά�)N9]��� SD�,���.����^��<7��]����))t7����|���e���\I⤌�p�+�4�m�!cE�Tc�ۧ��O�����`���4��BO\9
����NHk��<.Cȝ�#i*�y�YMMMK�,9H�l~}.]�c�����86VY�Q�榆�,���\�Ǉ:$bBU�Y��A�C*�dz�gHp�x��)q�8�;[� 󰱝��l�W����\l�G�.��+wI�l}��v�;��a
�Ӎ�Y�wVA�x�˾�h��&���@{@����ւ񕒜9KF
�-�:�U��]�V�ç�2�ko�sn��z�ah��d)����
��mN��e'*�[�rFXOX6�[�D�ħ�!L�iG����I�P�qT�G�}}���{o0�N��s�x"����Y�f���]�<�RdX��~��cz�Q�t9�H-tRv�H�N��=cn�a�f��fk���[��?��B�eΉ N�]{��&D������!]��Z�=q��o��e�~�8'Os�{'������r2�p;�CD�zݽ'i������܁�---�=���>�|� �"��5�͎�7B�=[��_�K��΋7�d������f=N��s�����0-]K�S\sXˁP\uz�����UЉ���4Y���xM=�yp�A�s	-b��wn�ϻ^n�34W�pc��Y2rEA�.��`�{C^���;UaG6hsl��)h�(�Є��G7U���d]266樫m��ކ������=6z������-�Xw�a�z�Rt7� �$�](�B���-��s�G8��YhU�� p��r��v!(e21���R0��~��z��F���VnYM����љ9�tM6{�9��iͿ��*�&#A�o�g}�Ɲ�q#6VL�┘ds_��$J`����y:o `��/wti1c��?r��m'^$m #����K Q;����ֱ{��1;J�uC0�0�{��v��h'a��a̧QJSp��W���=���{ ������q��"-�l6ȗ�2  H��f9V���
�K�ȋ@�h�
 �d�W.��5r3�{k�Ó�p'u_�"\��F�V��F�nz���CF�����}zvNMu��x4��<�5b����Ҩ�,ض,���R��˗/�2^��o�a)�\�X烠,��O�\	�����*�W��KJ���a'��d����H�4�%�U�Y_��DgK�TlB�m��E���iÅ]�Hٶ�h]�� �T/^$R� �d����X��\����^9ɪu�uM9�![%� a���M0fJ�3�:a�f��A�8,d��h&���X���dե�fҔ#ybvz V)��R!;����2G��[�'0B#Y4͛s��ϺC��@��l����N�.���� A�b��(��g�H����\U�r��ٺhONl�Y����K:�
��g��ӱ��X��G�Qn�Q���Vu�ƾ��0�CzL$�%�j�M��tG:��|�2g��_�����~z����' ���p�R��X%V7D|f��fx@^�
Ev�9�jN1���v�Td紊(pO�#���sl�T��c5��B���Uy(��&�)S��&�\�$Mw�s�zn>�	ZjêkG)��=]��wX��JQǖ��������nE�?@j�����}sa�
?ᘗ�i"H��	T7o��+�6����(g�׶s%[����圀����DS��Z��\���y(Nz�DO1hXaD�J8�\�����;w��������,É��6W�i�����e���|�>�@�	��6��M���WC9ɵ�o�3L�@a,,͠D}*I}��4c�r7Ǖ��cNZAn�Ct�ׯ��}��u��9i��
�R�B���qW����Y|��i�κ"��ۦ �]p�o��	HJ�;=ҳ��8��1�*Q�t������p��q�^9ȕ�6]����Ɯֺ�'�1tqV���"(}��H��l�0��h�0�5.�RO�_#�#��gPrgpH�f�z��`��زT�c�T��$1.��Y�( �(�t+AzvI���)?�hD|I��Q( �
++��9G��G�g[F+~����&�К��f��1���g0���G�D�t�jDG�����E0��p�S�}�]��-oQ��=BPbӥ$]�n����E�x�E�.�R?�Y�CN��k��l	
X�É" �XM6�����q&;�Z�`�������D�~w	4��<q���J�����uϩ2!���E�5��(�8vu_�q�qL��5���V-; �+
��cb��03�E��w@ˇ���1�̠�&5og�;8��9��=�N�Q��(�q������H��9 �)��|����ŵ�#r��Ǉ�z���s;�EͿ��-�PN[���Q�۶�:xF9Ҁ�
��D�x<ݲlf�9�W ��xމ��=)�<ǀU�_p"��0T8foZ����Ć8�' �U����3�ј]s" /|ŵ���6��i��F�Y�h�֊���n7a9������l����52�X����zw�0�T� ��ӳ���K`���/9����
�N����
/ւ]q~�4�ڠ���I��R�zU�R�%>�`K�e��@%UI����_������FI#��o[�z#9oҽ��w4h5�o,$�K��úW3=^0��b��'��պ9��՛���'��A��[8�����֒P���\��
q:*��WO�����5�Hl+К���<u��l@vyV��B�(��A)�ưi6���WC�����6)^�� <�]�T��:�E�y�K��DϬ�ǽ��5��;��_�ѳ��)�N�Ɗ�`�p�Ig�(y�n ����|+v�S��J U��)�q���g�H��} `��\n��;�C�<�����Xxt���,1��;eJ,��-����ӢI���^�%ڍ�j�oŵ0�mn�$�ܩ��(����wS��QʨfĘ%uf�t�a�ujR2�H�tz�W9*3XSQZ9�7A��W�1!�?#����Z=� T��'_���vd6��`����Y1��y'��;�'C����r�[΂̉FrD�:�(дTm�ZUcBgᓽtV��%�Ŗ���m�����55����mQ2�����sYuM���~B+�u?���=��}"xl�7i�#������I<=��.)�{�z'�[Us@��a�q�Ғ��Y[Q����I3Rr��D�O�ƺ�61�LZ�<|E�Z�C���2������<F�`���F��֚��N5خ&�^�w�	U���:��٠�Żkw�ZE�\�ʐ��w�����)}�	�j)��Vs�ۊ��X�ЗFRfӱ�3-���{�zb���Zw��=���͠���(:�w��v��qqX�M��|���-;������K��֖K��I��YV� Zi�q����c�|0q�l������Uº����4@�5D8�i�����6纜�B����pŮ�D�שr����錩�<�B�Qf1t���Hm�޴j�e� XUL�b�'\X}��O�
L����i��olA��(�2�~$Bc)�-�9#P�����{3��r�t��mS�#������Ps���D�΂��h6���ޓ��y��Zzv/�(��^Lb�^����0؝F�Q5�3�r�ӏY�)��S_���ꝰ�m�sCcb>`:^�Lc�b�7:ekK���=Un#/�
�zk<\Yv(F����X!�{J�����zW ��t�s����\ˎPF�/�&�(�&Oh�w��a�<��6��B�1/�'��ş	�~�rl]���0�����oA/i8��lz�E%na^T���dd
Ut^q(���M�����-�̸Q:bA	z�[C���;D��89�0�zq�!�4g��gf|uw�4�4$��.�I 4�?;[�Y��[8���9S�'�BHjH����b�pؚ�����T��1.�`5f���KI�YWԹ}�2{�~b#A�h����2�\<� �20�VۖA"v�?7�ۃ4�"��������iP�p�"@�a$;�����}�*n��� ���d��-��'���|�漾����u��ɬVKJ*�I"ܾ�Jr= �v!n�r�!�Zܸ�Q���D��3+'KnII�����(Зc'��1�"����e�
�o��0�p������d�.�)� m͟��H��#�K�9�%��zO�nS���Ld=2�1�?���<k� \�������y�����%����p��� �U��[%��g�V,�¢��m�Ŏ�Vg�E�:f�W�<ȭ,"Qs����ÑFk�څRh����9h\�*3����������p��t��|�ۛNZ�.S~;+��p���bkc*��|F!�=*O�M��nM_�B�����󲹎���[W���tC�t5@���d ��P0������
*<�L�;U��M5���q`}�/C�p[�ji��kd؛yy�C���`��$�S�[25����	��c�Q>�h���\��	�t�	j�{�Y�5]�<�y����5����� l.P���,�䠔�f������+�\8-�p�-�e?A�b��d�"�(ǫ��{u��#�J6]���pݵ�}Z�� չ.��8<�b[�,�&�K�`G�+i�ۍU۱��&�'�-lϗr8iP>�A���P軜"��Cl�-�ध))��+�A�͢�;����,��tfm!��Ť.@ڲA���y��w	p?|&��PG�&���ښ��)5�Pɴ0��&��r��}λ e6)5f ѪYط�� �0Z����p{}��v��!���[гVШ�y!�;hY���lȲ1���y���������"e~����Bз�M��:K��������էxJ�3�Y��G�WB�@��P�IF��L83�cq
�֜�.*&����0�lH��Y/l� m!hi~mry�nZ�����iƞ�2s�{�[8#]����&��2{C��y
j���h9
�I��!�f�6�O��	�=��(T��^7Y�X��i�sQ		�:��AW�ú��d��t�v�%姶9�B��ŗ�}����4�~��s�) �K�,B�_�U�?������qnv�m`��ڠ⎱c:�+�u�&���&^k�MP�z S1�w��jȇT'�A��m���|vw�jD7�@O'n��o�VE&�8Fy�+k>{�84�Z��~����������?9�l���;��^�����џ�X��	?�M�!Yǿi�㭗�s���2���Xq�R���Z�^u� �hB�}z~)��14~��F(b3�\�e�M��W�p~z-`|�&��َ%�X8W�a���9�'@�?m��9���Ț��{H�A �-���7�PkVw+ڤ�O���oHӒe=��v�%�5|F�CŬ�ڒ���-Z�l���=�A,���ه`��S�X��<�ۛm:���G��}�ټ��=]8� ��N�e`IU�l.��c�hp�{����e�d�Ѽ�A)p��[rΕ_X��W!�����W���V�
o�ɖW'r�n�r22�Z_�o����<ӣ�ـ㇭�(ہ�ey��.�>aN�J����3S36t������cT�8�d��j����$P/1�P�Sߩ�4-v�'sȮ�CB�PMj?(�0'�����*e�R�a�l�O��=�l=���I���
FYb�)K�sO��t��؜�/?���d��G�il��ϒ���䲟Ӓ9�2u����,�E��s���6\ÏR�9���}S�{/��w	(���cЎbG,��/猋��s9�+9��W�c|�{�B�D�N)��>@���:9�T���s���J�ka= G�P,(�8�����^��~�I��f��ps{��w�����RR���0&y77�n��亨D�iE��7�C�i���&��@u �:%I�� 2>ݸ-=-w>���I�0ψ$�^����LX��x�3��M��(I���@+�J�>����Է
�Y�}��wKj�9���z�Ϧ��x�շ�2�Bt���
}�����ث+
j6�6��!�#�c7��ى�YΏ=��څM��*�s�������[R��쎇�:�Ŏ8'���|O�w��ʋ?���z�H�<9�:r�1*��ͫ�Z���K��&�{���~���bK���Ǣ���o���t��}��I���~���r1��M��BC� ]����z�s���4�� ��z蜝��J�L�}H�5I\p�N]e�U4CZ�f1��cvGv�4��c��B]�i���p�->o.��fWT7Թ]�vmfˏp��.�����I��qHPCj����HS�'�zqv�.ǷAj�}aF���J��DχzAW���n��j��9���d/����;3�j�H����<QA@��m^�΍�M�H3`�}��I��̦��ר@�J���ũ'XW��Y{��f�|`�=ˠ��t���-�2�r�`�0���F0ڌTz�Qs&�9����T*���A�i���=�$��P�ej�������|dl��qkAzzd�>�tU�4(Mk�48I�4o�Y��y/�GWg�]�Vp�I���P�c��%_��Ž���&���$��N:�ň��T�f��x0.�b�َ�m�Bo?||�l��Lv�fsj���q&j�2gaFeNP.�3-=E�PSS[Lu��el�x�U�G��}������e �؃�<w�r{g�-�op�q�����p��н�|R�*k��܉�Re}�n~�.](�b���"�7��΋���?��.�A�n�ºu��Gkf��0�ys$�ʻqL�UEa:��^_,(b���`D�ǰ�@^�M��\6�V4�xyqJ�!��Wp�R9i#����%��Ka���?�q�{��� ��魷�4�[����LQr5rb!�gÀ�n��n7���RDӅ=�,*㤪Ho3�7wgL�|.�(�0���!7U��`@|�e/[@'bz3/��2�Ҧ��ϑ��Nn��������j�R�c��p��>q��#c�hE�=��_�@�Ϊ�Jbe�?YPn�R���K��Ka�$W���­�I@90=pYP�+z���ƹ$Q�����J̪�Y�Kf��Fֲ^�dj[J�fC�K�+-�����:r�=P�r����Ĭ�E�=A[�eZ�P����]��4�pJWH���4LS9�49���5)5W>E#~W�A�M��ܡN�׻7UMM&�>�P-��X�0�q*��~��k�'��)��^Ajj~�D����TMu)Y04��4�`�aq����Lſ�D���R*���rnQ��	z&P,�=�������{�#���H�$b�@���&gS������1S-gf�Dʞ�	���]����	�������=�d���\�?�n�����������������������������}�.&F�?i��]��@��=�ֽ�Q���u�e�˙а�K�S�={����L�ym<�8�+!��B�qO:�;)����C�#�7j4G�$�I}f�M�K���`eb�Z,�G����#G2���F�&��뭣�X���!q�挽�~(��F˭�	�k�*�����Oss����N��9�6�����V�xa痼�����h%��Ω�FM�P���ƐK�ǐ����hh��Y�Sk��Sr{�ݛ{wwe~�c܏�n��d|P�b�Ӓv��2g�<��}�NIL���=PlK:�tAe�@��"
�>�u��3,�,�9)�QnsN)"rʧ������gML���ه�:��z��?��r�������q�/�i΁�w������[��ឍ�>���q��7�{�_ޘǬϊnR	PX��P�;��ҕ�5��+*�eC�N��]��Uי�{Ϸ�^�s6�]��M��-R&�:�7��5%;�F��q�2�e����%>����}��,�#Ci�}���K�����K��@C�i-�)�c�=�T�;��DȐ�9�aR���G�a��C!�M�N��f]�+�\�Dy�vf�BH��$�B���ֶ?�2�);]Nz�KIj��A�N�ZagF�r�B�i>4��?zo��Ջɋ��v'�F������
�Yu�+�ϔ۴�T�MLu��qvf���ʨؤ���x�>�Ŭ��
���{&�Ns�������� yG�@�|\\�����sg	��mf�ŏ��Ë����@Hq�G(��άoqs�e���h2G1����K��GK�Zf:�h�9��b�r_�ϫ����l�a1��!�8�}gggBL��p]�&��o����dd��O��o!�����	����@>6��M9�l+�R�r���t�����5�gI�Jc��������[S�\���X�i��
�M���*؜����
ͬ����
��DV�2��Z���di�(Qa��|��+�_�ϑ���b����:���w�����
c]����'��`��8-D+1���D�l�Gu���t������Kjy�ZӃ�}G{jz�C��`{Q`��%��x�.o�l� DX�r���	�%kwӠ����?���͇�z(��N�2�A���j��~�]�r�o��SU(/�'̤�ncA��:�O�Մ��?�*[_����G�we������o�v�X'�
�p�W�d��[\ބ
�( m���:��g�c
y�Ajq���%��M<��'�D����@PzJsV�:�^M5َ󯣃U	"ZZ��*h#��"���V����+)Dg�!��h3�	|˸����0V�2����*~����KJ
���R�k�7݅w/&��W���!������);!����
�z�_�m6�H�Z_+��n���λ>"c�|�.T��~.�kV�
���Sn�ŤƗ1�m+�Gsn/_d-7�R~9�O���m6����� B[�W]��-P�a�"�ٯ�η�a9y�u��-��6�\
Av���< ڴ�)WZ[F�y��4�T�o��b�_���	��#���ԻF��I���_�M�v3�k+ hծ�ry�ҽ[ѓ������n"Q5����ȷ���`�5�Q5���*��� [1�?j߻�Y��'���%���m!�91)	9����k+�P�"\�[!�{Q�������󡽚��MX�5��4��y2�G�������شC4E%��'�W��dM��J�Mc����׈ VΡP�W� �y�J�G�,fm���W��M����u������9���+���NP~�
A�G�w�$B$���)�������\�OW,�p~�8_⓯��_������_S�(T*�� (�%o!W� #.�R���s���t� �����s�x_����A�'`!���L�U0f]��`���J����H+㚗��w���S��.�<m��$�L@��J�t���L�"3��Oa����(*�Ȋ�����&����Z~��p	Xi��1 ��o�C�_q&���tij"h*[P}��FezO����X��r�K�׾_|�ja]���ѻq�YOц���.�:�A2N%�hVs��}�]����C��T:�˯*��O�7\�3E �(�ׯ����c�������t@�D<�^J'�9�Ci �<���V�G���ݹ7��U��X�������j@y���`<�!\��^� �C��'�'L���,�OM޺f�B~Ś��?~h�s�\{��|1��,�������pqۨ�H��0N�/@�t��H
=v��������d�"���[�������߉�K�|ʎ�?��Ż�F �EF��o��q��0���x�����5H�2�}n��Qa{/��R2�Ex3�>�+76�{��͡FC��ٜ�����2�U�?�/�����Ĭ��aS	��mF�N@�vgtEL���7��B��������� �]����߽�;����Y_��qtnػ���@�j6,�&�cU�ߋ�'^�k7�s�u_OO?�s�����Z�C!Z�Q(/n?���ۡF�w�&�nE͗M��F �J�Hg�{��G�@{� �ٺ�3��2�c�V����$�T���~c��@���>�6%%�0^W�r��k����ZS��8�oK"��NI0�`�ay�g��Ъ��o�}�n�\�6~Ϸ�M�!����Um΋i�3�+K�c���ʓ���������T��K
�廇\Y�;�����3��-��X��쒁��ݠ��������� K��ļF��l�H[�vgj���;-�(�Z��˩��wF��b�O��t�(\�14~9�z0񋔆�`���hW#�LQD�y�����N��
���o��maN�,5������6�@Z��ֶ������F>r�?;v�I�՚��|�#̛�M��J�
yvƆ� Z����L�]�l��i� �{��z�v�����V�N�U`@j�������s�d���J`���L�[Q�\��Z����3�B���嵴�g_\Ӻ��������hÞ�وЪ�H��+Y�<ˣ����$A��{�ױ��ة4l ���Q~��I0)z��#˿V��n!�����d̚���4�G�k�>��Ą�ؼCQ<8ǅ�����k��	�P�v�p���FLL<mwww���
�L!VXQF��-���1���L�]�r�H��5�3-h����0�.�5Qr��~D��Ԯ���դ��2<~8'9�����d���qu�� f�y��WA"fH*����w�&��.����s��!���ҒJh���ҝ/Ȼ���nnktuu�g^�#��_/**:ii�y�E$�Uxb�S�V�M����
�� edd0��>uq^���`�S���0�1!1������G�L�ə=[5��笉�/�_�bl+�<�=ݥa��h�F쐕��W9�p`pql��
㔞]݅T��6A���cD�HL�e��f@Qnb/�콙���i�)�!�(+RE%����^���%��4Co��j�cZ�OƓ �͒ͯY6W5�V�vy�G�?�Lu"�֎�y*��-4ճ�32���W����H����Ļ��&�����Ӵ4���w�?o�`PA��;:ć9(�#{wz?f��h~���
#�j�/��a������mll��!�~��.c��[RɕA�Lv��v_]���jޔ�������y�ӓ�!#<<���f�u�N��ț&Ԛ�e�g�P����X�)��4�_�!a�F���>�J`NS]���79*'Zd�	����Y���b4Pv>����������Π��(88�د]Y����v�l���.��LF~�g�_�g"��]L\�Um�	��������L��7=�Z[]]���zݲl/ě"I�I:4����W�^��[=��X���'E�b��3�+ ��V�T�j�_���N?)���c}���p��H)"��x�ԩ��1�'���J����Qߏ�۠P��
��l��ɧ����Jt�2rժU�Zr%V��°�����'m e�>�s���:�C�{��wQ���]N��	i��W�H�x_JE{J�f v����������>��Y�)fć<a��(�3�n� i��6�b0���-*_Z�����L��kaD��lR6DP?<B��mI��5C���xQ#=���. RGc07I#���*��̞���-�Q���>��(
u�А���^&&5����3^���Ky4@����D���c��@���=k�/_�4=��[v�����Q���Rw�Naˁ�,Đ�^wf����&S�<�.^L&���i�ɼ�� 0�$Z_e��]���]tfp��;�HT���5�t�>�[���Ei��#��.���(/+��~� �w>�Ԗ��Hۜ9�@R�]:^� {�d	X��4�1И�B�5��I'�������X{G��\��Gܲ��+
[e)})J�|~t�p�ATDdd�|�,m1L̕�N�j����d�j9,C
3��[�̙b�SB����]/^�8mo��^��99]�(�F92�%8 ��T���]�� ����ʾ��m�+<��`�U���3S�/F7 ���?`hU ��ddWWW(S��C�2�6e���dV���T ���Yb(TQ�=�Au7����툧�e�ff��U�ώD7�{�	����j�5xO����pU���(��熝�K h�v>�lc3u��G��`2ГYY�1�K�SBR�P���xt_Qs����P���� 1�Ԏi�=B+����x'���
��#�1�]u9��b�mB�s�$m���@m��'OΧ5Tv����NH茏�$�s��Q<}�Jk Fh����L�u�2��1\MD?'���m>$�2P��<sr'yy��϶Q��4�@S` �*�"�s���'��3�)�M���Qvt���r3��K�ݵ~�I���m�,��cH���㴭����{�D"�B5�l��)2qqq���7 ��D�@|R�V�]�l>;ҥ��W�*4B������J�B��R�v1I �j�ʌ0����H��%˭ꦬ&GE�$�#����c0+�<��%+}�w}��{|e���T#�Eu���������⎺����I	X�?
�	�����5]�'��0��y889��O�i*( ��Ў�	�5�kIꝌ�+C:�Lʹ�z�e�ڟ��@@� �XP\��)�A���T���Mh��l�� e P<����#0�?m)�(,Wn��0s"��̍<���l9�BT���p;��A�&SR�y�f2����������u���!��S�"�\"Q<3��,���A'��:б�o����M�(7ZМ�6�цdp�L@��Nar�9���BR�I$��xG��1��,��i�^7 vy@:R8h�7s �:Wr����cE��y�e�>q�y��S.��5�;/+ �OĹ���j���a�n;�]�����qfgh�v�� @�%d�Aѹ	���$��E�]<I�����'oe&2�^�d�=I��T��x�g���Hs�pQ�该21��xV�i6f�E�����ˍD��"a=���Ǡ-�*uo��BG�,1�_PP���~󚠄N���!"B�Fjr��N�|���Pt0p7�u+�$E^Aa5`)�]P;�aeb�RS���u^�}Ro&�i���EBi����s�+8X��+B�l9��:�:�'OI$����J%8SZ&	E5۹�?ाLBL(�e��i8��#c� 0|�4�[��� ��
����n[�-�ߣ�0�@��Q���R�*�ng2�i ��=�|�_ ����1A_Q�O�'�,-M0\�������ݻA�Y����M��D����쎕���&��清���/��F+���L��N�N�Nk�,--����G}í��O�4�=P��~�W����b����ک��z������9�&}}�����ޢ��;���;F��23�{�XR�fW�ׄf$xN�:��ȶ�ZO�	�#\��5�5�Zx�$�F��Z�Ύ&E�\8��/�ٔD ��ڀP֍��XP�����^��B�-�>u����A:��ҁe��I����EnG�b7���HH����h���G���roNLL|���r�`������_��i�SQ��K��u�{�,�<�LN��&��&��=�O�@��>^��3~Ƞ����quD�z���ji���O�y~�hr���;��&Xao�篵��C:*�u�}��$a��<���/_���y!�6QX����ud�&m��REEE���M����?7M }w0O8��,���mx�>d��a��W��;
��O����jۣ�XC������8��sF�u���Z\'��E�4қm�9IF�Տ�@3I�o�G�����#-3^y�GQew�p,?�$)�\�?�R��f.��F��J�:L� �_d�7\�ag��|��u�C��l �<�a��k���ƺ������5�6�ު�ݱ'J�.���U���?�AxC� t��m?mrǋ�u����(˓�^gl5UIA�mf���	�?b�)��`g&{��t,����1*�
ᎎ�! 2��I�Ɩ��&�l�̤�V�v�!b��l1�+K�2�<����6�0ةP�8��l>6��>4$/.!��h���r���9�"ch��a>L�`X�񾊢t�gq���4�l�ι��Nͅ�	�YK��h�V,oHC�pe1�v�C�ձ�m��A�w�����o�\��ݛ%<Q���5Ђ��/��-E�K�x����CԧMJ� ݵ�ӫ5w�W��,:��>o]xw_��"���މY�V�s�BS6�$oe�w����{=�'�n^z���\`��T��O������K\a>$���K����S�6�*�yVI�w�����z;�	��[���I��_�w�o��_�^���;+.��m��χ��R{��@�%��!���=<��7�@�%��&�D�'�Hֶ�6�F�M^��u����:��c��&�/?�ٶ�f�N��p(؆����<�p��M?��]]j��}Pr��dYQ�|]�L��3|9r9��>p�0�A��7X�]���o�y���V�q�+%��ٽPr,��!m��v-�;�+[y��~��}}�K�1���hyz��H�8^[#dd������@�ٻS��9�`��;��Xx��K�hn#��_�� �;��ut����g@���ŗ/�o����n���o������?yA�)�
`%<�j5kk^�١9㣹�-�ʧ�o�����@�������y��e:_�(S���H�O6>�9���Q�{�o
�l|Qt�n`�����0����7��pk��n߫5
��}�a���l J�������,d�8H�����AQ�V6Bz�������p�͍�]B
��y�������̳�� �̹G��_��S���>�_� �D�η����T����I\�u��
�S<^9���|�`:ߏ���D<�}{��.��W�����t���n�Z��l����*`xy���!6�_�:����.GȼxiΦX�6P�&D��� �� �V>쇜ݬ�y���0ʻ�kUa�p� �R��v�ڐ׺�K���E�������${������zo��m�|N^����9�	�9%�����d����ޡ8b�f(�[��{>�<���90������r��i%������_�q"��}1Du���'�]yf�[�K ��;ͣ���8�2�]f����jcF�c>���������m���"����W�8�Ւy�ڈ8�=�5� ��Ȃ�)J���_L��y�N�l�S�۵�l�w��+��ϠA��Cbu�^&@�':���qq>�G��?jȤ�W,){]6�4��Y� *��V��&N����J�q��:=��?���'�x[DӏM�z��������Sޔ�{H]}j��"��_�DxG�O��7W}���I�Mkxt��Z���ew7�a��eu�M�dRݟ[k���H�o��}V>e֡��#��>6�>���ҩ�oӾ�<=�b�J$�M�K�\�Z���?�-z�]a��I�(�y37��{ץT�d�����W�/y3�
s%N�4b����t��<t�|�v]
�����F���TxA*������'X�=x�ܛ,�k�ª�yi+��$����a�û@1_AVm�~ H`�O��N�C]����G@���+@��%ށ�>AX���ޯ��OQ 9�Lɲr0�ｚM�_j\>S�k��9�|�h�I�d�����C.Z��2����]�{���E;��}�e\��L��x�!�BGy�h��s�T�'/7C*�G��Nyx��ٞ5 !�/��|Z�Ma�B����ޏ|�anT�2k��	`��_kƹOk6���n��G�V�/��7��b�~Ee�E����BC�WD�����^�ֲ�����6��{���5�������ξ��(��ln��	�D�1�)t�Kl;i�� �n���#`�Y�dz��?g�����
�
c�ྔ�/�0��/;�?�$��l	۟������ѱ��F��:�WF��6O='�k
l7��>�d h�ꗐڕ}��_l��f�����>���F�<�����u���S)�ˤ�ӝ��!��Dj
PsC醹��x��E���A�;�8�v�%�JA�d��R��
�9zy��ҳ�]���s6�������r�B�~�<�q�~����O�QV��7��9��&@���%g*����kW��]���4.��a�`N|�;�H����~��$���?�R��ħܠ��k���̗��ؿ�� �`!�,���aF.�ka@�#������O�#> f��Z�|E)�t0�%��o��k5�8��y|(�{�<��I@�w
�-X�wun�������X�c3�e�[�~��蚮��� �u�����`�ξI�d6�?)楝����@kp�Rz��Z9��a���p�n=���u�m�I�<��|J�<�fėg_��{��F���&h�=�hp�L�.�6i1�d�%$�X��_8���k^,��ټ��4wp��#�D�R�~#ZkK_Sӯ�T�!jx�@��x���N�n�j���7���OF%Y��ɛ}�����n��Y�I�z��/;tm~����ͳ��̻��:=�҅�j�oI�� J�L;$7Bc�$�"9� ����ePF���������/�i/K��x��}��ॷ��yn�,t�H�BEb��%^d�m+Ux�6�$��>Il�>㳑�`d�ʁ���Ep˩���v������`Lm�Mf�P��p�|_�/ ���\ܓ��a��jcjƼ�!tK:�,vh^Ŷ�f��E��렬-<�yp⣐m��˙�C�3ߟ��yK��лe��������c��릿Y�=@)�;����E��N��'��^��h�)�g�~#�Ʉ�yG����u�0�^i�؃���ޟ��y�zA�YS�����S!�ao�M��"g�`���P��= ��2?��o�f�f'[�m_!/a�T!>�@�Ύ�y���d�O!���yq��Tw;�W�Z�my���������%�E�ƍ��;V���^�I[^_�{��7�"�4?��K���͇5��W1.]�[�x����0�##F� <{������i[>�v2��G�8�jp%����+��L����?� ��\�>���W%owT�j���/���[x@��h��(�X��J���|^�_�P��%g���(���3��?����"��`^��~��:�� x��ڌ�}�}��ʁ�+x���A����ὭÈD��b�4�[�<��e_l��ح��^u�oc�a,�3�u�N����	�$~�XO����!/ю!��
��x_,P��.����Vrb]+&u��)�Iv�/�\���E����rd�A�L����ѕo�w}�3=Q�44���dU��F�
�8/b-��$�<��p��[�����d�=������9��^�� �n�)�R��(�Aޤ)A.o�8`v��|q�fq��{[�D���$F������Xc��O���e��߁�F-(�G}-(��	�-���hM�{]�����Q���F��4@G)�2��*?�(,��ur��Ҁq��h^�&����+~wk48uރB��{�|x5
�0�6D�݀<�Z���){�oY��DW4����6p�{z�^�y"������*EVkw��/Qhƥ9\H���xx5ۅz�.���3L��r�ǝ���1
��n	����:�n�Z])��������<��X��Xq���!͉I/����R]�mGA۠�1�j�^�	#=e��Ս���>�I��8e鰵�b����L�2���<����R��dHJ�.�^�Kʐ�/D�e��8V��x�8�j<��{q�����<�/�E��T��I}�A?���YE}���G&�ߴ".�DW1��4+�dm�>��+��ÚJ�}csm�ሂ2�� ����r���$�"�� (�
���Ƞ�AeN2�`��9B�H		����>�{�}�{�����^��?ػ���Uk�֯*U��!�K�|�>���u�O|����^������Z��OE�8&-q�g����`�$/��UJj�L��I��X���/r��
�3�Cف�[ �6�m�F�.J�(P*�;�Y��h�R5�W�\">p"���-�0MEɜ"������K��݊����R�1����&��S[s�#w�GB��w�z��p�߶�ZYZ(y��q�q�8�eu��9Y`1�w����p2Q��`C#""���1����o�#>ǳ�D��Rֳ�9l���r;�*P9� q:4�i˥L������5%��@![�}9�&����Xÿ���}Lx����<Hv�)_N���6N�7�(��^ڑM�.ܵ��뉫dĤ��ޏ���q�<9���=��)��Q��&��K*�|#�i�S�c����%����_�R��9�k��M���Y���礪�+L�� D��7��+ֱx�s���%�������	�m	7Ʈ�~@^����D�$!����0��7%�3*"܌�����Y� .�a����~E�M��`^L�G7�� ���)ϛ&(��t��|{�1�#[�,�6��4e�����z*���lI�����V֚�=��V��
�Z���K@E�u	X@�oR�&[Q7�(�V���+u�P�5�<]�����J��=�Z}턆5d������9r6����b{t�AM_;�߿��i��V�Ujxyɸ�S������ֻ������w����>�I�AG�����;l���$��`�)0b�ʘ��ϗ�T�M��2T���@��W�p���D�]T'�'�T�}����M]V�|�*L�^oj��$�Q��=��7�U�1�r�=���!�����ʈ�2��[����I�'Na���-��Ũ���٤xg�z�����g��U�7o>��Rf��j�Eǃֶ�k�y�'E���`���/_'R$��f�A8(XhX�L��Vg[� ]��%/�Lꥬ̮�T��7x禍�i�/��b��~U}���0p�&'~����q�Ĥ$�TI����@�c �c���P�_*��3���B��*vtx��X�WK����b��a�j]z�������vk�u�2��yy�k�I[ 9ΧW0�`1G{=巽�o�K�.��Z-j��U��`*�`�*ʠ�ƛ�yܰ:i %����L���]:�%�ɐ��J?
S�E	��f����,�l��M�'��7e�Ol���>m���)l������N�eׯ�N��W�Lкk�ޜ�?}�����4��Ջ����tf��!5~Csssg�����2����@p��7o�H�D*�n����B����|�1��=�o5�I�M����%���QdT�ߺ�`$��볘��$)�> �׺�q�+K֋�L���*L�ș�Q���,�[a�p?zt�Mxa�J_���6�`��m:�P���"�A���Q���{�/��L�J~�?pa��5�s?�A-���G�'MB�`��(�r���`=�C�%�I��~�q}���I��58�����In���
��I�=��c�2�;66V;C:�箏~�FV	��E��*/\�/�h�(!����	��N���( ��R�^h8m�V�Zu5ֻ���?����=Xuwa��z}o���q����ʻ3�X	�FN6�N�q�n��(����3��*��'G))'??M��7ٞ�:b�J��������\�n�u��Q�Ԕ$K����+�-/�RR����sM�� t)m�`շ�r��įC;�S����K�%�g�'=�OYs*P�U�o�Ye�n�cw��s*	@kq������G
��V�I�A�k�wDM��%��0�B�ׄu۶��:���!�#:��J�_���>Nqʦ�I\�'>H^���#�7&���t{�>����c,���MMMSA����=����f��x�Q�%����P�Z��2B%��e����6#�l�hnz�p]:p�����s�-^'�%�g̸|e�v�R&�`�t����z�� 6 �o>�Z�����ܻ _I]�5�z~q	>�C"߮l(}F��v��{%�M>Y���= �W^�t~r )^%7�֑/	�}����m��b08{�=��>������Ѫ)�:8���*�D��Dݵ:	��'���_�I�|q�̊i��q�1��$Z���� %�D���5���lRMpP�	Z�_�	
{�}gǴD4�l1�=�3�(U`��OB����S�,e�4�T��	�jev�y�����O~|���(��c�5��.�S���#p2<�s1�[�!ǎ���D�� ��~�[�!sC?K���Џ1��Y����2�E1�PU�����`" -#�]?���a��G�ېW�� E���7�_����L�� )FE�m���V�޸�)��X�:EC,�߃-���ץA'���8�4F2*Q(˴|�?��#�M4�x��|Q&zௌ�P�N�Q��~����ba--n�ys'��*}	�|��ězg����vY	�(�@'�1���eC�����8/�j .�q9�������ݤ�AIh�(��(WG0杳�Z�A�g/����.�d	�$��1�.��ԡz��@�s2�`ʳ/*�5���V;fQ~�:Z�"��{����kP�� V�ea��a�ꞿ�̿����~����Q#ӡ��򺓐b)p`�`�P�fЂl8�ֱCPV9G(���hM�eX�[@T�G8ȫB/�A�Yd���}������o4fL���4&Y�f47x�ɑb���H��A|��(˳�f���{����luEb��(�b��*�ΏP��
��=CN,����+���b��RF�+ �d�I�i�r��q1�x�4gQog���{��S�l�'�;��8<,&.}��4P&�S�.w������I�X'��ʼt�-?
Y�ܯa�?���^.b�F`b�;qaf �o=
)�x�a	j�`��� ���5�����_�	�3���u�2��SR���L������/KY�����ԪP�\�P\D[�@�{���;?�׈l��������W �zc� �جm��2�kGA�g�wy~tkG�ڭ�G�[�Y���.q�r��zv�a�:��-�:J^����On��{��n��8u�Q�a�����L�����%��V5��ѡ��/v�Y^��"hSa�Y�#�x�e�g��D.K��/�����	��Ē(Ŭ��&�Θp�s�/JpM���Ж�^�ho���R�sGǑ'�!�A�����#�=J�����c�OR}e����+��ݹ��F#Z��%g�����wkoƄ7ekdtU��q�2�*����9qC���N�M��@0u����ʯs����JY���=�B}[w���??w$ԧ?�S�iA���y;�0�����bL}�>��+K�>󄹹��%��O��<0�Z��)��~�#���dۚ��V`��R{�����jT�za>��n���l�n�-��Ź��=t��[ny���|j!�?\g�v9u���ߤ�z��V�\h��%�ۻ�љ����i_)n���^��]˧��۝���l7 ��}"_��t��7�]����mK�8P��60'S �eೲ<و�#��(!��3��u]�Yn�l�v;��U�S�"q�N�[���NKd�(P:ҥ�����n�{�\���>B�����۟5�Bޤ�+��E!������'[����y�e�O͕�,M�;Yj�GFa�vlp�U\t�(S_0�r�.r�b/\_�\i5�ф�§ϫ�''a�~x�;�E�͠���龧gTc��t����с�n��B��2���oܫy&m���#���4����z�y�W�����s�����x�@���<x��R��y��CJ�	��s^�h,��P�%���sQ[���&��G�ܡL�*tV��ǫ���ݚ�:d`�~���ߒ��d�6l�Y��L%<��������v>^��������|�~�ͱ	xw_�����D�IYz0����X�=ٷgg+)�{M�P�)�qL��A{���Dn�*���=/�caFH��J��~Xٴ�����ħ#�"~ﮪƾ�%%j��[�@'`�^����D2^��d[c��@Ѽf�e��SS�������`�n)�:&�[͹������XI��҃���vS�^�g�� BH�����j]�Ε�N�N�c~t��^E�R(O]�^�΋��G���,7@�t7��1�"��}Q�j��z����5�Qx��$��Tp�K^ań��J0��_�'ʑ~�A�j�8N�F�z�d��e�G�y�ȧ����HǌS*OZ�;�W\������"�vnTۥ�f1������=�� ܋��c�V��S�(-�2Y1�%a�/Mt���jl�JĘ?�|���J
S�e\3y�Q�,�TQ��K���@jq�=�����]��&v䒾����鞯�������8v}��P�[U�ߣ(�=">k��f�߂Ѫ2�͝����N������ݮrB`�/1Һϝ`��w���	�(K��5���h!����β�X�D�5φ#�푫�r�3Γ����>S��"
�P����`�n�[XJ�d�ݍ�Q�+�	>�8NF9�|��H�qMۅBX�:?�D����%U�V����V�Ǖ��T���Ow.��x�\�����-o"��ӎ��Np�"��h�/�mz�a�+��Ƙy�f9	��o0WR����c0�	BwV�$�]���V�*��m�=��~���|s�j�/aV���+�h�͂�R�w���w"���,�|�Z*�c������\K����Fy��yZ@1����]6GU)ڨ�!-�#�Մ/"��������?�����ZU�ܞk�P�?�hmח%�TN���7��1J��/,,��'⸾�KK{�!�/�vZb�����5s�@�W� �������C������g��w}�ϝ?O���IY��J�����/�,?wH�ym����{B��#�[δ�d��kM3�gΕ+W��xw}~��d�G())��\5��֋pL���p*;��9��Ɯ�,�7�Y���&C�lt��p���s]�X/��H�rS.�a����%���$	���@uD��T|5����gn��OC�׎U�jp�Oݭ�΂;D"����%zy��6���z}'���"l0�n�^���|L��	��o���R�܉΂�߱E�-�}�l��3G$�;�w{�݀��c[��K��b���ӥr���p��Oa%u����'{RRR�	�$��mwf�B��<�P���Ca�����au
���Ȑ�A�ڋ�i|f�P�ѵ�Ę����|����H��T@��E�{��jk;̽��E�D/R��H�b�xOk�w�|81ϋZD�Aj�� ѣ=7\_O�L�=�'�)l<?�wTC\N�:r�1��7�`{��ɓ'�[�����E���f��3�-[���bC�k�����	&�(�|ľ�3��O�$IzQZJ�@�-��Oii���!D$��W�G�����a��偺:RC����OpZ	 7�ؠ��H�Ș�؊O�=�~���	��(���"�j
�=m��|���+�
�϶�M"��	߁�d��$	)f��������S�q���i\�~��-�`�r��y��ڍ����].L���r�(k{{�&X;�#��`��-u�0r�X0(�N��������e�P�(����lœuTu��oAh�R�����f]z�L���$� ZG���U#�kݽ��=>=�l�5�L���f��/���D566�h��ބ�g"Q���=����ݣ��ޚ�����EN���jp�77���J���`�+a�@�m�3�������G���Eq���d5k��UH�<H��s�v6��|�S�-s�w�ퟥ:Gͮq�дLX+ru<^�#m|��s�	��75&*��;��[�=�o�kD�����ve�$�]ײ f���9�6)�U�^��e��U����Il�>������t$]ۣ3�bb%�Z"k&�?�2�����g��X*A7�	'D9��

bY_���)Y���%�� Yx_A|!��;�� !GwSJ����������D�Ae�e��@
�:9C?�)�ޖ��������.]�e�p�,,,h���َ�@��Q�h[*p>7����-�b{�g���Ucŉ�/kdtv��1���a(*��PfFZu�R}���A�d闓����U���!�=ؙ��E���v��3��a��q�0#�Y����?�$	v���g7h�ٓ�D�5|>_` ��d1&'��}m����H$R���Ç �|��
''';�-�7��F�^��K�Iutuu�2��L]`l�O����eH���G���ˋVy�zb����W���k
��O���Tuh�k��i����]y1r��g�s�E�JIH���)��?�jS5�Z%��M�g�52$��;�o�E*4�����Rw�rLLL� 4Wfz;::bhA�,�1Mob^��[����?�ژ�pSo	*zC(�Z�kq����@=Ka�ь4=�2�R�ޗۊ�o��	
rd��ױx
�z�9⼟*R+�Zx)q���o���}���I���PK   ��!Y�&�}[  y`  /   images/982accd3-ee7b-437c-8e9e-7ebd1fcbf7fd.png��W���x��,@���$$��[pw'h� xpww����]w���{��p�sf�L�tWwu�S�]���(�P@ ����2s��{����[�<�[��)Z���@tq&����醌����Q�ܕ�ã����0��Ќ�P"��b``�E��X����t��a9�檗�����EV�����*f7M�?!��ģ��JHH�`�s��m+�>=,?��8�B�ybѣo�h�I����7�.5.��}7�O�3�����1�]��fPz���	l5\B�zB���Ǡ�9�WQ���t��ԇ�t�D���=$9���y?����K=�`�?y.��d�bh�h�� ��;|4��e44Z7���A!Ɂ��Lс3N���R����BS����d�����_^��Fe�v�����t<����)^�"��y��(�N�Eİ �7�R���h@��`�(
��@�� Ё!ğ8��(	/�e$�A�]wb���?d)-g���#���(Dr�����C�G���!I�_��������{'{sK��.�f���P��z�>�7�Pz/x}�^�ʧ����f+%O)%�.V�>�9y 8�o�Y�ڢ�d4q}�o����V��؂g`�`࿘��u����_*�/M�ܛ�C�M��T��0=��������,�.^��_�������8&3E���1]����ߤaV*宣�K�W����?��P��|����������gi�j��fJeSk�$uQ��h�/ڳǠ��S���+M�x��}BM�9�+��rE�4dMӌ�����b�hp@���/fg�����Njy�|W"D��=P� �LC��˟@2b��+�U��=L;S[�1}?�	�c�'�z�ײn��Q��I�g���)�GD�!����3KWEc��Ǝ�YXG����w�W���qO�t���?�z,�����=#�Mp�����9Iq�����]fn�����\QQ8қU��X-�?�瞭���ܷ�Y�}x0���]���Y�c�����MY�W��Q����G�E\ж�aL��f�y(�3�_������ţ����6����)A�X�֕z�ΉJ+a��©�����\l���f:-��¹�/t ���'"�vy5��S��Y��u�èh�z��x�ۣ�ni{0xq�ʇ�|��_#[���%����*��5� ѬXX�'����K0y &�>�NTm��Q�׋E��j�@�	�����z�f7�*�������i�ǐ��	z�M��)+.���"}Ƙ�s��̥�b���93�R�R /�y5R��w�>�v������Fdt���v8���ډJ$J�ݜ��t�+�~�?<��la��綖Kц���x��+��0Z;H�fp�;����7.�c�sϋ����?L4j�ctҲՊB�뚚�&�n~��/H�X�A�uM�Y�����5�W���a奫�r��E��泑�'�'CR���:N^��#7�2�d&�o�ȩʓ��_���ne������;]V�	�%�R=r�G%N�UH	�|:��}�$�$SX9\:�H\�.)ah*-Ywkݸ��l7��TrCnElN9�����
��xwy�����=����$�a�V2?�I���)��5V��'<<'EI�I���%���-cO3:�u*b҈�Kl9�@V[�~%M���0`r�b$a�k�G�V����;-����m�'�{����6H��ca)��rw�p]�s'%���R�զ�ţ�L�L��Iծ���_�me$-:���y�'N|�ޔ /�B����(������\���y�I�f�f�~�ٸ�(ka��o�e�����{�)T�,K}!Q��`@6p���5A�`�҇��P_�3/A��8yZ,,,.1FF�Б}��'?�-_arFF��#��k\����~y�STf(JKI��efe�zQ<o��F8���>�!�lU�{�)�p�w���,.vj|?�!܉)_�1���ϼ��+{HQ�W�gmq��@WB�`aVN�)A,��<�:�^�Y��CJ,޸��o(ǜ ů��gwm�@���8Xt:U�.�3/_V�X@Bs���8�&�3�`^?�k�of�Z�0���%��2IL�P�������d�*�5�-M=���m�D��I@�)4�
�wQv".#(t"���k���R��,�WR�	 �ϓGEe%P=|��^;��_I+[kRk����J~��(�:I ����|8��d��%���z2=1�+�u���k!�p�P/>�/#�e�4�������5��D��t��*ɟ���8L�WD0�OD�(ɀ�6�a]V*�,_�r�קbC4�\ $�1�xJ,SR�r��z���oTgdS�[���C���m�:-���5�t��I
�KͿBʜ^%�*��'�����4f���Q(`���u
hR\.
���쳜��dMV�#�������IW=��x��1�ʐ�ߢ��3�����B�%L�D��!4�0+M��f�3���o��&x��-����Tl��d2��%E��`W걆���	�ε�O}�!9b��7���ʷ5���$˛j.�����K�8�j����#�psJ�{"��<|��[�v̆[�mIR+�?v��psL"��kDs�X��ݕ���)����2�_0E���c�3��Ȫ���ϧ����t;�	
�UUUlbb���n�F
66,�jA���IL]N���ē�E���((s�ak,)d o�~��oR��}�Ku=<��1��Y��t����K;y�V"(���n>��0��W+���,�P���sB.+ܚv�iND7J�M����w�r3����'{
���k�����-���4�j�cm\|\Ѿ�o�s(��+�cz;�7�������ⶳGԡ�5̙�~����@8�.c��m�� XE]m��� �0��a>�7}eY�՛ł'�äa�.<�L��ۄNm}.���0s������O�TUL��#�\�������.'z�	�:ڽa����H���x:N���w�ng�4���$�S����',x@���2m�]ەt�QO�ϧ��zkZ������ HS�f���`�eg_�;��l&F�� ��۪�� 0�A~�����{8ܙ%I�[��������灚��|��<��':�N��o��P�4L�Q�z�������4�c.�{6�?�2 ��U�Tv_�&y��v�G	?����W���4�apP;A��U�4�K$�ԧBG7�%[��r�6k�n4l4��i����=���d�0�����V���`���C��s)I�=�%/�4�u�9H���Q����'�,W��ЮY�B^ī܀��;��@��T烌(�7���v���98��Zݾ��1�����78HEC�xR�����J��	E'��=����Ϫ@*�^/+�:*��-�C������r�(�*�~3鄖>{�q�/���f�H�ܐyV]/�����ްd7��r�ߦ��0 �jfjn<:_���2CYV��Ç]V�v��+t��%s��k
/�w�{&[�s\4�)A�k�=�v���-7�#7DW�������"��yZ �2n����Ir_�ʗC��62B�̘�<�t~_�����Q�l$Ȏ����%>�=v��TpZDD���M�Y-�IF�/�pq�{Y���<���s�OW��Ef��iΉN���ߥH�:�0���(�8�n�5;�����;w�+�O�e:OG����\{�B��S��h8B�ޅK��NC?:=\K�{�����x�?#U9l|^}��r��'��c��)�=�Y��F"�쩅��h�n�x�ﱿ���ܼ��B��˧�pPx�����C�!��Gx��|�%���5Uq���pH��}*��^�{V��cq៞=����U>9��e�~�	��b�u2�++��pR�ȼ�굺�9J�ޞZdn��w��g�C����R�sB�x)�vb��/WS�֘Em?`�r,���]�<��C��H%�>�b��)�13tɰt�?}�2���x��iz��V;R}�s���7���&g?)�]�>^�>����c�����X6������I~�I�%���5EA�N���l�b���ͪ�\�N+>kr� 77���H=!��<���,�-0ߕ��D��II���"aK[|�|�3�e�_��z�;�hO���a[~���`�Lb��e6#H����M�M���*Hd��.^�$`�8�{=�r�w��K�~�y�b�x��>o\>l�{m�`/�y-w)�z)�ym����8I��N����[ �:x/�=<Ui~��.��*gM�E�77��El?x��{�&&nظ`X�iؠi��n_ن�8�p���n�t�Ab��K�Pd\;����.��o���BU� Y�%F��Bp&>�ß���]����k�k����ֵ�}�APy����5���K�M�K��k���r��jIy(C��EO��N�/��+��sU���ؔ�¸������Z�x�<A��u����d��:����t�`����zC�W��_e�.���������vY�S23cA�r����(hi�ظu��뒦/�T�չ�Z�M?ub�F�(n�f�-�u��>��f'L�������0��:����d����!�J"F����g��ɜǒ��9�*�a�2�F���������d||��>��hd����T��cw��J?~\�ή�Y��no�j2���dd`�n�>R~mH��D�ݦo�>?0�#�����c��E�jR��� X��<xkpE�fd��
��b=*�2 a�SW'@#��E�������|m��R~L.D��8��\��ݿ�Zj����'����ic�����'�B�5�% ����0���[�΅ʒ��Җ�3�I�R�R�_����)8��LLK�\����o�!�����~���x���C���?	E#z~��*�f�.ɫÕO*�q��ɡ�]4�+)j�n	�ܪ;/������g1e�I��Ӣ	@����n���v���}f!S��G,��"�\V�[��X�|
fa��"�L#K(i�X���|��S���r���^������G��R(���O���moMR��t�Z�8n>����U�!¯﹣�v7��76I���x�y_�B�������n���>?��|	J�+č��YSF!��8�|(��|f�C�V��d>�{�U�w(�xx�
�ď*�i��=Ճ���,��1B7�}|$������8%�A�G���j?�KȥBIy^���m�7�-.�(���EA3��3Ӭ��ot���m���Ә�N'&�2��ڣ�e~ge�'oY��/%���$t��j:�Y3ꉠ}�F��殺!��`��xg����ua6���T���w��j�2��KX�Rh8��2Yn�F�Ie8y��2_�&/))�R]�N,��M� *�� ���v{68?i=5�nD�2��ed�:�'3�h#"ƻpz�Bと}�R!&�����'4��[�oڮMJ�����������b��$?�_X�78���؋�U�D*�H$ǁ���I_�Dz�ɳ������]\\�L�z�����̒,eL�s���ꏈ�^K�G�L�?��.��a����贼�6��z�"��\�ęq^�_�*��q�h��{�c{����y�
q/mw���0��2w*�`��Ĕ�/ Q�4�����;M[
��L!X���kt��k��
�,	������D�qh�?4���r1�U<��֘썫�M��d�q`�+o�����4�3'^��S��$�vUGGG&9���Ե�`����_B`�����
�V��@C=��d@A�mk=�:i�ޙ���A%�oe���^�c��~_T}q$�B���".�g�de{��qX���.�􎏅{(~�<����r��ŢǴ�?L	��7��C�fo/,c��R���&kπw�o�ӿM[P߾Ϥ/���宥34N#�Me�O����l���O�MFe��z�Aڊ�G���p\H$��g ��4��[&�D���5)=�gRS3��}�
�f�fn�V�����T������bꞘX�.�g���^�����$2G;���M���
��`JJj3����2{QeU?�rS���fL�Z\�����tfV5��	�wk
"s�I��Ѳ#n2�_S&c;?0��{�6�}(��r�KZ���H�|;��& �����kdw�6��>�tC��-Kwк��R��˵���v�VzWhi�џ$^҉�	�:��l�s��am�ߞ��Cn4�	!�J]�����X�'Zī_��>�a�����zQª¸9�����B/n�Y^��.>��������4��� JBq���P9�W��+���'$�J�Z�T�L=�J�2B��B�x[7��_��/v�aTv~�K|闦k�g2��W���Z���صh�T�{m���:ָ=�/��W�%x�dP#G�d��(��4�K[�%���}�W�Tg.��� ��|<m�����P����"�y�9BIy1�s�g�Hv�v];,��n[���D��7X���?vi3��b��A����>_��9�ȸP�#�:8ty������/�+:�g^�~e'k�ħ"v���Z�����Z��{j�#���_���
�d�wJ�Q���N;�F*��*`S�"&��V����{�y��V�Hs�y�b�8\��~/7V���o*�֎j6v#g�{�#,�E�,��-��d�K7
�8nFA(�k�]%��TA������	����E�ʭ���Z��ʦi�D}/df��vB0RǮa�qw.�rx�pZݹbp`��<�Xx���I@�"W���b0;}�n��ZA䅤q���fM���~"onb�p�K���a��#����V�Ksj��l�Y�W�cBw���!ʋ6�\���3[��������|�}�ƃ[+)zP��,�UC�R�?9ϲ��=�g9�Rμ�|���@B>'ܚ�������EM��У���*���Gk��-�U��7��MwiF�K�����*,��ka` p\��;ط#n3�^�̗����D3/�%'�e����&�*�&�v=TWm��`���<_f�����֣L���fH*]u�%���tj��ҨԗRP����e&p;��p=A+V�2z�&��56���cf&xI��C�%?c�A�<N3�7�ԸEHij�R +��@s�)(`����,q.lؚ�E�*�۠��[����A@�����s;Rh ����d�x�g-mup��o��h�N8󜳿e-��~�pvlv�JL��aI�~��+aӿ(	3O�I�!3�,Q����#Qp1�;VW;4��}�(��O�Ϭ�z�/�,/O�|�i��%,���h��ƐF��>N��@8�C� �@+* #�\ ��sz�%����Ca?�����]���Ȫl�0�
M6�P��uϐRn�e�A'�W��B����څ�U� >�,䝚ʕ�=�	P�yO(h:?�]�\�@��zb����Se@Iy�y��yh%��SR���_:I=�(kl�Q���\8Ԅ~^�g씈�Q�v��_����AeL ���i|��d�c��ijfƣ"��/b���j�������(���{��q���Vl����FiG�&!��{��s���en�Տ)T���hZ;f�Z���ӵ�w��
	3�"*��l���22��)̫S�gѣi\s,��vAM��U#�r+r�,cT[e5�5��"��&����js)��ǓQk�Ro���h�6�>d�{d��T9�b�˒uڔ�1[���Qr��y�t|��e�3�5��l.����kA�޷{A�}W��}m7��}�;_�î�1PcE��.�k\0��Z�	+'h[�'��"w��O�^��3�#b&�t֗�Ǆ;&�*�H��'�]���i������K�C����umm'M �\�M�3.�%�G��2XΑ������H虙�d;`�[�Gq+�п'B�fk�p ,[�u��~PU�ɩ�ڍTc���eq�ys��9=n@����`�S� ��-ڎ͞�s|��9�)o�` 3X������ܺnG���;��RJ���ݧ��8���[;���+t�[�SR��)�������%w���ݜ,�=��@�����3�j���-�x��6�.8��4ᤎ%,�4f�=��30[�	�g*<?�����ɱ���UDw�Ɔ龠f��Rѹ!�Pg&�hg�����xFg���V75"�Y>�->���Ѧ\�ݑp�\�������Et�R�h"���:���3E�͑�ne��c�g���4�Au���˼,��-zc��429��/1"FA>���JX�����iX�n�]��g�����E�I�w����#"�?�yYY���t�H��u�K���sz@J����=�{Mm%~���lg��I��5݆�%Ɗ�0�3��FcI��1�`Y����Z����2��b��y'~;G�4I��[��eU������׎Z�G�*V\e�zM�s����^�!T�Y?��c����_q_���Z�) ��村���!?���w<���S��t��G�9�rc0s�$�5a�彐��|̯���?�vC������m�<��6v(��ZҐ�:��~K�����>�i�+�Ҿ"E!�$��Q��A���r�|����Ö��:��7��K�����Ճ�P�eWa?׽�u���Sޜ���bL����I�ZUL�y����\��e�۹�"�p��`���x�l�'�K�}!���Na�� x��Sn׋j����BQa�y��V��1_tbn;�A�l��z�����T�zM��0����¾^�2��B/M�8��7��f���n�h�m�tC��c:�L�.��͒��5�',���/w��}���%́�����MO�Kl&�œڬ� ���s���K��\Ee� �������+�k�RU1�A}y��~��M�O��:.h֡^l�!�����[���s}��/�Znv�vWܐ>�Z&{��.����)m�!���_��:�S+j���>���f*ii-<V�(Z�L>n$u�h`��5�A�GD1s�����z5�o��!C�����n��7'+�D0�\č�~�����$"tkpE���:�l��#e�w�p�is?��i(��a�?��8�%$З�%n���"�ܔ��Š�\Re&��Bj2�?���['2�\z��o_������P��t�}���#0�m����J}�"�_���c*ӦF���s�t�ڎ�=�.Ǳq1��KM`��j'��9�"��]E�J�迬��a���3[�ˆ���%�U8��|.B�
j�F폼�e��zk�(;����쪢"=e��BK�F�k)�������_	\c���B3�/·�bM�x��5mo{�_�b��KK�$��\�zHaT��& �P���9����Y�@�kZEE�	CT]?����u� �c"����������I�#`�U�Gd�R:םqm�z*�(��H��QaM�ڮ��2�r� �I>��;\����aGo��cf�d������l��t�k����!m�]3@���mM?U�DH��BF� 	7�wqOD���@�:�w1?��g<��;��%�㚰/�)D�*�#RI_�Fq�?lQN��T���,F�p%A�.l�
�~^á��j���gɵ_�q>���b�%8؝���@,*�H�
W���]]b�����3���Z�	=EK�"��9xk����ۖ�����r?�AYI	K]�3�g5W�F��Z�ZZ��gypE#��(!��=}(���gX~��&�/_�.)�N;ol�ޖ�رk9<��Q��4���N�	��Z���t>5��|�m�W�b!�`.g=3V
���3�z�c�_۽͈K�Zbw��2h�u�4�P��,�V�m��h����t�+]Б�K���� ��T3�|�_��������ݞ�> �$��3qm��-�p�~ 0���E8m%&/�C/4�uM�g��5ب7��=�ưZ�g\�Q��iV�٢E�im1
��NN_�}{��!��t�gy��j[5����v�E�X�ڲ���#��LH�*�zw�Iҕ����������$\�h�5Pn֔����%�E�ʢ~q��k�>ߒӠr/�	Cq�x�m�俙t�q>��M.�r���eu��LS�v/A\>j������2X&�����,{0dOy�#�oY��UJJ��-���q�{�F��CۤE�|YB�o����:�g8����������!�Y�>���c޺����_p0�0�B�0�� �H_.q�-��NP�qɾ��c�-��wD
6���.e����m�R"9aa�0�����IP�ԗB�|`�1��(��ZD�v�ߚ*�Z\>u�=ah�kq?]��'��=��&��Ňg�@�>Zح�JEl�,��@KK�*��h2�s�����eU��~�o{��e��ȭ������T��w�����qTjR#�7�$P	�b��{�dLwU��IS�ݵ:K�4{�D�l��?U�K��l���g��A1�a�D�RK�N�369��d��#9g,OΔ55�3�	;�j5�vmPa~����!���e�-�~l5���D �>6�r i��i���wY>y���ɍ�$��4S6�V�3i�&/I~��AT�_o=5�����1s��]����<��\�F;֖�V��ӵ��v��#7Ss����ZͲ����<Q��5XRUc���pRah�����T� ��KVI�]���'Y����U��+--r~�;t�}��' ΐ]ˊּ��f:���vQ�GWpskc�l֑���������h���/��$LH�C=� }a����Vg�⟕";��N�����J�z��UF&;{�DQY7�'���vЪ����YoƎ;%���[/���j�{\>}��¤�y�M`Ż�]<�"��**��03��ʚs �9ɕ����~�����(~��H7�LYƤ�a���G7ɽV>A���-��56U�K�Y�;��O~$�����d��c��y�'��0)�5�������z\jHr2%K���&?Q��wؽ��%�.�cN���~��s�ϐB�¹sPRWW_)�?�C�M-�z�����TGm��^욐�X�aŭc�F�(Z��O}xc�9����7h�Է��(���F�%��{y�����I�3߰��+l��]��Xܰ�+F���)����)`�Q�<hI��������Ia�S(�D6�c}Jl���O�I^�����1e��y�G?\]_��D�Tx�v�ȫ�Vѐq��>�N���C���mv�y��q�-���Y\BteU���^�=�L�{8�h|A����[�W�ݾ1����)H���r�m�NVr>%��Q�Chu�K�'�7�h~ˆ$�I��e���l���SD	I�Zs[Օ��ދDF%U]4=p/���	!yj�T�_��N��X���V5d�;��k2&	=<F��!����e\���>����z�$B�s&yL���P�$d�o"�K��%�-��D�a���p4�����''6�[�(>�W� /����m��7�_@��o V�R��>��Խ�,�2�9obleQEiU>)����qu�"0)�<��hΞ-�Č5N����V�Y�-ɟ��"&qtt,��|=���X�����-,�{1�����N�A�5��I�|���n]ƇD3;|Y��ޤ��Kᵚ-�ӷ�!�[���y��ɡ,s��	$m+QR)���i`K� c�:E�l�yuU�g���s��C:���R�3�=m!�r����ҥ�oS=�H. �N?�����_�%C��.�|u�:t�H����JD[],����r�z}�J��m{\�ޗ����lU,�m�h� �b)
���h�ؒ���L`lB
���W[GS.Δ�vB���m�<�����|v^��w�R�����֮۝��Yb+ ꀭ������*+SAN��Gb���z����f�V�M� v|�����*sj�Ȅ#mLJ�'�_>;/�KH���� ��_��:p�v� �R�xZ��6��Q�kL�f#I�3P�l���3?�qDޞAVJ5&�g�5b�����Bщ�]����c�aׇ�>��G��%���#	��Y���r�S)-kCp?�ra�ЖE�w5!u����C��y�C��|�5��71Ye#��=y��90�]��rk<:6��d�޼�QQQ��0̖Z��D�`�dH ߛ`<�;:򁚺a��H�]�j�W�ym�>zY��~�}$A��%�\�c�tDMj�\�*�oX��2f=V��tcE�ҘW��d�u�LF	,9�Y�@%SP��!ί�� �=��A��QP���[(�v��p|���R�m/��XN�")��`�+KN�j� <O�'�G�?�SSS?�Vh�6�j6#4�-��l7���C����hpQ��L��L����:�#��;�W�<�&x1��������ؘ��b<����3��z�zu�4Xe;n�m�Q�Ҵ�Ԩ����q���g��lN���t������1<����s��v3޵��-r���5�1���U/���D�D�!�,͸<˷��ɳݶF%Uվ.y&ʀoo����_1�ð~[M�����z�6���A��C�J���w7�ᱳ��~I�=���D�����!a���`�X�eP��Ю���z��tp���ſ��m�@��lQ�t��w���tw2���G͍��d{���p�H���5�H_o��uI��������~��qd�g�Z�\��N79�b���?��Qӌ1���ɔj�Z��2/�I�:�B�VE`
#���Ȯ��芰���]����b����Xma�U�گ	��~���e��	s�%�9�=��^�LT���}{5v	@kҾ弘�<K��<d)i�w�Z��~��2�떠�0EE.�k/�<(�Y'���2&1���w���eip8��k~�uz�DЌ����q��6���7�{X�5w��������=�`7+��"�;�K�F�;(�����!�׌�|/O��G��KR����-{�$�A����n/sɬ7 �T}��0S���,�;��h��rhx\x����[4J�D�糀
��R����j��g��k���F|��.�02��M����7���X�!��(˟_!m*������V���[��7����EN��0�}F��ӓ�v�z���vm/S�M�
`é��P����̯G�X�MfU}�苠�0���\�\~y�`k=#H�y��P�\�:��\aL�J��@�~�jȢ�\���^&��I��/ (�E.~���/����g���EU �z��A��\�(o�Ջe�iLo~C�bi�qq���d�f�H�E���Z�_~.U�!	�&���e>�2�@�_ױ�~��t�_au�	.�BE�N_��e�P���ey�;�6���|���8��'�`c�j�v����3�m��\�[e%[v:�D�M�5~8���X��~:�˙�ͦ�ذ��k���ډ��0��J����^�k�{���J{j�>�3w>:�|�9|��]F�ϭSE�'H��Ϥ;18Ȕ���o���X�ҹ�J��j��[�i�1�F�;31?��x��Gj��	qM����> ��v<8ތ:�A�b);��xq���ص/�5_*��>��&�����A�r1����[X4A���SV7ç�-�ȳ�Ê�N��6�������0F�N���'���Y*��*ZOX�F���7��Ⱥ�xV�����XK��xK]�{��z3+�P���{���Иl��Se0������!�� ��h�z��^x��4:�Iؠ�W��F������K��T/]��^��;.�i��}�"�'+�[E�1=UbS���ff�DF����IO�WUW7~y�լ6��͢�/�d��`;�[��Ubu[��]����JF~oII��D��[��w~�}���$~6�a`�������p����Ȃ��TP�3��s6Fntb]it��mѕ+?W'�O�q��d�w#��v�P��fD��5��V���U�jQ��Fb�Awe�����ȉ5��aY���Ԗ�x�\�M���,7Ϸ9���B]�O_�1�I�)������/���)��B-��������q���ME���~~0��D7�U��b ��gs{n_a�0���7u������-�%��t�ѳ��~�Qe��e��Df�aڻ!j��M��t�M�դ�̛!����[SS��XaTc��6�95H�]�E��;
���ȡ��e�����'�W��ĉ�����.�= m6^80G\\x4rbFJX7�Ka��2��?�lB��g�;�����CF2��f6o�l 2��?������O��C��ͷ�,��R�͘%��t>g �9��W%�����-~8����h��Q��Ͼ���_��:����iz\��i�$�)+X�-9y؉��z!��E�jV��$y[l��-���S3�`�%�wU�Ԯɂ�a{�!X��oap�9��t�T�]���`מd�$2��v�0���聕��b~�`��c�P�k	C�̤.+p���}*D(�`ؚ��R(z��0��h���O�����gE��*�s�_�z�Q�I�k��9bh�း�������y+*s��̭Y�wyP��S�N�J�����r�޵�4�,�3�qo�����Y��d�C���Z{۰�S|��+��ilT�4�)�o��m�>�sa
���{����d����M꤬��N��{��\7�g� }ot?Z;��X�53!wC��4G\�<߭��,��~KԴ��v��<Q�Ê��au��J�斈*�^�v�J�\	F�0�f`d�8��=e�a:{��E!v>����p��)�G��ѡ�'��ÊF��_X�޺�¨�v�@e T�)a�p]���	�!�ޘ�$�N���(ퟦ��J��wW�a=s�pQ..�_��hE�m$M
l��w���m��e�(Vo��S:�"��A�}KR��~��vq��t9.�31n�Dg&��X�p=Qà�����9r�щF�d3�IJ�k�Y�A�����'�G�!"��$�UX+��_����0-���:9�!ÙuQ.(�̺O��Q������t�UϪ�r�հ�a�7���/��d�4�>i��Ɛƭ�|ñ#��r�-��|<��ܦ�?_�>��]\�V�U�֎�+o�7��Џl&돨����V��|��R 4R�7���
��mA_P	�k���'��ǒ�N(1B'��.S!ɜ��؛����v��.��{�@�של�o�ݬJ�����'���%-�<k>DvAz��ZW������Emdј�����_7s�}�`.��O`��D��=g���0^����enZ�1T��RO|�R�������O�-����w��Z�^^���h $��P�`�0�#�`u�F~��>�)XIq���ѳ�W�\�Ez=9���}�Y�D��p��x����P����
�4b�z�Ί��><,�k%�xW(ˏ�+#n��= ��y�
{�N�|�}m�vBx0�j��3/��:���hxt�X�~;�	�&3�>s�_��7wh*(|��5��r\;c��;XS���YU���۠���Ki�HA��Ֆ�A�h�d,�
�Ǚⷂ����voW��""Bn�xbg=p\Z��
�[JJ
!��G|�aK���}�Uu�qy4]Hz_��x�TC!Y[oD�j.j�l���qz�Opy>^3�>P�b	X:�p����cll�JO��U\(ߋLKx��<մ���S4rn4555tfePB�*/��z���I(я��_�k,X��[?&ϗ�q��&a̫�ZM��w��P7��d�Օq�Ё��Ns�����;+�'��s�kk�OWjgϲ�������^Ū��9��T_�^k����jB�����p�<���[��܌a��ϟo_S5M-,�xx^��gZ	�g�+��\?Zݔ�=�!��{�/�oG�i��~B0&bc+J@�uu?�spL՟�w�׻�����C��~o��@���:��������u�j���Cs����#ŔC�AT~gg'��[+���y(��ƾKNM%�ۼ�HZZ:�ס���3:>[��ׯ6I�	II�;N�,gO�o^O���ޜV�Y�A8W.�VY�+�ܛj���R(������deŁ���p]��dU��]�G�$�F`�t��p�Bs�����k�7��J���\t��q��q�j�C�(k�E��m��3Z^���ˋ��R��!e�%�!hi�n-�y��Ã^x�f�U�p�И�ZB��QE���5�p ��bs��b������w�!x���z�� �db�0|���,���u��D�E�4ld'hi+���k������������mfq���:,�o�^��3��
<"s�yX����/1 ��ǐ�[��y5�P��*��bM��!�XF���9�����
*��Z8��Fip6�6�5��tMm���h��!͵e �G��|��e�!�]�)!�{�E�з�8Yi#fo_�l-�.���~6��G���z#� b�ye�DDN��_�{���_��>�8�zK�,�_��FH�����ɇ\���gV�|EG��<�1���Q	)��H�������v�ɿL�T����e���
���OG�TF*>?�g����=�u�^�+g�{��#����Ys^iRÈ��B����K�Ķ4��BeO}�4�a���y���n,��S����_!Q��
J����B���K:M�f�����]}V� �����.���kk�qg�͵�O;���D����
�4�]A@ HP�Hҫ� RC��(�{G�A��A�� -t��J w�����s����ݜ���}�=�<3����Бk��Ln�Zp=�.旐�/9�oڟ���ƶV����"���2�=��$ߧrNq�9���2w�|w��ר����T��&Ӷ��MR�G7g�{,���gl��W1�X���_%z�"�����-9�`����_^ِkf��;/�s���9B�^i2�,��&�m.��hN
y��2��ry��/��ƫb�L�����o�V.��ug5�"��x�y�m��N��'�)�)���-������az�H��}��Q�Ļr���3Z��̱�g0{��	��*�V�/�u*v�����1�|{�l1��.j�ɠ�.�[�1E��æ���(���$-����=ط����k,4i�||`��3Qi��s����師��B�S�Er&Q��d}rN��	���f@�g���@)[=�?�2�ݿ�&*���+�}��Y\\,"*��j-q��n�%&Ջt`-^��o��W ���7V��ƪ������۾�HZLѰ����B����QO����Se2��><�����h����&���������S��ތ5��Q��P���-�LHi�Q�]ޗ�WA&�3Q��Hr�U([+��<մeҷ����$;�k���X�ys�a�� �b�c�.-�Lh~tݟ�t��)y����]ccc7��c��5������F�P[����~T,k�:�mu�t������[y�|�O�l���]�*�/�b�$�(��Oi�`���q��'^�e��D�-��$�q���Qjt;����`�	�G�؇���s��8H�3aTI?q����`�39�����RBɝ�L�������x��l)���*k�V���ې�O�W��L�e��8�s�K�ɫ���@�S���-(���ȃ�h���O�e$ě%?u�1a��Sv�m�cwĚ��La��X�ZkV���s�p��T��93�::����w���'�m�ȴ�4�������kWW�t���t��'~k#��=��l�cv5���ו��MT���"Sp
QśUo���a��'1�O�=����{Qk���
����7��Y�zEE�~�7a��B�aޑ![gG̈́~Y\���pe,�d��w=F�+m9�l�Oj�3����4X�mxL9�	c�������r�^
��_
���.'�Z��8��������C]{�1�<���7�D������)�Ϋw4����d�,�f�/���씙���H�Iv:.����˟��Lyeanp�⹫���y��+���1�	��je�\}�bO]����g+��Q�Q������5u��b��d��=ςPp+|=v�;S�C9U}��TX�5ex�*kc�~S6Y������W}=��ӭ.eZ���&y�sx�0r���L:�/�(H��U�^+�-�t�h�Vii�?4��(K��>c��(W�����8�ZA:eE����-*.E���3�[�M�z�uk6��d=5��]w��xP{������|�P(�w�t��5twT@�����M9��n���&cuF���ju�Y��0�k�rnM���S>!-��;DF�.˺n��ڻ{�;�5�#����{�u'���S�j�����t"A)L�;��G@�t` ���hű��o���b)��Z��jas�����R�<���5Nt]M�c�y?N���d��2��a+��Ɉ�)�|+��)���ͩ��.���\��lD�Z�[�����'Jy�o�Ve�[[�U}Bm.ȮU��g�^�3�)�f�׈��,����������!�x��ֵ�Ͼ���1��l���P��lױ;>�٩@O�˯'/'.�S7s;%U��1�P��^��c�vD�񭣘��C�˃M�������]�k�,u�o
;aC.J��~<���zÕ���������h� .���(��,ش(zU;`�3J�ZI�U���e�ƴ���{�Q�ՐLk|+A{�C���k��h$=��p������@5��{�p�U�1Z^_�'����KH�k�^teY\�u��P���i�+��g�h�^G���UCT�J��/�k��y)��6�E�'<R�za	��������]T�|Rq�����1o�֑Z��Z��-���%e[)p��#"(����JJ�`�7�u����8F��hx�}{�Z��)9^�"}h�6>�$!+mo�Y8g��l9'&6��\�o,�H��6f�,<ג2S��=�7��!(��������b�T4t�p���޿�O�+y��gf�SU�2U)-�!�NҾF-%�{��2���w����U ��*��H���Zt�|o__�f�'�`ȳݰ�^�������ԴTۣR�m5#7���z�0c��E�8׳�5�ظB~���z\�b!�c�֙a�l�ܖu-6duoxh��d������}G�=7�5E���qs�=ѽ����$7���K������)��/1�,3{e���+�,IIIrb#�m�'%�������i���ui�[;/�Bo����`���ǿ�"�&��f�}��
V��]Z�^8��9|.�sĘ�ƾ�q������m��r��˨��g3���O�v�gEEE��KŚɥ��7=>�W��-J�Fvp<���4q��m�e�\�<:�����A����M>>��s?r���g�E������k��u���Wűz��L�����(��:vj�j��f}@ژ�ԝ�^�E��	:�כ�%&}��!�UUؒ-�ћz���������	�E�O���y�2�F�W�����~ȶؤK]437	����܉�8ڙa�a��p&RD������s«��r�e��1�e������	���Q�<�f*�^�$�S��RRپ>>\����/�/��T�j��+!�|�"����#*-(t�ǚ'��#L#�kx��ƒzx��E�l���z�o�"t�L0��x�gD�&�X#"�jVPPд%$�(�������r��֝�bQAal���/���B�_�6��YT�� ���@��+��
%�1Xz�Cj<׎�Q��R�1� I�e˼�F#�<F�Tvo��f�ƅ_��|���2�-�[C���:E�ׁ����{e�+'��-!�Zl����u���>D�3���P���>]/ 8?�u��7zЇBB��s)�*-!v����i�^:���MuJ{Y���]�"�����x~�4�Т��R'�R~9� ���{Ff�ERR��������?�l�I~}�޼��4�B�*9[�0V�z�U�/�<'�\~���,�R
V.N�|���W�R���ba$S.�|����S�._߲�ކ�s]3��w'+�+�����<h-�4��|��.��gW'��q�7�s�?�p�|4���]��*���2Շ�_K�f��Z���z��h�s뱝ݻ#B�㹕p���l��������1Ny/0G�Z�Nf-�+I��sj,��¥Ug�d�J�l?G�.����,?�wEi)PD�I��ܹ
��mw�v|Qt�y���s7/��0��}���N��«V���弪L\�nf.������o8�Ǔ3Sw�ϫaO������W���mgvTU{���vJ��/���Q�S�Ҫ�2��-_3W[�b����w��V���hu�x�hXr?5"�8pg.��[���e y*������\1�/�4��k%�/#��⾩��}��GĹ�L"��><�]������+��e� �i@
���:���b*��ꇨ���Gbn���(�A6Y��i|�bv���u����A\כ�����*&E���+�q�o��?��r�70h�K<Zl"�GW�KQ�oQ�:C��*Vڟ�1�l{ܰK�.�?#p1ƽɜt>�~�Х��N�&�m�ƮYK�c9'�}a�x�k�A�^'�����~�������.������*Hdff6��qRڇ�y��֛�`�	::��i�Z��m]���X��j����5��0k	��h��L�S�+3�K���n^`��L�7�t���A%l@k�k��V�n��OgZmA�C���l�Z�(�����ȕ�yߕ���α����C>��|����Ze���9�Sq�(��˩���k��P�R^����n��p�@Ս5���KUؙ���>9M���[[�����+@�I_�����w����0\�s��HW������G��G���kp� �'�ؿM^�h������H ����uʝkq�{"�56��$:KMW	]����!a�Ȇ��_G9,�������b�A��X-��=]]k����t���x{ץk�G�a�M�;��G���U�HO�����fC!���C3iǅ���xxy�^���m�A��ee�4M���Ȟ�nd4�m@~eP>h&���t���{K4��>�/t(?��ܽ>H�Lܛ�{}�`�Lf��뛎�<)lt���n��I���z\ߘn&R� ��ܡQ���{�@�b �|��÷�Rls��V]�����f4���
��T	���*���*vZJ��xLCN+|���o)�91��62� űKo�c�K8����W�����F�a�A�m�Ɇ[R�4�(휗+}2� �*��M^+��n9<˯��Vڗq�%_��y�uq݈K/F k�D�C֋����}%�xȒ���o���eGgqX��B���W����y��Oţ/�Z�g �އl��K@�&Ox������xT^ʗ+8^��������s��zc���X6�%���P�Z�	��Ǘ�\����@H?��g��\H��\��s���L������_by�����g��t-1R(Y����R�4�m�y;��8���㸼�V�����r=�v��TO)=���6�X��\��*x8���n�cd{�۸�O����9S�4��@!7H�MG����i>{�\vM���]���u�ܶ9�5E��jk{{��JN���Ae��)�fq�Z�x��[B	le���۸�IN=�+V��x!�CA�*ЦJ�w�{�6�s�w7�-��ͬ|�%	�VLMq��4�(j��U�1�95;�ۈtť��+C��E�'���/7���Y�y%�Z3n�c���:��
9���ٳ�T�j�q�h����}���r�ͣ�!1��d�����Z���8�?���%�4All[���
�=6�����W�8�}<��4��Y�φ��s�;2�یL򳒲��P���ɺi�_�.�3&~�g���>���4a�	��_΍�\����<�'%%e6ό07��ݽ1]8Z�O�T�`V��ds��Ƿ/�)����/(Z#�e�	�x1�����c�N��r�Of� vP&�&Y���r-�_y�Ʊ؄	*X5Fڰ���|D�$O?�΄0��b+%%�����R]Ĵ]�3�h�ƈU��I0#��{ǘ+������݄���o�Ĕ��l��M"i����ʼ�X����n��:H!(��|׸�B�a�Uj����&����N����[����AK4�\�f�_�#����S����;|��w)���+5�;2�<)��Zj�>����\8�F���������KVψ�
�N�*!]f��g�V8L��Vm�z�&�$N��Qg�-�A	)9���dN�Q�-�>	��S��g^�/[�r�sȋ���8��l7)�!�^|��� [��$�y.�CU�~��}�V|�Q@��!��xГ*�|g�ۂy�ש�~6daA�H(;ؕ3��W�Yf��+7;y.,�Ը82�S�>�z#_0ao���'�N�V�?PXd�&�S�;x9��i����m����m�HI��}�Q�_JI9@�+[��/bS鱕���O�KY�|0|n���W:�]ٵ&<L�����[#E-��3��ɋ��J�s�"�Bl�GӍ�_�����>�)�=��� �Ƙ����r�k�#Oó�KVX�B��.����>��I	�����X NQ����b
����
���ι�g��'��pn�.E��,���u�����-�ԍ6�]ʲ͆��/���Tn7ݑ�w�t�L����r_&������Sz4SR�ϟ��;:~����B����GS��S�z��?��oI4�m-�QLwA P�������*>��`Q���~ 
v��0�E��0�B�J(:��}󿛬����{�,��W�ڳ���0Y���p�������>��	tC򆤸����ԃR`i)���5II���AOP���������D������E 9�c �	���99�:�A
�f/����l�y�tt7U�=r���yz�����9ہ��X�����KJ~_�JdD�20{{���W�����o�玗��#������I)9�6� ���8���>0/89IU����� }����&��4�tU�Tl#�PK   ��!Y?S��� 2� /   images/99226213-8268-43da-ade8-d9d07cfcec9f.png�gP�Y�6�3�3
(���J�80�d$g��AR��!I�,y�$9i����LJ݄&������y���s��rW98���k�u�k]k�C���.�\B d2O�VA H���$��̓�_~u��Q#�7��+��w|��@�� ���f��
|󆋔�������DrX��8�<w4�pp�Hŉ� �2��架������ge8p����9~�����9~�����9~�����9����D�a �6a����s�?���s�?���s�?���s��W��
?���|���t�+�p�����q��ds���,�r3�A���7��vaj�(��%'�	�ψk���XRKj�^ی�����~��Gz�޼nq�"�s�lz�c��*'��B���G��*����'�t�����Ð����9~�����9~���Fy\G!�~���AN{�8�֤�M�,�-�U���0/��w�Dd�-�h/j�`��z���L��qe%eP�Td6�`�$!{+m��+�H�0/0�EV\&.1����2wV�6Rer��t��=	���n8X|��^�V����ϕ���-¯%> 6#�
{q�$-��6ﺴGDW`�3�O�5wr�~�;�VNYv���.�7N''kg���}��:�w4&vy
|�4;�k��:�[�$���L�Su��u�w�4���Yz�+�,$d1<�nە��f�=*�����o-;+�s߾k9�����#����0I3��\�#n�-�1�i2E�=�]KeS�g�~Q���z?K\���N}��N.'�M��x)~M�銶w�����2�-#�z!C�܁�����k�U�<K���5,Oz-�e"l�k�xͦ�ٻ��Ǐ�U2�+u�D��uLǭ?U����{3Go}�5$H��67�Ck�g0܆�����<�s���?H�&�����i��rJ=��k���p��ҁ�Ɇ߿Q!aYP+ڭ�ұc�����X�."ί�b��$��f�@�ى�a>�[O��w ��[� _7+�����~g�EG�+�}X��$�qf��q�VB�<��C�����B�o����Y�xj������g�bh����>�ޓ�̧NLPK���ߨq�nd�����B�[F,���O����o��)<�j3����J�-�}^3�S����q�o�'<}'�0M�F��`7�bqmwi���~3��քQ���dFK[XQ�����5����b&��-wd����^H8c�V�g=m$�,�l~��"\D������ӕ-��/Cny6�*�)�O�|�����8�??~ZK��ɳ����[rm�2�#i_j>���1wY��l�[8W.5���P��D#熆�L<������"����Q]��]s��蕄\�y"���;�˰��G�v$��T��Zۭ*H_ݥ��<�>�e�g���P~8FoY"4���i�ɚ
�29�
��g�'٘,�����%|�}��ݙ�F�k&�{ټ
/���\�.���� B�v�ώwt�m.���v���2Ln�E;�3&�e��Y�zDU0�GѷX��R�޺f�&�]0x�;S��>	,	M;R�v�-�)�Z?3����Q��Hs��H����
�y�٩3摝je��4���%{c��E�[::4j���T�/��~)0���o lC�{�݌$O�4{!0uUe���1c6�s��a]�Z�~{0�X�����,��M�4-�F���z����;�N<"O�?�4�q��|�ɗ��Z�+у���[��*�������^�Q7�~����w�㔭�S'����:�X�,�����������K�b/~0
آ����nXn��z><Sj*<�Ij���}{��J��⃖��.���C�\�r�J�l��2�|�-5��u�I�>6k:��y`޸?-3��׺8;K�{�H��d���A���G˝�����ȩ>�ZhO4�h!5n]b�ݫ���R�4�W<+�Ej��7i��BS9n��;xZ%�	?�8 s�<n�%̝oz���(��-��J��/��jX7Z�����(i �_N��Z�û����y�soձ1w�7������2UOZH�N�-�Z�G�(6���oEuE'�pu0�*�S?�=_B����"�/FW=����ټ�*x'D}�}�6�
�����u�:�j��:�lГH7���3Hk��?V{�X�pEn9p�-g1���a �������5��!S'�[ԗ��<`uy��mZ����ݣ�<n�LKǳb��c��`Y�4=�t��?�����>n�~=�-?�1	�/s`|��R���x�g��i[k�����h����__�J�U:ڀ�z�L܃��._{�(�%'^�� �N�c�e�ڔ>���©��3p�B;�,����L�:6h�z���"�Qy�*��hu7r+�Z���y�6��s���Rv����Մ��eܹn���Y�ۏ&�>��[M�L�T	8��J��q>�x�%�ɦ�lx;��ƙY� �ZR�pf�u=wR>�:	��l\�����������(����`!�x����s�Z5� _*�ȩ��@�a�=v�0]��0�-�7�;��ձ�i�&�6_���<�Ik+����>fͨ��ѵ�N0CBK��R��J���j�u�X�N����{���R�6��t����`�g	nK�3rT]ݝ��B��6�|1��`Ba����9Ob9o4Bz�5b�V>3�s� �8	�c{7?�� ύ�b��.�l�*_����N�6�~?y���nTy�/~�8,'i<#��Q�n)��������h��ܖ���7��}��c�:z{��$6N�����:���g7ŎU4���4�}	M�M��f�5�����S��+��pz�e�� 9��BEؑ��#�*@hL�N��o���M'���E�e��h��$����0!���d����}) n�+�~�D�is�=`x�� ���q��$ bƱb��4���/9�0��������`6�������e-w��俀��� Ä1Koc�r�o�v�T"5>������?v� @(zP,{��9�/Yw9f�k�:ͭ�V��H�}��9�Y�o9Z�t��=� ��q ���[}�0
)���|���� X�E�������ѵ������M���Av, +J�X�<>��zFk`jF!(o�ӻ�U_;�����6}�`�p�=�5��e��������؊w���ǡ�����&����'W�Yɚ�HI�:r�������������Իk�oR�k�[	lJXN(a݃���-�������_<V��(��Ow�f�b��g~���ٗ�޷o�h��j�����铆�R�+k���)E��0�GwU׫��<�ݹ���Yh���.Gu>gx��l/���u��j�$y��h�����S�gE D������i@�V,�(��8,=be)���]i_Q�˸��|�FO�������1��U\�>ơ6t,��<;]�i���C�&?z~>%f����V�_���x�f+�,�`�����A`%���Iك~�llZ(/4��\g*�}�~�a]#�1�IK�
�o�z��bAz����P���}ε��1IŠEUUt��1:���0�{Ӿb�=�N��@��[������^4�7r�?H8qpߺ�yZ������s����~�y.�~�y�h� ���!~�2���0�����a&P�so�!l�;qp5	�RPW�hN�>���Bad4ڴ�h4�%ho��r�Ǔ~�}��ܼA������~NGǉi�_x��	C�����  �n"���P��;�Y�th�ԉ����M�!s��y[�y� ��2ǬK���CKF�4�f���ɾ
/��Ryp�`���t���!3��z�{F�Q\�[o�h�(�A��&@�h�*��E����U\��Hvѫ��Qx��0W���z��7!��$t��2���,�mO�����xj�ǋ���p��q=��_��7j�
���S� b��o����@�[�_j��(o8Z�W1 ?"�4#��ɉ	�)�Y��E��<��f>͝�M(-���}����E]u����&�j>��b�}�h�`�r��*� ���~�
dG[���s����'{k�����hvPO��L��_����/z��O�	��wK�D0�P\R����=S*���Mx�vh1C�cܑ��U������z �
 ���Wx����ܽ��aGn�s
��P� �����@���Z1��{x���+.~0>�[ ���큖Ԝ�jWGwynˏYC���ì+��֎������<����jEmX^�J�����d!�kEE-��������A~QD8F���İw�&~�p.��B�� jͬx��� q��E2�@S���Z� q�1sv�t���+,m�@���l~�5{�R|��� U@|��40?��m������F�O��f���:���pi��+0G����$`�ׂ��g���Ϋ���>R�Y�U_���om�MT�xy���]��;=;+�� %Y0fqiCܱ�>A����V�<��P��3�7�mf��w����pg��j�@�i���a��R|�R�0����hh�2�����_w��f����������Oq
A�j�a{l��������}PB�~`w�>��&��(��R}þ�E����o�9�X m%�s+�F�����ڽ���%q`�y���S����9�$����i/F0U��g{���O=�٣�;�^a��SBR�pt�cݛ �d���[����ef9�KA�v
��\��|�̜$�JN��N~u|�k���\�6�d�/�1fTpxog�2���?���'0]��z_[hId�߯:K!\����%8����}|/��FV ��((�~��rV�ӓʏ�x1�A�ܪq�ַ��Ԕy����� J��R�eT��m�~�ǡl����D8��\ЃY���}����;9��}�rR�ܷRR	3ƒmͧ{��8� �(��*��XD��b��2K��z�
���ݵuK˃�)�Qî~ȩ�PNh���M�,)e4��+����gp�X.xtd"��U�gS�xmخ���%Ey����ۇ����ع�����)c@��r�?{�TlH���Fn�U8CFf���������!w��|#���(p�7�x�b��6�ii��}6����b��?tG��g�K�R3+�or� ?d�G^��2�e'}5��Yb���s��+�_������5��ܤDV9�P�ׯ����^�

��3��ׄ!Tφ@A{5�E]S_EP��GH�l��%��a�y� ��#���L��RT�-�X2$ز�L�ҧg��Z9m���D�\�J�+�rO�ijJ����I>-��y֕R��1�#��s��j�"�饻�FoP��9�*e�F��{}O&vd�ؖ���] ���<a�%'���FFJ|#(��\���-���XcU
�{m�.|�Fn��@���:`;��߂!�:�$��I��-����{�	�+BQ*%O{��N��d}��K	�����(��r�������}��`���6B'��rV�FYv�w-u��adх����ވ}F:&9"R?��@];�X���rb�SW��>��'h���Us��M6��i!Q��oS{9ʖ������?,rUPȴ_YK��Q�QZ�����ҽ��d�cc	2��]�ZZ*		�q��^�k#>�xlE'�
��TyN�����_�?[U�ЄL|�ܷ�����Рd��1C�^�J ��8�(#77��W��1�G�`"H�^os�>������_M}WW!�ӗ�֫���Q��1�Y�gUl9�_=$Z�,�XJ���Bh�>P7hM�$)~JF&=��(���`=���ֈN2��8:8`���_�v�xˁ���]RD�;;;�����bL8ʇ���^�N��[X�����d\�DaC#�:Ϝ����Z_��{t�w���I`u.@f�9J���Q�jk�?G[�܃�»�49]�����­��Nc��FCO�]��I A0�N;i<����KV6k�$��%�.�<���:��==������*��pGx\-�w��G��v�fE�#%2TTb�����7������A1M������ڊ�ܗPE���͈]?�'��B��hg_{ܓ67��V6��/߃\^��� >��zm�D9�̮]Y�3K������?f�f��9Ɠ��-��M~g���_5�l-#� 4���lA��ʸհdc�m2��h��"��ۛ�)�j������z)<�>'��)��K�anD	U�_A�g5�!8W �F	g���'MZM�vy��@���5"���9I�/0�;ux۬�.����A�N�*Ha��46�M��<90�QZ���_��k����y��mv
MoO��t��ׯ�+�˼?R���w7&&���\��}W��2�
�E
�I�Y���zC�Vq8�VO��z:III�+/��v���|y�}�.�2(u�٭[�~:L<�R��%��5����$�&�f d�@}����A�q���~��a"��b߬f�+K�U��S��t"��LU���Ch����2Y����:xP7�op��ܑ����?��k���$~6RH|(v3��7�~��s����0u��8D�T�M�Q=��7����}����ct��is����F�\��h�_xG�u�<07W&+�H 6�ZI9T�V[-��8��kO���"@��(�LN=���C3zCqPgHb�+)1�\�輏����}�>��v��0~ܚK
rzg��%%>�f7*2==�i�N�8\��5���?;M0���Wa�B�_u_M�/Xgm{�^]���<�<���ֻy��綩.�g-��R����oH����? � 4����j�I�l�����8���1����m�\T�q>�gk�01-1[����������z��%(����s^�d}�<=�����8`��XPK)��O�GEP�,�A���/��mis��;���k#=��E/�]lJMO�̮�0��m(�uA��:%���;��I��o=��0Fo����7��������� @�t��Vx�,��g&����<��.d���yVOSRn�Jk))�'�cHS�{�r����u��&[�{=���3WI��.�`D񵋬 p��'']��WM���kyz!n-|��E���^�sJ�X��.%���NP6�h-c�(���$mm�qY���ujj�е�������1f.i �[ix������N���1	�����v�w�c\GO���0̟w�)rߙ���W8�M�������:)�q��- �s ÈL��V�?J[��Ɛ-��蘘��'u�ZxV�1���c�Ų��t���3�e9�J��� ���*k�,���pt���:�
h#,|�v�r�[[3$qq�]��}��\�n����oԋ�pT�A�対��]�f�5A,&"�a`>S�!������x�!��w�uX�&�@vq��5sߠ=v|��� "l��q|_�[�?^�Tt�1fخ��K���Jyh�@$����<
��,|ji}�������F�`�^⯰��w������H�A1tt�+}c?V��Q?��'px7X�5ޕ�h�o��DN2~�8��2%%4��������f�A����i�!(��
u $��SR��tt|�����C�!�Z@/�o+�{�i���hbR&'�(
�e��қ�1�̋\S��$9#J���*�:��P�J�P��\�h��\�2�u�Jaa^lT�.�p�a�� )���f4����W��ǝ�� L���ό�z� ˤM`rI�?o�XWg��}����Ȕ���"��'�3��VT�kZzh�Ǟ�.ZP,�_��U�ЧOd2Y_�C���jh�f���z��!䏆�}�nI������P�#Z{(c���������b0�@�bv{go�8?��~DD�ݾ�Bx�,ϴS]\�_�M7�w)Bk�MV������=>	�����ק���6)�q����o�����v{�Lg'����Xk�
�����?�ne8��M�K�n��Dw&9"�LBK�2Bc1;�ާ���ʐ��3t0ם�B��n@e�**`�RS<�A<o��$�����1����W�I;��V�_�pp�((�ο{�A�w�6B&���ق���V�����*�Бf�]w���♹�0���V��f��jN��:�z��Ʉ�Z��m��l<���_���X�^���ʰ�o�Txl�Vj�-`���xg��ηe��8�����m]�@���6�_����Ԕ>lb���mH�hV[�44���Ԅ�)R�y���L7�܂��(�w�A��bP�T��b[*^dL��+烲��ꊠ���̟\���C�&&W��RdL��Í��0�F��uV]{9 �^V�~~-��E:�
Sz\]N�G3D}�,�jkڬ���Z�?qssu����0{j�(e.N�����a�`�+?���:�R��cN�����g���,~���FQ8�io%G����u9��F8�h9����е��Y�t��qպ
5��c5���S��oߐ�a��J'>�i��Q��jZ{�"&�j,����|�������@g�����K��%����$PZ��lE��Q��O��M�`�(�����11���}��4�V��0�x �s?jC~�E���*�@tԙާJX� Xu�:��=�:���΍��X&���s_nnL�R>�XB�,~�r��Iw-�����O$�6�h�ր��Q��F�皺�)�}�ߟ���������-Q?yr�P���X���51��Мm�u��#ynh�V�Ųk���c͆៌���4���x&��Dz0�G⳰��q��I]]�T��F%� (��N׷Dh�hB��<����h����\

�)OQ�s��������LK�ӣ��p/pL�&�U��V]�m�� ��a�� �S4M�[˓��4��8KT*�4g�U�=��s+&*�Ã-6Z����6mw��(����Oc��n��89y��'$AN��������7q���;��T� #��c����V�/ϟ3�3>h���Ş���#7�{+���_��� ,rjKv�wP8�_jjR��kI���K C���I��z��Z(��wuq�gap��G$-A�I��c���śx���@��׵u��Ζ�^%8)o�K�L��`�z"#O}��Go��)\�li�[�����Y
��Xik��JFn��--7�5����E��pt��]_w�Q�~NT�^)�w�'��؄K�� b��h��j]���͖0���=��Hv9���K6a��k�K����4�j��JKҪ,����eg����s�y�����Ѡ;�ɨ�'�z�i�x����0nϛ��b!�l���-m/�.���D��2CBs'X#�X��;���p�Ç����BIC�9kXY���˝z�M�JI�xQv��D����5�T�[IA�%:���B�l�A�F����A]!�zNR71���R�������z��*M�.O_��Ћ@��im5������h�jg�e
?6f�5�Ɓ�m��������}�$��#�r�Jˎk�]_~����WRD��g{��wvFs���㷁 �|��!mk��/���0Җ��q"��E��G�3�Jx8n�+��_�N�uaH�4��ڕi/�[0�T��&A�S� �0�GR2S�܂bKE�6�t�~=j�%P�90+Kek��tHH��"qyy�.n�K'��YpG�F�b"@ߊ߸y�#��{=�k,�']E�ȴPe���"�������h+�.���"q8�-�7n�fXXZ_��y"mHZ+�����L��vF�5g{�Q)�ʤK67?�%���%(9�i��?/�B������3���А
R��S��)#�����m�^\҅|9�X�{_�P[�ۉӒ��Z|�U5w=�1l|0;����/W�c>؞�-M����7*"n�M��h�T�1�,.r2r��/�X�Ud?*)��P��S��'  ����~��e4ZI�e�������h����sIL�5@1�y�p��6��l�;�K��ixu7���߉t�*,tbz,�D�d/]A�n��&Y��\��\��)G�e��Eʏ�2V��c[�U]�����ڭG-�,(ߺ�D}��,�"�2+�����BMM�x۱͗@oM�		�ٯ`�����-�IK;i25�_����;�(_��u�f�dѵB81u;������p�CY��9jN­wH��1 Z���|Z�O��@�L
��q��x(4����h�p���,"qgU���u ��9��h��~`g?�T[ۜ5�P��< ���/���d�*�u˿C���?��gW����^��q/����\9��HJG�;��ejlx�		0DF2X\�p��Z4�e��
��Ϯ�L�_bT4� �h�$��l9�X�*�B��И�
*�Е�į�8�fnvvН�Cz�-=lI$���dm����{�e��M�
�M#f�k��X��p�z�x/�u.8g�
�����AIO!)��T�č�Zff��y'��܁D'�x⋲���iQZ^u����������sq�	�Ѕ�v|�wr���M0r;�(��}�����z�:K|Hp%k�[� �;q�|�1�>.]\�$4t|תʲַBSh�vXL���b��Ћ���\ˊJ<��
M�ſ-����>��3	ڞϩne&�������i>ܛ$>CfP��d�_��Q���Z@�s�?�����Dc*F�[k�.\�{hx7���u��:�l�+����i0�qK���(���v�3�4W���N�I
�M����]]�=�M��"�`ՙ���b<^�86F���j�*��r�N�Ec^;�����(���Տ]����<�#Ǒ��;���n�&2j��V�5gKc��Á�(̇�[t���T7���2F`.d�/���ė�O�a�	1j��>�L�}s6�mss��F|����i���Q��1r�( >����g��鍉/�'.�;T������2`ND��)�(�eF~(4T��L/?YHIq��p�6Y'W��$�{]���ϯ��`�#G�Ǎx���2�m��!��~�9�r��҆�թ�MFɬ/P�i�����bԨ Uj**�����_u}��ыJ����>F�4{�)9}��P����4����ќ:�����X#�]1�CR�wa�UW�-z;3����|"i@_��DI���Xr��B��U�B��.����;�z�;��A~�ݷK��%i�6���T8�����:X��x�=��4�i��Q?�Bݬ|�>�@��h���֭3ۆ�/�i�ߦ�_�>hR�H��'>�W��XK˛k�ܮ��ZZ����������X�5��2�k�vq�$b�e�"Ū��l��PUG{c��l�k�Cӊ {� ��n�4J(*L�vu;�^�G���Zd�" 8.9x��V���FD�C-���j�C�@&��l��J�M*+5��k�9�i�.�e<�!QQe��;C�h}ԉX^/�E��ep��E)��G~�j�n��j6�����O}̎��San�q����O�$�
(o6#.zz�����bNX��[���M�l�ll�@���s|i|ӑ
E<kKZS�M��ׄ��<36�[�O \�Lf�X�h����_C�_���X&��,��ǒ�.�FƛOa���a�{�OU1/���7�@{x�OSAM�Q��w`�����5�k�AA�J������>!�4�qF7��$� ���t
Ž����)�_�� �܃+k�q�='��R4�kr���	^m��[5�,
�|��3/��#�E��wI8表~��1���.�(�'67���
�}v+#�J��S��Ђ��0��z����T��g	�\��?���{��x;��V@g*��1���`�dC��k3�J���CG�$a�'�Z]�����Eig��P�>JRP~������.��QM���|��fa@��Ȼ>^Y�6����� a�&'�����[���p[��"�Q�7+{�ui�kC�|6袵��Lm1��P�⶗e섆׸Y%��* !_D0���/�oZZ� ��]N���Jq�e�Ǹ�k����Zi��b|���:;-/�O����������]�^����DA��?�V�����d~~q���¢�t;R�-�`��%y����QH���.�qʌ���6�鋵.3EG%^��c���$������O%$,^�1�!
�T"x/ܟ��ΞYT����; '��hJ���#%�8�]@�G�j0��82�+%2��U����h�˴�@>L�lĠ��m�0��T���B�}�6�ݕ��@����ԙ�k���m!r2$��������k��0:L�B�����A&`t��sV���l7 .�_��*��"I�+M���N����&j~��ϫ+CT	V�����F	BN	�@8��S0N��)���<�h?	`��[ b@x�>,����_=���	v�1x��e&���k�}�_Y^�b p�*�g}l����y������,@zl�9p���D�'&�$�&	;�gxه����:��NWAD^��!��wMG�Ga���̇�x2��K��X�f�� "ˣ ii��[�-O�M,pB�e��F+ˋ���Ê
�����P$5��N�v�U:U�['�}ț@��e�����+\Ζ��wL><j��A����tt�A �<��<��6��a#}�۬�3(�-+�ҷ������kkׄ��)�O�lA��NMk&�͓\���L%H��k���=9��u��O]YQH��ڠ��d=�%b�a��r8��(�N2<u�\n��J�{���� ���`W�Mn![:<��^�IlW��w`�'��ޏf�wu�^�g�0�w���(�3:���p�iy07�	��Z5CO+��^C��("�7������DS�:	�Q�Z=n���$l����E0�(lʰ�44����P���-k|�v/ņ��Z��)��Cl���f	�!:-ϒ�}ך�����m��M.�׀vJ���V� �g��������O��I�t��cq��\�fIHI�q�����-I�c�#��4�4v@�_�+*��A'z���fK<�k�a�{.)�N.�0S��1iP������@��<��Z��u"�pӧXX'Z�e���,$�]q�L�Rݥ�V�u��[7[`I�\i}��#��$FF2��\���K�`����N��xp*.*��w7����?}"]�0��X8�+�{�t�<{�,F�t`��l]Mʳ��?��Dm������M�<�
֮h�<��>���_R$G;}<�َ�ш~M'���}���}yAi�,׊FBw�I�̣��e��O
��VL�m��Q�����'-~dS�N��t��uOο
��j���r!�	���t'�7�}N]�GU�����o�7��mnZ�W�����2���3���%���ʭ[��s����L@�h�)��͌��[�>�O^�1�!��AI`�9!��d _�[��V�s��_'ײp`,gc�礯/,�kğ7d�=�%���OC�K�����蕾�$���w��sUnѰ�{�S�)ނ}�x����8j��|�;���a,)�m�m����I)�=1X��N��������%�=�5�<�B'�b𣞫 �*����H�
6l���G����#��8�Y�x��h���9MQ�Q �D'�Q�~R��?�ctW�b^v }	k�9����Çɾ���{J���A'�G������|J�y'w������W�_贮��(h����`g	)(��.���
ߏ�Y[.�v�����	��~4���$%K��ߡ���y�,
�k�/�ΩU��ԍ���-�MA��gB�U ��*���
�Z[�$����*z�	���g��������@d!�s:�9J�Xٛ�����R#�S"@S���E_�n��+��NH\Gt3���z��ʧL��r��q�Qt� zj�u�=�:�&�6|��f�J�֑��(��{��PuM�w�ѯ2�(��8s�W�py��	�$	�ߴ>��Z�b��Ǹ��*@z<*�����rr����x�^7t��<��Q�}�/��)��o����]�q[�7Wl�����Z/{
���F��{��[_J��>  �#�N�%$����C�#��*JI5�/�w�K³���;	��mp~��#H�If�꿠���P���|��4�TUf�'@�T�mI�3|���(��Gu�������4Y��7�����&0H'�n����H�]Mqz��,
���Q�IuQ��@,�C,V�e��W���JȾTT=�b��@� �FQ�};�����Zd������Kqv��-L��$}�w���2V��_���4/{�aRC��xYZ��X�%�q����J�ͳ�!1GM���K�*F��I��;Y���2�i)N"����둯9`�g�݃/-f{�T�}�����hj��U)Wע�JK�lN��ᗾ5m��A�)x+�#[ڏ�����#���5٠'�����_�9Վ3>x����O`()5X^��t�g~E=��s��l��p[�"y��Hk�4������B�]�0R�}$~|L��  ���~�~����4w�)�Xָ=�Va�!�^^��#���}дG`.ɔ0zlu���ǿ('�m���3m����D���f1�7?t�T� ��i/M Q�ꞝu-h� �Z���\�,��a��M����u�8��i�pt���Xt�ũ�J��5�nA~s�:+�_f��!���l��� �Y�I�\���.�,�z�ɪ�����o��d��;2´"�ߌ%P��{���IlR�!���<k:8���XE����4�~!]�g���5��yd�L%�����-��]��w�{��(g��_2�U�e���E����~t�קaa�}Z��/2����v�W�g�Pńw��x�{X��Tw�{�@�U3_%]���$�j���9���_a���\�UAM��ў�!h�O��1�"�C�g��|=�{/	s%O��/�U���������XŤ=�����.���4�4�VR-���h�%� ��+˜�&��;��^�Wx�L>�e��Q�5<vH�fB,] �����;t�a<���P�R�*��z���C�(^��89���8�(B[�	?�C�zY�o
��=/c�"t�?�t�+[����ɲ���>�2��|��I��r��;N��{(}���|м�0yeC����n�%h7�!�dkLn!�%N�Z�	aL��,���EB��Wmu'䒄�Sx��M]>��g�g�NN����� P��������ꊕ���ԏ��H-�����fろL��E�=΍���p'�i�H�VR�������T��'wsN��7���٧�DA��%�������@Cq"��İ�YQ���� �=ݙ�e[�Ԩ�7]ب(ttQ�nH��LJޟu���Xzf�~@0��.��I?Z�}��ӭ!��Β#B����޵�t	�j��Bt��>�W�����Ԓp6�x�8�Z3����7H�\��c.�&J����,�Qh겳׮�D,v���u�O�$�6�����$z����={v��*��א��	h��$�w�f �t��,��_����ٍp�ٟc�K��L��0vp��T�. N+���m�]�{� ���m�'���q�h^�.:��/F�k�!_9�)"�I���H�J��ϟ_2�:l����o� �/^��^i���;1�j�>�=��6�K�Dr�.$0>m���;�	,6��<2;??�Ț�!���׷�͸�o�����;l������x�����㳝#�\ۏ��S�����^��R��>�L�nj��#ܜ�:�?-h-���)a��v&\���K[ŞJ���O���xɀ%�Z��?���cw�X�|�4��O�4�vh:��EUS
�zϵ����
4�{�X����������� @�S�`�)Ǹh&�z�.�����O��Ӝ`�l�FL���i2�Ny���y��F�21��Z{׌��㨕�Ќ�i��˵�ҙ�".���e��E�(�]\��@��+ ��\�T�RxKk�+�#�dZ�+k�<}���p���%)t�)���P��g|��#���	���ieg���O�+�`&�[k�*)�Vgd�k���w��|~OD�w��5��n����5�OP6 N~#���K�(���3���/R���.k�juI"����8Y��.��C�ss�����ș��2�J��	.�a|��;#B��m����B���dL��u<6�wK�z�yHē�*�&��L�����~o=y͕ܸ������x��~�Z`�Pp�o%��V��%�~8�Нm�[4\h-��kp�*�9���ص60�����闱��G8�aDD %�[���Z���(Ι���s>��y��+�.�����(q˯��oEv��d�]��(w/���{��{>��9�+@��tgK�9mX��ɞ�e��ޟ�/�{�O��|v��q��Y�9��nm�\~�{"���)"���|nO>?<��vz�����*�M�z��X�ޏs�݊�ޠ���@��gy��I8Ԥ�*_Z��Nl��y𜻢��g��Hj�(7C��x���&p�b�M�no�i&�Qi[�g@�/��0+8�qh��dٚ70�~~���p��+]����]�>�,	�\++�Rj���Yߞ�c�4���n�����f�8׶H��������Kw�.gYVWq��<2p��3��^v��K<�����|���C0�{$NZ_���$Tq���{I�@����ڬ���%/��@k��&j0�ss����5h5�ݴ��Ao�͹�ϙbQ�Jt��wF\�b��7��DӅ�!��`�R�fg�m���>��+����a፝��̸d����;�a��K>̅V�����ӣ2MT*�{	Y�����Y	��W���@<�cC���[ݎ��V��w�;���9b��
�E�%i��/��s��i�~oRW3�+�[�ML2�w���{���#̖��д���д=ר� �E��NDu�sV���ϪF�)~�_w��>����nH��>:&I@�$FG�UuC|��!J0���@����GS�o.\�鿨�h�Tij��{��F_���+BA���2��}!��U3��2}���_&�^�.:R��;9���i��L ��=;%e}�n�K*�{�ueŝ��΃e�:�ϕ��ؔi���d{{{U�77��@�'��{�B��ZU��Z��T�*iE����B���{Qt�l�]-L\�R?�a��<?�ɾ�b��s>����~`n�2_���-����y�(ߔ���6I�Ͷ"�i�+.qpH���A�!d�U� 1q�ư����qO`ڛ���B�9�z������N���[���/7�+���иDv�!e� �|�x���+�j��_g�̸z�;���xn6�@W��^�@�Add�a�u�"���2⿸n��!�%�c�0����,�]���^�T�I�T�`֏���)�\��@z싈L��6=�-��H�<wmm]�-�����O���x��֖薨��'XAԻ����-��'�s/��<�dC裹g�g�v��'�
Y22/�ڻ�<=�
��J?7�����w~k%O��77�Y��y�S��ŵ|�{��g��9�WQ1@!���}����"7\\�������CsN�CsJ�w�H�&;@v��J��x �1%dc[l�2��g�Nb�&�!��2�#&t���R���V�'�ÎC��v��� �U��Q�Q�뇱�����}N8�����¨(��?�L��J{��dS����F�^�+XbH5S��R��V�H^bJ�Y��/�a\ŧ�l�A�\�w�	�P��z�O�A,�K1����2���F"H4��.�D!�5r��,'�}X~W�ʜ7�r����ωJv�Ƣã��y&�Q��g���ggA��
 ����I6%v=Bpm$h(�~F��"pc��ɧ����VB�=���y�4R�d&#~�"UX�8�ʃ8a�&�T�ʺ}�</x!ax�,��-���@�YTb9�t���U ���;�����r	�^DIADE:E�KP��[)��V��ne�ai�.�����g����8<��33�}�=��y�O�|��,�k'	���P�T���{f���ec�{�ʏHD��*�/��X\��uH�%���ү^���Yȕ;��G�3��R���j�=sPr�B�]�{泛S����
��<+�$�����^���F���O��4�Ź�&C�\1���с����Ξ�O��m+Xl�����(�:��ڝ�GW���.Pvo��yR��p5'��:b�_Y�@O*p��Du��Nt1��"ՙXP���f�'��p�bvy��EF�D�*����w�?����!Z����!�̽�e5�h�z���&T�]���R��ThLR�9�X 7�����l�����NC/nq�i!�u�O,K�K�+�urf��vk81�ʄO־���#�Q��ږ��9�u�0�X�s�]NW�y���U�p���rIx%�b�	�\�B`� �E��ilS���H��Lޤ]<����h)�kf��?���<�e:@��U�紜���u��:�����7ׇ����.	��?^�r������c�G�۳Y�[��Im	j�c�Mv_���k��iV�HP����v����_�:Z�';�����L��=�C�v,�D�`�����`.�PR�h)+IzY#��p���|ՙ/�1`�bl���՞��rX��<
�xJ���וH�r9�@
�9��Z��-�X��6���i��mP���Ik�D}�]�onu��AU�X���^��S`�{R�n��<�澁��R�7a}���~�+a��k��!�v��1*_�vKn�T��>d7���Tn�}sbA,�%yj��T�!�`sݖ.c��nL2t�w`ʢ/�F��#f8,A����n���=j��z(.��v���:�J�͆rqm�V�� R�;6���他�
��Գ�_�����v�N�\
���$�[��h��";���[V]>?�����1�J�N�?��/G�+��2��`��vw�+*":������w8�y2����zh]'�nWex�Ӂ�s�o��"�-A�%�jC���
]�x:D�2ER��^;�Y%������Y�8)w�ʷ w1=�W�������W7�b��`��Wx�b�vw��_����$�V�*�=H���>dp�3n^ǎ��������xNg֍]Ѩ6,��G=��XM�g�|�@R`�&�#�������*|i��%��P1��P:�0�̧�VC8d}_����%w/o.�}��6�\��"h:X=�_B�6�4#H�b��x֡�!��$�p=S�<�QC�А\��>翻 ��R^�sv�A��{��C����c����R;�����Nj�&̐wpwޙ+���o{�5��$�e��:��qK�9o�8�L�'_rC�|?teJ=1R}[�\�QE�f�7?�j9���V���AJ�ȝ�Ro�T`]��D[�uĖ��Ỹ�����(uv�7�'��-�w[Ìg�*��L��A~�L23#p�����ٛ�:�$!#�Q�t���f>�P�ce���:n�R��uH�Ҩi�M#-�)?�_a���3>��r�.����$�н���3�y��F��$p+]Q:E��	�_��6�^h2Y������B��
�f��S�O=��%�v��T�.�����l,�'������M0�͕n�^�&pX���[ ��
�eʿ�`%���ҥxJ3u�֏���+�R�I\�߆2�bѹqDn�܃G��~����S�p��#���jSH��>N .T��+������~��?�U���Zæ�X��HI"`-�?ɐ��XHov��i�"���AoT����UЩĬcUSw�+Y ��q���eN�� )E2R{���ϟ���gu�_��\h~�(��(n/<�:��Q}����� oԕ���^iW�_���)��S���=�>A SR��ʼO�r�0�?���+ʚ��ߺJ��n7�oq <+PU�P�,cN%b,�*��\�8��ܜ!_��l�µ������<��;�l�����c��_���V��y:�$�^�ٟ���`�(?�n����9>9��6����k@A�SjkJKk��\�MsYX&c �&�+�Rb3S����ŭ�}W@�g����R�#�����	4��87��W�8�i�"�.�ꁇ���V�����-U�>XP���/)9c��x���U�:��r/�>�}ZU�v����h�Z���a`��Z��Y卺���c�W����acK��Xp����6�Ԕ����n�H��U�',>��7�nni�i7s)�ھ=pK�Ǯ�x�wdm��~v�}j@y�����cƨ���NsC�껼�D0�sڕ�V���}��b�)�[�L�])�FH2�w����2MȪ��>|W�� h)�h�?ɬ�c�
K׿	S�G�bAA�4�@Vf��.s�^��w��C=O�<t.M����9�-��fG##E�����V��V��-zn5f����MZeE���d������X�]���l�H�+�$|q+�Y�!oS5�GE�yr��x����G�kD/����M��yv{j�uu}�;�&e}R㒦���lf��=\{�g;U2����M*�.ì-�_�%#����u/N���6ܘ��!�	`=��>���?�(rm�j=g� |o�
sq��\@ѨUځ�1|7�����O�]�bN�?�Z���,�T�$a+JQ��{D�Sw�b{Np�D[be������^<�ff�}^wE�_!2�$JKH>V.<���݁�'����� ���0WP<�xo��U�9V�l !��j�VE�����	�:�~JV���a���8s��_�|�tg~f�1%�.�θ\<f��r��B�#�_�`_���*��7F�#JJ"�"?IJ�&��zIAu�Vz`����yHXϔ[�A��ʕ�=���K���hA�"�2$����mO��]V��[�y,����~1Xvp��ZJO���P�I�j�?՛���~���qh0�]�vv�=7u���j��=�T��{:UfffeT}_]�:�HV����:�d��t�>���\A��I��	�xn�6��{��>I:Ï/��i��h��!�����6�#��w!_���8ި��,E��:��'n���
��k��-�3��9%�AJ^��,--��x9�i�1DcՐJ9Y�g�6���콳p����My"����p��v����ڵ�]�R'�E�s�у�3�jχd�/�ʒ	!�㉝jz5$İ��j��E}֟�󊮲3Q�k~�]6X��1�������lyg^hE`vN	�K,S(5�&Z`��p��k�����,Ht�颣��	�%�A�n�ey�\R�����s[��d�7M$/�9���qN��r�}������T�6������5��L��R����&`$�e��GP����И�:�kH�W�v���W���\�°�ܯ��q8-<e�_�"���ú�~_�������ڠ%����S���K������N�����n �������:_1��*�t�_�O��˟a�myn7�\|��@�$ �	
���4��9�Y�������acl�z闱��BC{�):z�_��Z\����șt���W��y�ya� t����#�|���R�4�]�҇^�O��g�ӽ^��`��"�AqK�U�T�຦��M�&��jF��c�}�6�g��u�~{C�'!!�b��?��� S\Hn ���K��]AFy�O{O��13��/x�~y�- d��+��<N�e�O2!Jܕ0�s��S����8�?���W�������~<��n����9c �4�J���q����p�)}���oyi�.�;b6p<���Og�9Z�O	B���>��֓3Ǳ	�
��|{�x�.���J�	��|�>=zqUf�Di��s������y������P�����Bd��nD([��x�)��γsx�R�*����BՍuT�\�^$�O}��"J�0 ��,x*Ͱ�������m������/�MG����cy�M[��J�Q.{+�-t��/ar�[����V+��"��L�e[2��h��
cVr���TY0�D=��Q�3ߚ����M��P�{�:l\ 7u$�V�����~70��Gs�W4o=qj���y����7����f�����1b��D���XTbd�T˩��Y0�[\��tB����C/�`��)�_�'0��d1%���I� �y�|��ı�EX�,�+��H�vu�=�7�rƑ�ii��y9Q5N�s���:�v�L�n ��7����4�f��(CƧ����v��i?�#�����Iۅ[(��9^[�_<� �{p��2�v�d�{��|�)�)����1��$Q�2rEV����@�C^G˷,\��]y(��m�����,�Wb�����w��ff^C�C�Fs�2d�F�
^$�\�++�Zδ<2@]����\2��0��¨+�Pj����F#4������*�ǃT���P1M5��>��eQwF#�]�P`��w0\�̬�&Es �O�������.��*j[p����������D�l�l5���R������4�D�ܲ�Ng�t`����/����<����ꥊ��;,D��������!J>�4����}�s�r�����l�;o2�MM�JA�ƉWe>O�H����-�1]���j�k�[3�ƽOGmq�#օ�2��+����ػ��СV�d"�������$O��@���V9�0 ;B�11	�f����ZWG��LE`a)��1�(}|܇����C��o�뫬���Q�p�/X� )��n�\�(Ri��:�=����f�~-�	�[j�Se�$��{WY�����ʻ�������z�v��`e���m7ƿڵ�.vx=�1L�r��@����vK�z$c!]*\�ݸ�j���щ."�ә�%�d�EQ�c���\n�W���j7$0�'$�~r�E�N**E����?aT?{�ۖ�,=ѝ+���ji���]?'������L���~��m�e0�����:�������� ͆����}'!]%:rM@�8j?R>����m$��~��4T�`�f����촄_�Y&�jj0�r�s��)UB�'5UKk>��iT/Z��>��1G�%Zq������!7~Y*dr�v<�%�	��O�wR�6�}��t,3��H��ٵ��УNH�zc�1��~�-30��[K����D�K�Y����c�)�Ƴ��iN�t\�&��B��K:(��������M�|,�_��3MDw?WK?�r>	�l�[�|h3mtL���v7�rѱ��0J�'7�hՌ���yd��2��[�}��*>���?Cg�Fg��{	
��Xo�#"��AR<�/7W*������j��� �3�)�~j�<X����)st��}��?O��N�Q{���`pi"����@M���/���آ��r+y�� �'n88��8������{tq�Q�L��`@�q��w>vf1wµSR������i�́��^����+1 !����U�k2J�V��� ����F�
�Ry�;Y�O11��v�_p%̿��*b\�;��A2KlSIme��6�������V�"�����+6��u�ȫ�Ulum0�'ǽ"��SS�~��)�r1�U�K~qd�˺���i��P=;Zp�x'&
~u�n���&|�
����QYw��7?�bLZ�[���Z��k�U���ANU���7?uV�t�?׾�؛�\U��£�Bub0}5������{Չ17W#�$��ibl�(���h7���1+�ۈ Z������c���?0�;!��6<�uu� ���Ɛ�GH����&��B�1ܟ�S���|�i˪v�x��6����	��dn軉sS��0�N�}�ÅI�,�,���b����i�!���� =�l�g
`�|ߋ���'���N+=ۋ�%�M�0(�M8m��4+�g�!%���N����i)7��Bk�h�W�n7�����jq�����+$�1��hL�����K}� �eU�!�Rp��6i(h����_��s��
t"2(J��������C�z��Ps�߰+}�wAJ'h16v<�n��Qا+�2�b��s����_���?sD�$dO���M�ڝ1����b�R�s�ׇ�%�.³Aj���W����X���V�7���#��]ó�h1팒s���x��W�\��8���pMM�ט�@ʄ���'��F��!��=X�@W#�\*�[z�iC��{��4�I���?b:�w�/n�!eE9��{����3����E�b�H��`-�+[^��Aly���չ�Fͱ�>�YJ-���(��F%��/:�dp��>�/ ��x+C�^i	���q]I"�9�B@?,�b�{����Xl���h���B���i�;b&����Y�J(+t�!����Q��J�Lzv%����Q��F ��]���$;(BO�Ř�q���yJ���FY~ ��T��s6�â��o�i7�f@~<[���c�>fwu�5��`�
��7�$���%;32*��DCuL^Du!Q�y�C*��W����P�E$����W[@�H�G(o��~����������	L���P0��b`��tH���]NG*ͨ)�^ڌ�����jH�A��z^�xu��&�aK������#�Q���Kx(�	k���x�u���T]'�v=��Z��=�DH2�����ю!��\6�}�Y��gDM��,�5^_w儾���d*�ۡ71��[���F�+��>��2��1z�V�.�'�t�2���,YԵ��BT�ʾ���f�?;Y]�^�-6]��p�'��Ƶ*8}T�����݄ZqSdi'N� Fql�i^��::Fʑ�}��t�{w����եW-�������nNz����G׀Y�,/+�n��e4�!?�eB]���Gi��4-��e�����3�~}�!��R����MM˂Yh�δOmIr�����-'1��
'��>��9�n��$nnjcMҿ�,�1:�
E�Ʀ�g���)r�\�����ec�j��n
((*�]���ϳ����G���9��,/�����j�t�j�rt������ͬ!�؊P��6�`G�gᣓ�P��Ĵ�y�'A��G(uqޖ���V��%9�2]�=��k��bu�5A�{H�]gwp������7�!#Tw�m;]<�� #D�Y�tB`J�6y�ܟx*.frd�Re���j֑޼6�]1}��3b��C��(/��ܼ�i���>їH�|$��yfq|�'��M�.��,�_fNM���?"$6R}
��9.��@\��=?����2�Fs;Pmj�023H�tv��`�}�������=���Ѽ�#�d��
2��ݾǏ�����?�M��s�!��bFjB�\��O�J�r�񣝣	�TDLfU	 R�r;I	]��t��F����_��n43#pp���<ݛ��BÅ���s�0	�\h�����~�L�LKН�^9y���'�gw���O�6� ��P�=��!Y���
t��9 #�}��s6G-�硰(&^ݫ|��{�sQ;�??�iv��귯��jT�{�����d�ٴ� 3������*�,������)C��kdEG��2$0:Y��\Kh}�a�3���5e�u<\�}�-�#%��)�1���M���Ѩ)ٛ%��"�Aj�~�0����۾�K�ٺ FH!}�`T�����T���L�9�G��|㪛��Bc��EF���|�I�\9����Go'O/;?u�7��>�#����� �D�������"G�B\X��:UK�����DU���_G�n5 �%��SqJ9�tb_ϙ?�����j���u�yX���gCE���M�:�;ɫK҆�ӹp�`��Ų�.��zL�? `�E��~�]���}�g��L7�i���JO'V�ȟ�-�L��h$rKCS��2kԡ�=d0���A����ht�J3j�~<��}�^Q��6�РP��yy����du:��BQ�">q�c%��Sn�t3�n
�@����Ё�z�T�""G
���dyu��I�:�Zna��c�a�b��I�2R�g�Ǩb��\\�ڳ���kS+�1٣���(��.�H����b�v����>u��ϝf���7Ǥ�p�<�BG!���M<�vO��NIɰ<mi��8����}�������W>�u��#3k!��3
�MZ�΀����8���<�a�Td��r 쭿uBr�!��奬�X�m����&�z�����&j�8����A����Ŗ���ezŬZ�}J�twG)����D���ҐŲ� �u+������̼������w%��| �b�	2<s:��D e���p
��5eܘ����!Jƕ�w���͗�>�U@��o��/4A�o2n�|y���P�6����0�z�����8�EeQx�P<1��~����[�g��b����a9�$j�n�ru-��=y��=��5Zu!�	7ξ�7�i��c���!DI�2�X�K�!�][s��w9ZT�(�ى�|�N#"/�2@�a�����P�Ú�Q+��it8Q��;R�#WN��Z�'�)� �	��B^M��O�vg�nIJ�h�Ҏ��#�	�7�]��?�q˚��q�5�!::��I��%srl}�����5h��0h���"���us@�*]"J�si�n��n�oM����u`
Sj'���f�~��h�q+��i�ٹ��l<�X,G�����u=��Jz��1���p��Rɏe#r�f��6��C���I�de=�v�2��U�E�������8�>�@0�-�b4Szo����Z���M0���_�Y4���ai47/M��T�cb���{o��#��D��guL�rۉ�YBDީ E�!P!'.�O�u�^�XLy*`x{R���?:��ۼ��7���1)RP��|(J_��Д[�kux�����tEEE���c@�<>�V2�+H��r����S�����ǒ�W�>�	_v3����+s�Ю�ANŝ眸a�)p*��H.v ���1�I���En�3�
�I������Oo�b�t�u<��\rW����0��V&����pd���[�ۨ��eSa��I��mU|�N7��!D��S��D�ff�,|]:P-� �ws�CR��lT���M��p���u���}��U��ڋ���3��D�������bP09M'Q�V�`�.~͆��'ׅ���B���^�U��(�8�}�3/�n�ʿ�!_Y��:����P�<��W�^��z����7�4���p�GU����	uvu�H=�H=��zbS���$ڶ�:7�é�Ԭ���آ�_�=���1n0ra��d4��z��F�"!.h�I�Χ������6�F݉�.vZ��<-B�{��'�Į���&;0��YoX��n��){��Jt���g�H;�W��@m�<m�R=8OS[�\Z�ȵ�,��j�g�c�O)�1ZS%7�+�>Q�˂p���ӳfoH����AA�xL�<,�m���.�B^�i��1ϒs��kOy�<�!._~8-����-gv���=u=L�~{i)�q)��F�����gVK��K~w�ܷӥ�-3������7�R���E~@~��g�y��N۾���B���<b6��,"�bk�'�C3�B�AY:>�#��w�Q�و�P�B�_4��qX?c7ư�)o��U|���|	��o���V�Z2�h<�?���U�D��o�va��?y�7P��_����W�x�^���q�װ� �:�֬��u��Nb&D��|�%�]�r�oENR9;��ȏ��߹�8�������1�,���	�{�oLy��|���Eb�Ϋn��%f'Sm�*O~_%���^DYu��Xy�)XHz���Aj~�(�h�q����~����0�v����2<xx|T���,!��)1�g�w\�L�G_G��`"`��[���*��h<"l�2j��pГ"=nNBt��>���SX>ɘQ.�U��HR������ގ�l���M��n����uԄ�b�� d�z��Sox�[~p=��*�0��z g��K�����/Ưr֐�_��a��_�)B	�-|�tq���i�����W��Xd[�Gw?���6*h�z��x4�(�݉g[���=duGr*U�?V�6>6�L�ݒ�����_ۣa���	X��n����V�̊R��l�5�+.c⿜6@�����ƙ��;��yC�^�-x��VC��WI�n˹��5%�\8E�V�?K=.��埏��>���$�� �ԛ������r�o�u[q5����O?���DM~�8�۴���=Q�,�u�$�{��H�i�:�9�����Tkn+�B�D:S��ϖ�ͺ�5
z>�W�E|���^�H�VK���1VFRϛQ]�*���-C�PX�^s�����B�t���iːV���;7^�6Dbt����/����#�Z*)b(�(�!H&nn.P��w�×�x����xSS�`�%�RS���I��P��оJ;���2��c�������E�+-���P֨��0�e�1�r��̮�^q��Œ{���_^���\;o�5����4�
rΈD�^<�j�V���[`�����җ鍍|u�t(�P���C�$g��q�k�qQ�)�`���G[��[��B�M^�Pp�DFy�{�����>�0�E������z�gޯL\���2�V˪���x���NK����S EQq����$�[<[X�m��tk�a6j,G�����S���b9Y\Ћ&�:��;kW�d5�;}��#%��,M��mr���11C����7[�/X/w���G���O��]�u�GX���W��:땓%��-��;9O�yAZ��#ڠ�@���8 ���q����Q�rλ�O8��Ū�v�+�2'�&u�pQ?�2]G�4%�*���>u_h�a�k��p�Ͱng,�5Lo>��x���ShS����;�D�l%�؉g�)o"��*횳G;��_cM٦qJ��mp;�	A����}KLO�m/�����3�*79�
�jN�q�e����e���mw��	 ��ef϶����p�׬wd-��C�����Nl<�Ȥ[����� �"N��	.G�pt��%şf���)H��ĸ�"7W`Q -�C.vH����q@]�x�jd�!��� s��9Z��F�پ�Q;Q�W�Q�̋���3h�5XcY�`ڝ�MA���Dc��dl�^���*����"�A;���iFT�G����N�]Y��)�Q9,�4�����4>�y��g�on�vN\��C2sN���"��$����������J�j&Hm+7�L(I\)_t�}(Ğ�Xf��T��j�UW�o�9��S������GGY��r�ŝK�5c+G���'-�J��J^���}�J�i��Li��!K6.�����T@Hb�#�K-�)�~68(s����6B�F˼�UJ.s�V��[�Y�B�N9Yd|���<��Ȭ�#F��{���qv ����"�dGs�0���>���i	'.xo75���aA�ؠ������v{�岽I���M�%7��iT�9�}�snX�h�7(���ѵꝦ�	ӿ��{$cŔˋ���r�����I�U!�mc�
�G��A,�?zR�/_����@�#z�^e�."�n��i:LG�����A�a�����\�{+'���?��nZo��VI��9Y,B7���@EG���v@P?"��Ŵz`��J#�T@��~-WįE�H�9����F�m��Z�R�����J7^����;"r��A���.R�@	�C�1ж����mm�\X�g΁��,q���-»\��/M�
�F�����9i���$���x��ML�(<�k�dC[n^6�Y�~���t���9CT�T��:�V6҆&(mdt� ���m���!�G���4�%8�� ��̓�?�V/+6����Z	�o����w;�[;ItݖB��aPQV�-AI���� �����n5�s>�^9��.��5��@+�,�L���Ifo�b�j��ˌ���+�����OI��;Vbb�]�q����K:&S��Ϲ;0u��3��-d%}��E���� � ʶ�yq�'#)�f4���  ��θ���,�����֋�P'��Q�v���"��KpqB#e���14T����̴��#�5��*�Pv�����i��a�a� ��gb�
�\��S�o�1���� ���w���m�iv�Y$K��&-�;b�</��fВ�R�d�p���o�o�b��E�>r��4PY�L�#�g����S�z�?{X8^��B�[�Q4��TZ    �֕�7�������G9!(�(���ZP��G�a�+^����r੿6�9�O��V���n�
��K����dBU>*���s���9Y|��!�)|4�AbΒ�1���j����w1�7��r�-pO,��7�+���ȣ��[	@��'o����fB�ŕ��x�I,��� �u�nA����DS�`%P�
9���x��d��ø*s��.���V���YɃ�)�E���{�E�JY���*�||'��N��R����"�;��YG�l<�Rt��mHS9g�^�,�a��b`���=\���ѯ�tB�w�O��Khh��~L��uy���� �,ʉ�JYq��
�y��m_�~��v�]OĎ��������� h���娼�ҁ��J�6�
�(��&����`*��<ˏ���LJ�-���{8�h����i�T��M�9�F/����Ncz�k&�b� 1I����y ki,-�p������x��L�@_xT�<���>�pM#rif��m�,�lǂ�����~���:.�YϺ#�� ���]kF𣰐�**��Q�Z��vʼ���u�D����^��n�����b�y�d���M�l�Ҩ^-�w�e�(�x~���pg���Y�G�8[3_���]��`���Nօ�>L��Hgݮ�p��Ąہ-����әRͮ��T�p� 2�:��P�Q�/3���~T�߰��^E#����<��@h�dQ�ו����	|uhzx��<��r�w?K���'O�Δ;w���~��!G�����uU0���?m,���(,?Q[
dܷ���qӖ nTt�<?�$о?V���(��P]9{}ܬ������נ���N�.�\Ov���Ǿs3\��ڸ�~ �iA�1�G����X�I��&��A�m�ϡ��-��Lq%�i�+��3e=NFI�*V�Y�7�O<9"�ac���1�L�)w�M^&�.eX �Дկ����j�����DD�SO`D5������%`��Q�j�I?����`�$��`�� �n�wet�����(��K[7<���n_11��!�%}��b3�PGqӏM�[h?�ɐU�[����b�15^\�u0J�U�V�����}�yA���	�K
Uj�>W�;K� U�܆�-�'�x%@׉HOײ�U�8��jm�8�[gLdt�h9='!���]!�P��]U6��H��j�f+�JLǛV���U��8�:�1�M�4%t��%t-<�;m�t��h*�|��=(�K�'���i*Aǌ�8�EF�;��� �8܀%�&�Wr�L~~�V!��R�B%2Q/r��dnC�k@�U�RwWב�󍍘`�sT����Q�o��,�����\��w�,&Q��Ѷ��Ƹ��&6B91����P���<t�y^���uT'����0���4��p��i���`Z̔9 \V��9Pԯ���6޴T�<ݖ'l��$��d��2��RS.��E�1��)B�7�#캊�7/`]~ ;A�Y� v	��Dpo�����*Ɔ�8g�����M��n?r?��,A}!MTaM�h�MEN5E�*��<���hV���.���婤�蓒
��?�+��1m���N���h|*W�Vjl��ԝ��;�@�/$D�F��%��=��)�I[PR��!!��66�>��;�MB����o�Pw�4>^�ML�ء`E�����v��ˑ���x�n��Z��8��혤Z����m7�=_��p�׻��{��iۣS&��%0����Z��c��){�-:��D�@�a��^��	]!���3-�6!xO#��7�.8O�Wn�eVH��j+	A%e�~� �b;Y�J�
��a!
�GǕR�������#L�y��q�`���N�~�')�� <+����_7sd��Ɍ8��� ����Ӧ%� �復�zV`qf?n�M9&H��j\H�B��MUC�5bl���eծSS�v�UӃ�^�-��nωUx��k�N���^6�UT�T���u�
h��x��ǃ��.�>$�yV� �0�_�ʷ��̧}�4O���D9Q�va�>Ww>:Pр6���O�n#�hq�Q�>�׊��jV�@آQ�Ɂ6ѫ��b�����'(rNǯ����]:AP�Ol�ٚ��h��!Ѫ��:L�P.S�I:�O-Nt��-a#5��!��M@�N;#-��=��P�O���#�ӌ
_�ĸ���#�O�n�X���;GXnj55��8����~��U���^?w����B��w��	�л�� ����Q�Z�'n{ykG"�f�k��Ō]�R����vp<̂�=��=ᆛX��/�X~�L7Y�}e�c��ƈ"��
v�5K��ը*�q:ݒ_H5/�h�(�98,�����
`�ffIHjoy"E��<=O��s{�R��H���vff.\�����ꏖ��_�^���a���0\Z�R�7�"p��Ӄ��y��-���I&T���<}@Vs����n�[��c�C@�h���Dv�=q?[q@���PVn�p�,�V=�'x����x�۠������9���V�����9�'�Ϲ���Cm�ﾜ0gq !���[��kk?D��(@�·V�D���������_r;���%�"	�I�D�ftT푪��kh���5V���-�vz��R[ʏf�29 ���G�P-�=�'g�&������2�Dk�O62V�$o��3d��O���4�߮�h5��U��dz�;Ob��g�
0�F&�Gp�	�r��Be��"���m�
�67'���':�-��;�?�D;������5XOԶ=��Y�F�^�tE���������À����h����7�٠Ɏ���Ɇz����2�(m17����C�n���[.w&1�k�f�Mh�.X�f���1ݿ��eh�Ȇ1�jn{o�e_�Pff�����6*BK'y=�97�%pO��HV?�m���A�����S�bo��{��Y=���aݝ�"V�������E�EdJJ���JS'w�_{\�?�S��K�c@�YO�RG����N�"���2�+��%���������nO��*��0�Q8n#ë����}d����@��N�TI���߀՛�&]�d#�@�9:E\�J<�k��P�r���SV)l?�t�J�����i�`#��^g窜�d���s,1gϸ�����wn��(�Q	֑-�tq��B���`ny;	�����G�kif#�A�������|�v��Y<qόi��hW�d�����n9�����T�ҥ�����c?Rz�VJ��C��:�Z:*�8�>p�h������������:Z����Y�9/y�qt}N��#)\�I���sA��+C���M�/��1�8��ݜ:����8� ���KCh{��.	��mN�ڿ�ԓȫ�r �JK:R�g�&�E�J����jg��	����n��|<;�V�M�j��ng���@_H�huc�)�Ӷ�\���OZJL-{g'$ViS�u��s��[���(qH�~��a/�BQ�$a�m�2���?�T��4��~j�B*�N�w�� ��|��OB44�TW�W���FrwӀ�z�`��=�G���vT��{�m��X�Y�v ��������E���0��1�`\����ЕA�ٿ���Y�sw���ym���I;x�c9�&�(���z8�g�_��=�2��o�
mJ���P��/c�o�gM���?��������[j��ں�J�S��i�aRTp��$��(�d�U}�ͱ�i�M�٪$H� :M/��9YO��MOM!EV+��>W4э�늛:;)�.����^�����#��z�2�����i��}�����F՞f�2�6<|�I�FJ�E0D�]q]����o��Y/ʁ�EU�6�"GZ�F:�C�e���_����ڭ���2�+b0/��t@���E��'JF~�����(�>��5���a�Ձ����ۀ��r�!C�w�����Do>���B�Ѿ�v�T�S�]荷K���$��D{B��x��UGG�rSu=ozb��������3?��*�9qvؗ�Ϭ�� �`h-o����Y@����d�
w5�B#�;���PPgS�ө7��?�r�r{d�[��,��Yq�����9k�C_�#8�3
�裣���Y8\u�p�9B\��{���}SS�B��(S+��ՄAդ�Rn^�\^Q!`�����y�%`o��Ȁ��H��<_��z�j�!����R�� ��8EޫJK�}���{��v{�_������H�F-����l���5,`nn�d�G�/iU�_YS��f�n|	�G��rҿ�^T�'�z��4��U��L-rh/���R��ɉۣ5�5�9!@2�w9 �c�e�Σ[�b&ȹ����˝��3�s/��#��?f��������r���j��y�HL귒E�[0����e���K����e,T{F��H����Clz:�Y:�'}A�L��\���ѷ�>t�P'�������xyaGiE0=��97 �z>R��{�V����1v[��CDŅY�j�$��Y��q�`���2྘����	�k��@G�ch�ur��0a=P���%�a���o��<�r���60�uKb""��g2"������|ǃ���\�DK��N���7�@IU�1��A�r�w��E}Q����C�:�_��n{�v`��kJµv:O[3wmD1���u��F���s��d��g�?��t�]���$i�z��*0 A�<f��_u�Iw��+M*���3��*�KF}�ſK;�Gr:���h:'A祬�lH?/;�.W�.����c�nC��C����K#&�e�`e�2x�᭭$�����^����G� ��j�9�}D�,�M����P�"���"9@�T�O�Z�r2g	�����BET��ɮ����9�A����
��R֨��rҧ���-��o�im}IB�ݷa����S�d|N�U�d��F}�J���
��g��qڬ&��3= u� ���d�0Q[+��W!��2Ն����F����0eӂOrkf�ڱM����7*���xLi?$d�g8+���,��+���-��Q6�ͺ-�����I�ˏ݄ޗ��v�V�	.o������ݐ"`,Ks�$���Vƍc�` �́�c6Z��TbteU����5�޴��c���N�m۫<xv�qa	q�g�1܅���������2�uع0t�d��{9d��FI�p���t��0��u}7j�nS�<�M��������7�R�T���b7��ka�ग��ww�rV^Q�`�:�N�Œ܏�Ry��n:�y�+����FDཱྀ����x��R;��b�۵��e���ߢD%գ�;~~���0c��5,�f>�����I��p�����̇�`u:TN�BB�����P*͌���5��������mZ�8��V�d8�aC_s��`z�������eIvܰ���R�qF�Js���j�VHJ�+��jಉ{�5.΅��g�/T�0��H9��.����;��<�����04+"�T�l�+H���t��1�(E��t� M�
H����A��������K�<1yvޙ{��;3��)�C�%��<E�e#'�8���8aR�%��p�&��rF+:n ��u2�תk��z�<Y8G�zEEm׉�;1��(�9)��i���X����G���=E"�\��]�UK�'�l��.޴�7(��9�88XCB"��k�s�K��Y�i���<*Y.m��C�� �x"y0}���Z����Pob�{K��{J
���p���#t9�@b5g�Ͳ��7$��%��r�~���<�II1,�8 "F�#��ĭ�<O�hm�w����\Ά2쭞��sl	���A /�.����S-Ʊ�yĚp��o���x�F��FZ>�e#�(�N���D��@A�2^��%6�oLbk��W15�]@76��)�����ߛ`�}�8I�{waJEzv�KM\X��y8�PSC�|�����������"��{�ap�M!Rh{}��cK�*zyܯ`��`�6l�=��h����V���O��4T�KW��S[Uz�}0���Z�Ͷ��F��\����g���Ȉ��9O�S�V;���BMήG�Y͗
�b\�����B�l��)���.e���	�d�~0���W�+����?�c�]��f�>4�u".��l��/����D��Esө�c��BY{|�n� ~I���V��N�nQY��6M&&�����C�~��8��i��Z���Ы36�t7�tnY@5����m
<���F_4�w\�捖t zN� ԕ%���{x�ۦF������Fb�M�� �<�=�%v�KRH�v����$K0��P����|5: ����	�"Jn�}�ίB�Vo�%�D�FF4�͓&;��c��b�a���v�${�$�X�g��E$���� �Vz�������_�NQ�����ݜ�W&����eNY���Ձ��ӺD�C��($c(A���e���3*��Rw��W��;!��b��2-ҷa�4{�xX%�$����Z�Dj�f~����V���䎼�~��|�R�����+x꠼�J���%��CM��~|۲�5O���๞�����ɹ�8�7�w�V�6�9ρP��уM���cK*@b�\�޶i�FX���������e!h��G��g �а���΋�~����\�t�wYF?2]�n �Cw�� ������Nܡ�BAT��è��1i��k?��B�4�`[��W�S�VX��ş?�DϽ2޽��w�����%��|,2j���w�7A�4���S�.���i0q@�忴��ʋ3����n�������U~�y��rR�?�u�<��tK86�\́�� �ŠF�qG�/�q���Iڻ�Ѫ������b�pY
�i���,MH�����X�Ngv�::8�Ļ>�h#Z�c(`Svt�ԥ��͗rv �Y9����1�-:6�+�Ӝ�֢�Uz?����0ޟ��Y2�K/�;.�=&�.JJ�Q+�#���r��hW�:*\ĉP���nu|R��=��=�cc���o�'�J�?w!{o��H�YG`U���R����镏?�����;̨���g���z�6B�6t�3$��A��H���zA3 �9O�C�.��ď�њ����ƭ�p���}�^�w�ѣ��	7���~�Ue��BM�:�7q�8�M_P�C�(���z��_1�� �˾�����'G'wCf3ʤ�F:Kڒ�E�![�����әz����W��Jf�أl4ZAbS�4m��)�[����/~{m�,t1԰��DD,��� U��7lGߊI�Ӳ��~�	$�ݸ�b����B�L�q���É�)�$W<}�i�����	�������"�b�g,��Jk˝�A�"�BBaP���q��~�x�4ָl�������Uh��SK�N+�<�m�r�P:,���J��ԫ������O�o��DD�c��Z�g)ҍ�I��޾�I��g�n�l��r{zvFYY#D4��l�ф�k�%cÊ�S�XB���%�n��DKn/�I_9
�+Nc�i��79�v}�bB�ϲ�l��m��`x;hy����T(��~�$�c1��Wc���S<W7;&�s΁Mk�Ub�L}7NL0�	��(}\nQЅ=�LK�$ߌ����c���,�\Jܖꇬҿ/�EF}�q9���i[93[�~�mj:�{PԱ�d'7v�
O��1}�TDa���HQ��F3xz�kwg�����&�R5y���$%Y��D��(����R���y�E���뫿�.�hu���Yƈh���c4����Z�����߅�� Q�,�8�hП��� ,r�5~{�:!�-�����}�+��K﷋����GY��E�{�,�P�r�Z�µv�ŋ��ب�^|k�����!���{B�r�7~��a6 �}u��Wbj���2'��vᑟ���i#����ST�X�"b���~Sîo�tC��X�������jf}�lM��a�E_p4Ɇ���y��Ҵ?�N(Ei��U��B_Q�Oo��5�.0?��W236P9�C>�x���.�_�ca�Eu�67�i����Q�xz슼:�|�v�7�_��
�Ѷ�[�|��xVԞ;��^H�w���C���Ӿ6e1[m�0�g�s�P���M��4�1���`���ˁ{��l�ҋ	� �� vP^��	��aߠA��K��}���8�8�Gܹ$�^rcB��2�N�� f�u���%h>���EW�a�i׋4p����Y�G��^�Ǯf-�T��������}y=�,�*eVQҟ`ө���q�$���q�w����@�����Bm�
�l]����d�%n����s�COA�����8Q����x�=<�u�����\'��.�	�JI���z�$�t4�5Q�_p��!�=K�|���W=v�K�±� ��cg!�]�~��AA�����B���6�y�V���w8(�Z(��V6�额v��ފϵK���K�Y�|�1Rػ��ߎP��r��&��P��<����갈E��[�t�wD����I�;�jF���yc/Q��`+K+2�h��\
��.���r�:�`��Zb�X���ŚTib��xgB
`�v[VA+t����]������@��$*��ǆ� ��#��.��.��準}�M�!hEޒL�3"q[�v���e�G?�D��on4A��V2�(�qlY�c�(��H�L�,��]\�֬���i��¤z������4ɫ5T�&��wYD���:�z��O�W�l��>�P���W���w�S�I�NPV�����p�)tDu%+��!�}�F���l����9����:�C_�p���Z����z.��n�J+c��ӈ����K���y�h��
�'6�}g����@f��������=9�K�Iv'�$L��e������]�s��SB�y��v�E\�7�B��wJ�}b���E$�4"i鸳�O�r�������Ob�:P�����B��v:��K�	��@��7�=>�m(�&�a���6@E�r�E�c`��U��������E�ӯ��h�B�ÍEZIc��RwG�s�S�En���$]�tjrD�n��Ŷ����=cά U_tɌ���&@�b88  q���Y�F08���1�[ �x|����x�;�-qb���'���us�Sn����q܉u�n�!dkϰq�~��e@�hlh���Ǣ_�l�!:�㝇�����K�8%o�x
@�����}~nl�!��L���'
���5x�����|a{SY��2��gP���x	vdа�	w��#�IJ������ P�`	�-ЗM�|�����	�|�އ�a�e���u����c/V�b�ޙ)v=X����s�oEm�6���H��]���aUA�	��l@V�h��o�$�l�/���^_�����b�+�;��aE�oT�B��zI�<7N��йW���.��Ad��V�i���ǋ�	2mHY3��g�+Z������
�3�,�;��I�d��N�L�b��j{��
�y�ڤ�^w""6b�������;=�e짤Y����*gAڙ/���9��J�d�
�ׇ��7{b�ݺ��,m�1�Qo�8��3$��g}5?�H���WRc�G�ñ�i�{�(�-�[��������o�h�q�����[F)��H�[����|�p�������E]�^f8���+t���M���,9�H�[�0���twgĝH��-F�j{"�w��B������1��� '��I�c��(��;eq\��zn슈�d߾�~�;߃?�z�J�=I�'�I�[u����F�XП�9��\Bͩ���g�T�ywR:���\t�K|}����j�7���[i_�/ǿ9_^��~��(U�߳�,ӉKK�Gq0���b]�~�u����:��k�]9#��P��Y�������W��}T��y�:)K�rDq����܊�I�pɩ)C��/�6�N��a����5��m���}�����(K��ݑ1H�1�����1���(Ov��f�!{��N'zZZ�o�^��l��N~�f�:�%�V���B��VL�J.瞇Ǜ��vvq�g*��abd�	"�����������/0)c�����Nn� �8��muu���J��׆�U��h}��W~׍�.;�z)���\����\�f^��4�;{C����;�X�C��xx��g���k�՚[+��{�k�n�̺!V6�T`��n�f����;�\��.��Ǝ9��^֙�n�*��h���k�:��Yп`=g�Mu?��I2�d9,'�z���/���3H�����#�Ǚ��E%( 
�ru�s�%6v4OsZ�/g���۳5��s+���[�Lj�}�kS,��dh?���&Ox��;�I�����ۛ����[[z����AR&t�_ъ7ܰ�H����/�t��%f��l����Y �/`E��9�}�DO����
�s�4�W��g"+���;�j��>p��
6���ٕ()��~��m��{E̋��y˓����V=�է�O HF>t��k7VBkC����|��lt$: �����⢞5=�^o��3��s�Sw����hh�Q��`D�~����C%R�O�I��SzI����/�wϊ�UQ=�?��c'+�$1�U]=����,��ie��L�E�E6g�To���4�ܲN+��%g���f�x���jT��-!��ِ�	a��C@b�m]~��4d���؝���[�f�㑕�X����>���a�m�S�Z�f惆��U�"8/8��s�	m�<���j�}���W/��m*z�.���{t��H�-A%;vT>��JxR2��;`�귳	ņ�ev�~�	�q~_���oB����Q�3�x��c���'���*]���#��s��I=��e��\�H��z�t�D�{`��qq5!���ƛ��[[�7���}1�ЦT_qZ�d�![ ���!:�F:�M=
�r�D���ya��{����b>p֤dۑl��#�
�K.����=f��*˗"l��j��LG�:Q(�V4��^i�S��s���j�
 <��rH|�r�y�
S��9�)G7��[I�81.���\�r���'��tXa�23��c���dLA��s ��@����_������X��P��CF������b�B��)�az�J"���ޮ]#�{�����)�Jzazz�;ү���1����e6zU���b����i�&��ГD ��I���,	�.$�=�-���tR��q��{=qU,H?|�1buu��S#�T�;����R1L���g���]�Nv �Z��]���;3P�.]:�>1��nn��Y�Ei�fxlF�������glc���:2`����hii9mp����?.FŒ�O�f�LHg�L���Q��<�J@��T�\���V�(��q��������8�
Б'n-��e�@��<�ttTQ<�~un�� ��\��f�O��.;�0 �^��YR��[/����BE��@>(�����!?�ʙ�X���`2p���LN]��-��R��d{JiΥ%�j�T�eS��[Kg��<�cI����gYE�ͱ�Gy	J�(���c�r������g�q�P6X�)�֎���W�e�o��2���'���
�h!�t{ʷ[�����ji)�|��D_p��2RZQ�ޖ����K�����1��s�Ʊ�_<Y0^;�B��rF�Ui<�.h9ʶvׁ�O �z[��H�ue�������@!Ʊ
��������t�����LT���U(,�b�l�uZ� Ӳ��'��S��D���e�Y�by=T�ʆ}M��7L�P���^�D�d7y�CK�7�-tL�s������*�p'������;�&�=�_p���%&g�z�]��HG�Ի�"��O=����E7<�쌉 R8�<�xWZ�;�S1��Y6;o�L/���^���+�4<�|O��ʟ����-��N� �(9ߖp�0S��vH����5�z�`e&������_j��E]��s�<���/�Ѽ���o�<9!I;���k�n�$��	~��J�5�os����'��Yz����O(p����J)�BN��+����iy��4�O��x��OcO�r�lU��'��3)��f��q,O+_z��������Df�{��ŋ���s����\�k����]&gr� ���u�8\y�I��۝�/�
���lw-31��c^���Y�l�kg��L�D5p}@*����'�C�>*�;��;���n���x$z�d�\��ރ�F����迟�p!�w���n3��N�jN�-��q;��--�X������
O@5�O�;�-�T����_�� '��?�ݳ�Z/Dd󪫫���������uV�Aa�S����[��k8�x�F_����B�}���
w��P$�ܾO�La�����KYpt_!v��`J�2V}���S`�Ì9�|�n�dkk����:wGf�ckѫr������r�>��+De�r���yr���ι���oPmz��g��Rl?������(F&8�Rן<y���]�L�P�?����)��%<�n|{>����.V#�u)3��������wc���*���0[w��H\��r�v�7�P⎟�u�x龳�qϣ��3���ll�f�F����������P3���n<<�{�>��j�৷�{��F���\q�o[�ך���0�xD�s_F���dV[�py��p�YeIx~��}L.{�c�+@�
��{�(-�]�������_�گ����U!8�=H�6�,*}��G�¤�5��72u�0��E@QY���%��d����C��Y�ɟ�VL��G����u
d�l�ɂz��FNm<���o�wv�Cf}��Q+��`J�L��I���c��
�����Uo�d/�=�i�4�?��m�;�	��$�ہ� J|�}�����5=�&Q��{�>$ܿ�K�����aݢ�~zN��rp؜i����hw��`��W	uz��&�dJ�^�	����9y0w}�,�ujj[��B�� `�U�@Co�����R?}�յޥ!lV��ى�����N@�̎+����f�N�T�k�k ��ԇ��1��^�R���
�z+�ى��Y��~Tbr�n�e�&x[`��j��!ڌ!+:2:Ҳ�>:َ�l6 �)��th^^���/�%�ZVɡ2P��[{��܌��q����FƝ�(B}�˪ߚ�D�����K6N�m�S�,m)<�Kφ޴�c��G�jl�P`����� Ս�zH�'�����\���:��%!7�^�A��5){	G�ͮ:g54�DI�F�i��䮍�,�s����5\�����>4] ��5^%S��̂9�k�\�/�~~��R\PbmTI4FA'm�`-t��3���˛��V�_��Y�_v��*��d?On��b
p�����f�ڙ,�yъߏ��u΋�0~ZIួ�_��"�W��ɧ�Ɇ��%�����p�&��p)�N�k�\T� ��L�Y�O�h�k�0����`����:��:����$���jݳ1�N�X��~���Ώ��q���S���hu��)�)j�hE(�XF\xc�g��d����I���TUB�o^�d֎��γ���&�4��tB�����q��=�4�D���q��;&�AfL���]a�&���׌�ǥ�����c�y��b��/������'�>Ѥ��kA��T.��a��m���mk�D��޲�#7���6d"�=Y�����I��|H��)�U?��\]���@T~�诞�2l��	>	�7Hє7�>��<
��R2�ܵ{�>���#4��~�`<��eq��+ O�U�����z.�����K�f^5�8�#���0U��}�Hř�h����l����X�M�9)�Qm��;�B@X�2�� �(���ut��O�n�X�SVey�I��x�X����'+�޸�1�%��'ՏBtXW\4��B��Y��B�ж��n߿
4m���1<`����{�0�l���:�Rl������=�b-�;[���� 16��Â�.��=���'�25--l����D:z��~ �t�+{�*�R"I�3t�L ���yo�n�"WA��Lrb��Mw%ŵqS�Yk"J8T	�����TH�uqTYzل4|�V��R�ʷ���N��������;�I۳�j ���<�P��Oؤ�6�	4ɏ �`�E2w�9�M�09&�5$�f� �/�x���AcU0=�KֿD7��Y$�T�,��31fZ�z�����G��T��Y�2����ۇ�y.֘;�/%��+���V?������z��cGPt�vɪ�f���E��^Jn�%���(��0��'�R�}#�x���4��+.�Z�i*N�7����̰�� }Ķ~@�t$j8�uu��s��ot��b����j(tP�
�����v���Y(CM%������l�A<���3���I*0����Ke��~|�Ě6;eXFHX�%=��:��0^��u��|�77���:�;�w2y����R~�}�=�J����/��9�Ǆ�&�:�����熁 U�m:3-99z<�z���,��I�}�3�d��Ϳ�l�D�_Α
��>�I��{|V'=�1�cEsI!�����SLv�=�Ӝ[<<ڎvksKdU�:8x�Ib� �t#I.���v���,���F����\�q#'?l�t�F���e�܋Jl��ȑ�`��JG#4�̴�w�����չ(�F��o�d�bɊ�2�PUˏ՞5K�а�N�� ���h�}����;�d�����
c����G*D����C�ڂ�ΚD����.J��:�(�7If��ZeЈ񽖞�`�G���z���݀$/T���k5Y�h�]S.�k��׺S�A��2��BS�����&Zd{|�@mf�p�t�c�7��Β�Za�2Y]|�kG���#��[�����k�Z�BY��G�=�Y�B$����?��rK~�@�g���]�9!:?���><y"I{��{��o*��l(������9����Z��[U5��m��v����)l5��������#�D[�/{guly����T�r�!Ŕ8Ɂedu$d�֥=Uq]���;���'�����(�c �?�
*��Ř��,����`c0���g�h{����6�J7�ZX�,�Y����Z�`j����/�O�J�B	ސn��NlO�����_�G~9vz�TQi޲1�9?���J��:J�c ��Z��Zk��@����=���;8Buz�s���yk�u�=�5�����2���S�5����ǩ�3;ĸ}�>t�b�J�Q�F���.F̊ X���°� (n����{*�M:�5��G=�������}� ��9����(iQ D��"�-;mu�Cgo�RhV�ߓ�(�9�ü�D?���vNn�̱$*)��k��y�n����ٓC���I����_uP��� |c��W���f1�/�~�@�Oy�W=�tg�J�5���)��Ϻ�=9��J�0�-���	��&ܤ!
�7?'�
^������O�.���X����R��1�ɝ�Ԙ�r�p\_��Dׁ�]ļz����}�S4N ��C��3�T����iL<��Kɟ�53��+G�����}��3�A�����n�2~͍_��ؒ�	��ۓU>e�������t2 ��Ƶ-�9YGM�VV�\e��
I�~e�>�2�g��������tKg�f�R��=��w9������^'��_ʌc&�����pL����<p�A򏧕2hF᡾ӳ?hg�=�����P��F�������|�:��<)JT��QT:�Qgu���ֈd�հ'�O����9N am� ;]�����y]��l��&i�t��px�t���a����
5E����OW��q9�H
<�k��5+h��>�{4�o/��Q�2rR���H-��2��!�;S�
~��f��d�7���ﲲ�j�n�g�
�~�V��+@k�A�駲uX<��gB���c��y�¸ǻ�y��C˴����Đ<0w.��Z8E[o{����[eC����	�<FX��"��3�?��H���_t��/����5 ��ޢ_[V��7N9m��z��Q@� ˬ����� ]�M�����vT���{�RmD�ZZ���hG�9�b0nyp��&I���x-�$�R��{��;��?����7@M�{ɟ�#�i��"g�2Z���5�f��\�d�\��1�pNR���7��'�s)�$�<�5}���ĸ6M��:Ĳ���Ѭ?K��>�$�o�IZ�\��E.B�jw�~�2�w�A�s^��z>T�8�s�.4�RH�S)�f�s��1Vso�`��]�����Zo��[ u����"�b�Ny�M��xΜt(�����P.���
/���T�&,��T�&&Q�O��(�};��fW���NR8�*��~�U��T5�h�p�$Q:۞&�3��c�݊�\A�<#�\��ҋ�}Sܯu5y�m�~�O���I���X�������m��]fΤRCw\[�I��br޵�z�Rr�����L^�*��׍@���iF���^��A����;��r��E�XO	����)S�+��D�,�����f��=R��A�`Y�u��ʊ�cIa���Y>����V.�XTt�Uu4�@m���)�Άh�*���$���t�a��[ź���I7b�|��am745�\!��0�!1*�f؇M� M�1Ԅ(�e.��"p������̢$�n��t�.)��Ϲ������OZ����� 9����SU--m�,��6�j�2�'�������E6{�<bWR��$TB����3c�!���mf�|^-ࣤ�{�yN�8���P��ռ\��ڛl�4�Ɲ�P��c��#�r����#��t�/�u�X5u�8���_0�9��x�tB�)���$��<My�tzbׁm��z��1\��o��y=�/�7͠Hr�������mr�2��c^x��˄.����ܪ[r�:�jYd��
�=�Kj/\��4�|���/5h��Y#���$�� �aZ	"�S�f����a�kT�����ȣ�W�ːj����&��� �נ�4�v�u�_�O
�q�7^ⱆ
�����ퟝ�j�մo�BCE]qmZb����_��0���t���R��-�n��P��Xz�VE�_3{�Bﰊ���/+�kn���-K;
|D_��X?V����6w]��2d+I�t��9��YG�t0y�U1)�W�Z�LcW�l�+�a*d&=�����$�%�������Ը�C�~�T-�+� j-]�L�e���G�/�9e�~��B{���1��3��,��?U���"��@Uq��>ˉ�����V!��~�#x�\��(bk�Y��W;R�xdU7��7�w�7�����CЈ�a���o�1)�܄̺�h֑4�Ƿ�"��)�v����2U�� q��^�~�Z���8tih��
{g��0�����яJ~�&R�3�&��Y�PZ]�/[+x��i��&i
�U�Z��:N�X2��.^����5���,�T7T����&�Oׂ�´lf:�I�f���N%�8�b�@�}�\ŗ3�]�ת������Y\Uf�1�b�k�A2IU����u��K��@�n�Hڱ��)Y㏎�M_��B��"����z�Y;���;�9J$#��%����7�W���V>5=a�@��뮉I��Q�ba?���[����z�x=��{��
p�R�X�p<�=-`W���+�f��k%�ը��8����`& 7�K|6/�a�u��u&���{h�Q�A�C��O)rV�9{���g�5	�]�B����<������z��I�Kܕg ����|�O4~U���Q��9�����*%5U����Q��JD�}�M�ζ~�E�0YB�2�0�Y�"����U3�_��0wD��.���H<��C�7n����r޼�����]����[���b#;��8~ Ϗ���G	ʧ���x^��l�Y�t
P��vZ0R�I��u0P�3�q�I��+P��Е鳓��;e4�R�|��7�)y�n��)Bmi+�b�p�����M��+��b�hS��(E?�W�@�2H�3�f��69d�x��T�m)quw��=rcW(8f��=	��saw�9��!v�ӕ�>���U#!�p��t��t�\�;�H�A���?� �Oյ�~с������ /:V ���!��	�� �M�� ��/:�K����er�	q�o��<��k����ʕ�m�1-�M�;�0��X��)����c�S�$��NO��c�V����,�8^���;TYc`���?I�l%)QJ86J�id��킧��%�'	/	��ǭ�t�˟9�L�p�F�B_�G��lx\��\�ЬC#��$���m'��vr��g�2�؏Lk�i8�a�3D�;;J���AH���p}�d���ܢ!tx����!F�Sv�/�q	I���8B�Q��K�����1��ܾ3����79HИ�[׿(�IQ�a_Ӡ�(��*��B3e��_	gg$a�@ө��4ŕa76nȏ-֙A(\_�2Fǂ�W��?><�ڎ%|-H���4e`�)���������E(��zw�ʿ �ϣ������t:�X~O�zl����|��K�	y� ��ǎj���}�f�Ȫ��9����Wt��xx�z�>�����>	�c�Й��P�4ZH�D��$S�Ӕ�v�L�+��T� �l�; CHe�26f������jH�(�=X�b��~i	I�A5�g}^*��~��i2�De+���Z�:#�g�Z�v| ��w�*���mm�>��]U��
F�D��ȩFG�c�r.���L�v�H�Y��Ҵ�n�$A˅qy"o�5o$k���K�B�m��<}l7��+.����O1�Y����\W���d�ڕH9N?m����]Ԣ��o��� � 6���E�¢��S����9$��=+Fɟ�G����;?���ݱ�OZ@�ˤ��5E�����B����]+v�r��;s���=�37��!\zj�q�!V��Z���� QAxw�{�fv��k�<h�C*hXh_����~��ס'�w�J��ì�Wd[�?�� 1=(�7�g[dϢ�6�p�j�|���ܵM�#��抭�f��e��JKt�,�j������ ㎉�R������PݐFu<(	%����҉��!!���`^��^+_b��/ժ!c���Q8�٭�Ns��P`����X����?��HR�+~��(�����s���ruU�`F�q���of�D訰�hJ�i��'iә� vzVA�돾�e�ȡ[i��n.Ls�GZ�_�u.�eQ�}H�Y������#����~�bͦ{B�!$v���u���<���m��kSe����{hv{����M6'4&F
��_�]�bg.}(AR�����2V�g�Ũ��ۨ���T����4yQ�=��yE~&�[OOl���'._����'輒U���G�k�bI�	����ֿ]�7�Q�F�D��8_�+~hS��>j�n__�_B�x*���X��{��|��
W�G+բ1��䕭$pQ>=,漨m
0���6_e%cbsP�t�ix��	���Z�c.dޢVk�p�t;�����(�#*��Bw�f��+I��8� "-���L?J�O%n1;���O.e�㭓E�}kr3�	Ð养Z�E�]۵�E��!��u�Yl���*/pvd�|�����Uҡà���*S<�Be�Xۓ�@�+�zz\��?�6W�(NB������|�f~Dgd�6��9�-�Ф֬���2�b�;��tĹEl��O,���NI�8ZLH@��w��f�H�4��j(f	(pY,����
��e��b�U���>5��?
�a���o�jYK8:ݕa?�l����l;q���z��G<
8�<�JH����,��!�z��&��nvV/rX��r�i�(�.n��N��RT�^N^J7Q� q�����X����y�c��v�,�T�^rN�F3�J��j!��9(��Kk�k����,,(�G����׫��	��.Z��D���(pPp�(yܛ����h��:5v�;%����\�[J�Y�z��͞��F��>���K�e�+b[z�U��L�������[ぞ[+�78�	Xg
%��p޷i8O��UX'���_
$�+����ιbpS�e@�-v�y�Hq�>���tK/ը�-M�Rl)_��w�D��G���3���� �*DC�dX�i�5�}
�ߑ��ӻv���@�������d"I���x��p,-e+�}�%7�%��t���@�M��3B:����/�2��&[�M�����ݥ�k��H��<��b`��?�3����4ڝ�S�6��/���[�w�2Sr��������i�������oƋ���l����~�M�S�Qɗ�.��$���n�*����M �c��ڳj�2��R*�)3�~�+������yQ�_�з���H`�	���C���_pS�znSƘ����ף Ni��~ee�)>��5�����Lp7~�\S݅ϑ��	�c==2�(4�  ��e!q�UK]����BX��C���#�2q�τ6�1��ץ�y������eFr'��eĔQ.#�d�LtR:�!�t��jj���֯�F�ʻ�����&T�v�K�-A��C�Ƽ@]��V�-u����`3�c�އ}W�J���C|�3e`2��Tw��T�O�����-�>��,򔌝Q�IT���.�[�Y�^�4�=��@$��ɼsk�EV%LɎ�4f4E#�/"�;�왻��T��,���L���>h�H��";�"ՓX�-B�d5��Bůl{�SR���^��h�� |\�?�u�Dȶ�L<Լ��
�%6#�h��he�*��0�VA�DMK�Rh��?1�I~�c�d��a+� ����3�C���m���5]ro�ی����F6�ہ�7��J*7��մ�A�y+��Kd�;�UV��:[���Cv����[-���l��6Y���q@kq�;.�ٿm~�C��V2�TL{&�(�5�i_�CH�Q�`�znx����o}}���'�� ����R������q���Ld������:��r�Q0��L�(�á�#Z�T8�Ax��Z�fߴ���
�d��]��� ����~.>]A����-��7əx�?��8^K�C�	�^d?����ٓ�1Ɵ�>On��2]Wa�t7�v��XC7�%����m�p�Y������K
��B+[S�Xhp^T��v==j	,G5��K���Ȼ�7���)K��� <����;i��R�f��׃`�׵����BipK5���J��"�UW�xee�
�K��L��J�m��'7^C.��V6�������rAzo՗���3W�[����kP�p�-� �/ϧ���|�uE�!M\7���x��8��y?C�G�����7�"W�֢(R�@[�����s�Tt��O�3�o-�v�.����?���c��W��ixz	�j������ŖD�0�V��n���R���<��G��O+�8�>��?J�F�a}ZV���b3Y�g�e�uA��������.��@��X�_0x�������8�tZu���L`;o�f[���_�Z������7�s��lf�m�s
��u�ض�"�"�DF؊���z�kK������dy��0E��(������3NE���F-\�����!��@�K�u�C�k5�%cL8I�w��W[��:}��֕�]�>_�����&��o5S�j��\ƞ��}���*L�X�,���&����W�FFg/�≛��+ywH�v��)����syĖ}����x(�1`��c���m&
�E��5�<�6xgL�����8�'�2�7��kC�C��:�R�u�_C0�{$=��Y�3��T�`�9P��ĀGd���h�'�a�D(3J�.g���q�^rn�}l:��Аʽ[���%Z�#%*�!�~Ҋd_��b�?xT�y�-|���N��J����+e����f�c�#�(�tP>:�_+u�~U� �ԫJ+z7���<r�:�1��v<���1m�.x���'�	z�{@�������)q�ʘq�B<��M��J�H1��O9�"�i�=���^�L`��9��������_�	F�>'?����L�W�KЯR��T�w�ק3�KL����=��ոI���q7D/�߻�~�Oi*p7L{jJ��0�pTU�OMk��`�p�_��������C��H��@V���rm�08s���!��WP��-%HR\A_����h#�6��Y�UR�����#�+e���C_����bu��@��c��[(K���GШ��M-,w��7���G��z�o�N���N��(x�:�}$@�,�%��B��
�V��0n��uBG�#h����\��݈�����zV�z�Ks-�<�QGEr���Y����_�b����(����{�Z	���G�@�263�22]�1�R������d�Q����732N8����yq����E�<Y��SY�B9]Q�6�ua�(�!d+�n��c�W���~jr&8�T�y\���E5o6��0��D��nd��4�5���'@�D���Jp �|[��C媟΢4�8��fYV�H�z� ����X�~�Y���!���G�mO��Sx�U:Da���3�s^���U�a��i�qq�Τ��r��jL�Ī�$܎hT�v�J�g�pJ��J�f�ػ���I�АL�oϻ.h�d�p�r�	��5�j�u�Q��1���E�&���\��N��$W�[�E+���g�n�`�W\؟.X���c�Z7=������^��M�uJd�Bb��{��G[R�9Uڌ�a�����g�����S[b9V�=�$��#Ѧ���CѸۋ�w����T����_��gD80 �_NNm���VH]��q��u�E�޿�#�D����q�P"F���P�[���
ݶ���L����)Ӝ���7�n�J�@��Ѕhb+��wǒ�����A�0/���#��?��:q!�q��u9��o��yH���Z*z���'[arڎޢ���UA�s���hiI,3���/Nr�&-���V!�oM�տeR�ra������fz]���~��B�QJL���Lph��=9�P*���T���އ �ߦ���&��u��Xb#�0u@XلQn=@��kCUV�9��S��y)[������G��iS�6�9��`�a�َF�ov�g�����X��Δht /�i����W|{���ѓ��U��O�`�t�Q�@<|F!j��ڶ>�@Ql����I��O6���yN�
��V,F����b7-�6�Urlڡ��Ș�bl=����2���)�0�)�f`���B�?��)��A��Y�bܯ�W���ܜ�����/�E]�׹�Wu�Tʓl�{yr�.x�����_S�d9�q�	@������!U�lo�rriZ�d���N\��o��j�A
��Ӷ�+y�}���f��.�𤕦6��P���4mA���J���8�o15׷ߘQ{����g��+B����f�-D���TuU��J(��~G�cͪZ��/�Ñ��*�w�

ȷӽ�3#{݇��El) �ԩ��P�I��6�U8�Y��]�Ԭ��u�7O#&F��Κn��x��T��a��Lپ�
j�r3-$1�e`�O3F*\��xk��|1s�j�P����)����W�9k�U��n��)^P!��;�w5w�{�8����ܔ_��=�t�pkm�?��ub�O��^�WSYv���׺�_��l�,Y�ȩ�pK%�U��@���-�PXQޤg��Kv��v&B��b"��Db����ֿ3����ן��X+v]���R��uo����������TQѤ�o�I�Y���O���"z���\��bF�I��DǏ��B�ژ����"-�}�|rj�����uX��]�Ol�o�ҁ&(���\wj19'��M�~�ൗ����{s��'qW���Z4b8|�<J�9<���X ��E0��3>�'D�t�If=���(_��D˵�>*���$�����+)X�Dɓ>N��goN����%�M�t����Ì�i�������`#��pYb��;���D�n!sdij;V�����_u����Ct��7��2��F䳦�4z��K������Є��gXTW�><�L,hb C�ĂR�EQDA@�h 齏�"
QF@� �m�H Aa�(�0 ��9�P�������z�"ל}vY�^���>� �n"���'�U@�ʾZ:v�%?��y��RP��O�WP��֎8`8<����5/�Η�㖜��'�_�a:ߕ��x4��"ںOf����{t�ݬ���o8�_=%�m��a���{�R)�ڑ�F���g�:T��(���b&������M��~]/��HO)? �-eB�C�W_���*������9t��S`���s23q=#�r��������E����M�:�W���d�<_�5��Dj�n[
�����X{&���c{�������%��,�oη�ǁ��Q�&�������;I���I�\H�w���|-@J�I�^�e~�Ț���F�5_}mi-6�'�o5Rג9��ۈ��Gm<�J�����d��x���,�Ǔ�!���ڗ{L7�ن��ʸ����?Z���&�����?���촡-_�<K�(_D��DSO�.��#,�:��]�'X�]����r%��ȣf���88�v��B����qX��PVN9��&������쩆I�0�}R���>���ށ���U˾E��X��E�5lv����������M%��eiE�ͫ�qgG�߁���cv��2�އ_5d�tD	l����ui���g�Ԝ�-E���j�W�*K���`�����.���S�/L[J�XK�d��o��� �6k���b��_��}5����� O��{��ek�d0�mW������=�'^�l��A��F��eo�5Aphg�Xm�0�'*�!]˞[�R�bd�>�Y�-̊z�l@��`�����}���>��,�_ԏ����gfLp�>�%�ī,�̙z�j,�ZA�/n�z 'Q�<��_c��eJl�hRIե���)�0_~x���|���=tl��ޗ�G��� ���]�7EZa��N����}�-y��:`��:[}K�} M�@�N�"��	�f~žڠ�;P���6}�}�4���/����ν�Ik�*n�+q�����=�l��� ']��_\=Gݽ%��/ᨹ8��F��kL�E1��d��:(.�w��%�l�M�� �����]Ăj��d1��fy��l�p�K��2.:�������U�����_�����w� p0o�֧��(Q� Ȧ	�����ꖼت���b��~����N$b8�nT��$�B`����y���h{�I��]��?�� �����A����3Պ�pG}�:�p���GŃ.Hm�8�� 4�F��+	w�VD������oF��׌!�.4H��3��{�|i/�S�j!V��)�I'�5P8fʔ�a�t���n�d����~.��b�X(��_۞����KY�)�P.��{�h4?�^���d��
�N���ehz%�pt?�|�'�EA�;Tc���M>��Y1���"�/�&&ZР�gao���ԋ�Hi��EL�?���DYc�;�f'4�
@ɋe�ɺ}�)�H������5�t�������������g���b���;�<� WՃ���noP<A@i�'��pbq"�jwN����"�[��ͳ�a��%���������]���/׌�����J8�p����K��F�����G9��v~^%�R���+�*;��W��N�f\��,�n�!ע* �_S8z�'��y���`=p(�b���mY����:q�*�/�����:�">}A��˷ѧ^�u��MU٧��4���?�M�iz�K<�~:��]�?E�l�,�HE�.�3�����2UZ�;�}z�X�����Gf7�K�jX����ʲk��	�3ypFx�|-������D\r[Oe���vԄC�L�u{�Ꮏ<:����^I���{(�O�m��9�yth�O>6�	j�~��Y��np�}�9p�0M|^��X.����X��	��?��(�����`4E턬���.�+O�{ ��V�VkBU�Nm��k���3��gW$h�ݶٍ�耤k#�� ��ϛE��޹����g�oVs�����065�0�9Xv#��O��	k�}��9 5W�Y�M�����.[��w���h�\r)�p]F��O�M^ �tw�A"���v�×�0#�P��D�n�m`M� Iz���T���0h�����Ur�HQp6��7�\wo�<�TB#�O��q��U6�����,��znE�_([�G�L�;����ǯ��N����paW]�G��	$ɜ"��%�;��g3~ʓ���K���eb{�p�숄��yW������(H��N�����p���D��ǧ�׽%��_���p�ǃ���|V�P�~��k6�/ݓ����?�ޖosd�5��'zڏSv�	]�s���v�����*�P��ۈw�P/����vן�_�zۉ%�`"Ur��h���x��J�݅I�K�vd��qw6	%�H��B�n���E��˚���;TE@�S�D��M{t<��I�&�V�����F��
����u�����#�J�����A�a
�	���6��N���c���k��k^�X��m#¹kǳ�XڂMBW��{_��_C>Q~/���K�g-K���� ��� �&�r	�G��������fzP)K��;D���A��a�9ɪH�q��|F����O��r��3�,a��3�"i<ǵdP�ZN���Hwp��(+_���=�����ˑ�7�oSqr���dm�+X�T�v����� �+�={5@"0?�+U��ܕ�,~�qy�
�,y����>�0�܂ů ��'�AcQ$]��ߢ>?)e��ζ���uo��,���kk@�� �Zܾ�����$R�B���/Yso��;��D�BN{������2Q4g�/������~Y<B��kO����GQ������ϧ�g߰:��?ڊN���q���ώ5��;��9�+m��yK������L�ܼ���n�r����R�D{������C'/�n�X�;����;����;����;����;����;��B�9�6�R+��л\���^���R�pE��͉K�..����쩝�L-|A�U�v�ԓ�z�E�b�'�%v��7���^�˭���{���{5�ސ�CGVZ��7l������]�#���gҶI$\{�LHw#ZY�c��YI�Q!���5x�H*��n�L����ZH������˓�2�F����H�݉yVf�n\���Cs��"+��u�_c31����1��59g��_К�o[ۚ�E��_K�NL9�ipTCz;6���s�؊U����չ�9�>7��\;�ҳ��h��Qd����T��엀�t*�0�X�Ŝ��>H��A��-g�t��-��5#��5U��ji��ġ}����ڶ��~700�Ԩ=ňgcx)����4�>�0�9����1g�,�,��Ф��ϭE�@eW��n�ų́�w�	��~^�۝�~�`O/�R��k���w�㛨ў:h�����ō���bK������:m�(�AJ��F���Z'�/���G|=N�̍���^&؍��/=7��Ԍ��^�D�@��r3�h�|��G��|�>��a/7�� \5������2�ǱnV,i�	[���p�# �m2�4�B��o!�����	��k��ԟs����;rK�ml����er�#2c%�R���̹�x����&*c�G���a�Ka(ֺ+1����u�-�D���^��v�z�ў�6[�٩��Z�}2�VIav��E�;̍�A���I��w�Qsʼ:��b��.�� �^ݵ�3e��p�թD��;i7n�X�pw�d�o$�NZ�9c�!+pv�>6
�Cvp韮�������y	�I�#��H&����VWt2_:��1����F��3�a$�Y�Q7�C��2��2!v�LW|� ��t��v�;ג���l6k�R`Ppg&d���φ[�:��������S;�xǟ���j��[v���¹�Bn�V�Z�l�dH�GG�9�82��ue�w*C�2O��p�3��qj;����qP�ZN�O3{zR����-��+�z���n�[�F_e�AO'��|.E��M�!n�K�M:Ag9S���F�?am�1�rN�α�8hNJ�_|�]bE��{�n$�������#}ֿ<�=�>�(�����ư�W� ��eN�Bz�F[�#���t{@�����,.sl�+Q�[5|#`���Vy�"�-���=���������ߧ"�=:5� ZX�$"���9�'�{۾���4J����nΗ?~�reB���pe#��0 8(�}��a��֩�وY����~��'�2ݹ�ΰ���7����C���|�餬f�抿0o��&�ٙk���[=��\� �u`7X����k���_�y'�>N�3�v�x�XH�I�����e����GK�ʿy@/uo�����pj�������'�_)7~ҋ��M*�՞{�-ӱ���������ý�䴁�T��G����(�z�c}����LR�@\�j��TK��LS���/p����������-�:~�w�����I�y�h�A�N,q6]�E�V�]����xt�ˀ��m"�/0]�T���70��5��&]��Y�
�|��&N�.9��Ck�mk�����dT�⦾Zց��Dh�E�ȵ�6�RZB*�+�?:W�vs�q�a<Un<�����0;�/q72��κS�Y��t{��}k!�V�/�k�w�St��$f��6�<> �pE�3�3���h�����Ў����3���Cu�[�����F��7�Gb�{ҀF1O�tmT2RʉM���Y�:�����]����뻯�A-X��?-l�w�[�ͻ"T�$D�+��.^���� ���T�����
����3�`�a\Xf9�=�k���و�^��@�*�Aѿ�	?l4D�_��/A��Al�{��!���ީ������n��Og粙�44B��	�@�3n4���jh�$y�������bi�:vƝZ/f�yw#��{��*?#���PAN�ӟd���KH�2�~5��ݯ��OJB�� C@+m��+�3S_��C�j�)��T���{��9T�=l�s��zK�P��Y�kՋ�����c^`�)��W�����b�]5Yr�C�:1%�6,�Ӗ~*���DC��
D�Y�Hj�o�_��xd���!ڿZW���	�G~s��'��a��I��NP9�'�h{�q:�h09ikg!�Vm@�=_��R���ݛE1�$y�&L�nu�3�=�og3.��A7������}v��kx�	��RL���E�I陏�i�0�X O�� Yr¯��1�¹�%��1�P��.|�}f�)����vZ�~�|�Z����ִ�*v;O�6h�vw�dP��5
���t%:�|ZC_�����80����Z<Y�A��e�zB?x�iwGX�7 B�yS�M�{ib�5�7X�@��}PS�K��U}?��
sd��4-���N������Uv��̼߂\h���A����I爙��N�)���ߓ��+0s>O^�M<��"��9���0�;W���#��фi��9���|�B��"���hL>�2`�E� ��S�A#�ؖ-��J������l�U{�#q
u���ǟ;e�x��A�l֠~9l{=�Um�Q��?a����e�]�͙�S�J��NF��D�O��z.�n(��:X���|�Y�M���>Y>�;f&��Xg�+�K"����O{d�ٱ_C����9�0G�m�H�����0ˮc�'m\K"��H���Z��f�/���j-u��ؠX���F:*o���3�
|J
�*�O5~�H��r
	�=�?Q�[���9$H�Bb�هC&��Tv��Ǳ���T���ֹO��c
�4s����/�fm9��з�F ��k"Ǣh�N��(4N�.�㏯�� ٻ�Dd�)��'�Q^�>^�ItJ}�P�;�^:d����.���m�ԯ��n�+Y�4 �#k�}[a�%Gl�Q�v�q�£�oY�REhc��=�q!r�C�|��[�`��Q�.����q�6Ŏ����o�q�-�O�q�)�3�H(r6���Ab<.�A�_&��z��˅���t���&�jBk�ܴҌ�?/_�v3�1���Wo�tѮh�<Y�zKt[��츽�F�3G�T~�_r��2�F�!)W��Ls�������!eR��c��n���p�:.Fa�S�=�/�K�F� T��#_ـ儼��w3�:)����3�j��L����)	}��"4�m1�:<9ܨ��ѓ)�N����Frz-4�F����J���X���E�}oh92{�N�1(����T\}|�6���K,αj��m����E��FUJ]�hP�A�t�k��{|�\�GP>c]�6���J�F�R��q�@n������c�}�{S�Y��pr���0#@ [Ef�][Ψ���G2ػM-L.�~�S1�u���]^�q���hx���p�nޮ[?�ڰ"�]Z���"\e�Yy;�f��<m�Zv+.uB6<���:6��+cl��Wy�xg�JYde��}�I���x#1���O������#����rb�We��.�=�/�<����U������m ��+�+�\M�@��o'���zųo��Z��19v)�P4��N,{�P~��X�r���c��e��ϫ����c�B^��2�p�I_/����©M��Έw7���ƙ�柜9�w�t�jA�L�o�O�3rm9�M1�-�\��NO&�j��X��oOx�L�o:���e0��U�J��� ��c�����}����{��QVME׮��Z����j~��k�\P7��FUM>�U=���6�H9Bp2kcu�*'����6��ߪ'���|!���av��v`�3��zˉE�P���5���i�Roْ=�	�&��A������#��ڜ_\��a� �j���cg��	%��x&n'ì�'&�O]`b��Sī�]�(
�(6N�c���?c�ާ#�9f�~��k<c�b���2~�b%�����a x���oS�bsŻ�:�!�z7Qǧe�{S]S�u�\a$4�Ӫ䔑fw��=cO�ZU����E����6|���
ob,��Jy�*{1-��}\�ݗ���B0Ҫ|�K��u���/��N�G&�;F���m�/uϫ��� �p���5�;�{8L�,���N�*T5ɢ��C��VE�j
?�������p��t��ޯ��_s3@�a0gR�79s��q0���v��V?��ԏ_@�$U�w����X8��3+����}������$o�V����AN������}Op���j)�g��B��������A]Ǽ�;������)��p�xu��H�~���/�H�:W��N({���(���ۛ��N��Cۻ�N��o}�e1�	D�"}6�(hv�ޯ� \����&�?ͫޜW�ܦxE��N����Y~HF��s�֯���;a�+7��\��Y :C��+rW������I'[�����i#��k�g�E`�QM��
q&:�
4�-a���\%a��i+t"����u�	i��J�h�$l�q�y;ӮwZ�?ڱXе���h�,�U*�� k������0?h�%U��I�|!Q��RT�����3	2��T��ɌšMá-�o\��+z`�'���b�Z��X�0�a�O�ݨ�<mzc��Gne�;c�dF����%��
�,�ыQc緙��5��ˎ����SS�bw�5_���R���7w�)1������,^j|�撡4�i��kۊ�9��1x\�o3O �n�i]Y���	��</��99��ƺ�gbL��(ur&0'�?��#;�9�k7�Qp �A<�x�\��=`R��>���beE]����[�2��)1�>r���.��_�W�ɕJ�| =����ޏG��j�f&d᚞�`���CC�T������8�#��t�V2��T�xv�wt�xX�q�KUE'8`��ܛj����!G�i���&?a���{��i},fm�N����F3(�و�]D�:�Zd�>��{Ã�;�	+rf�_nv7��F�*Z8��Z?S�@GI\��xȃ���`��R�&U��������6�8���O9�����5��%!W'���9 "�����t�	��|*���@W1�ZX�f���en\	W!�����Sl>N��s �t[�����M��T޻;��/a�\O��Z.OȞD<��9��0��U�<9�XR8;h���cI���E2�do	�h���D�� �n3us�ޓN�Q�F��)�I��U�"�����a#�Q5<��
L���I̡�����&a	��2��#���@����p��dt�b��w:Gz���8oº=H�M:ꉸ=�+� Q��!1�5�C��n��\O�0��#��v
��Q��+B���]���4JOy����==O�'U�e �\`b�[Mǻ�O'QK���3���P ^=1�JcxL�ĊQp�?Gd�m�wy��nl<��,1U���Hi���&��eW�m@��<e�l��X�j+38�[zSAB^@(�f�z<�]���L-��\y�{���C����M�����޶�gW�Y�$t��]�J�u��o�C5pvƵ3	����!��YeGu~��
�jά�C�*[�;��@��n��8��*L�fv6�(�st�7��{�R�?\���BܖԜ�f�ޛ�:�.��]Y��5��I�3gRZ~��t��������R�k	�j�8n\��E�نǜkl9�<�8hS����|Y�$%5/p~�X=-�d�M���OjT<  ;�;�Ie���	{�um^� K�x��/2�ᕹ�Xc��ԣ�rbc�q�`�ź�K�*O�M��EI׌�%ݻ����C�bT�	���B�vQEHr�Z�(��J��W�Ai����JE�%r���Y�Q?���!�&�UX#�1 �GWd�ťJ�߫P�����<���v��s�\H�vr�N��Tz$�j�&�7���_l�jdÕz��$& ����ح��q���N�o4U�s�qa�Dx�J<v ������@qo��d��NpN*�}�@��ݨ��s� � �!�D<��f�3L&�0/�U��f+Ф2��*�Վ�P����P�������%)S��ݳ2�N��*��XdJӃ��4Ω��z|�%ȯ.�y�΄[�,�#FJ����v)ԗq��M��*���K���B�?r�b��aE�:��ϼ�4-�Ï��l��6��U�A�.*��4�;tŕ�k\��feKd	��?�R����u���w��L	솨��I�������*��:�� �0M��ÿ/hN�����P��D�B���1՝��x/ɪ~뎃�K�%��8Z�u�X1�&�4�D
�X�Ĺ�S��E�04ST�đi
���� �u!��IS���=)rB���2$p[�758�[�mT��1P�����fQ7�O�C����z0����;�ô��?�H����Z�cĽ �j!�(��8��jTUX3��qj�/mHID��Ӿ�?Y� 8K1��0��d�;� ��a�������;����{�^Y�܆�K����Iԓ;F0�w\mFRj��M����������{�Ԍت!�������
{!/<��,���Ow�}ε�����-�9�5�C�
�>�LK����:��퟼��'U�`y�n�HJu�9�l�nX���zѻ�[qOR��2{ȓhIz�hb�O{�#�{�*{�H��ڍ�l��i���F �S����QHX���l4��D�"b;��3���ح�>-�f��{p��ղ�Qgs#��	ĺّ@�|��[��s���P�h���ȡ8�����P<'Qmv@�+��2O�I�wJ�ЇK� }n�����Ӌb�Dj_ݰ|��x@)�^���j�h]���%$��?�L� �7@�g�����l��;������sM�$&�D������������.�<�N�b�K9�D@d��0��Q�Вs�Q0�Ks����t��t��HمF�
P���Cn=_Hf7������=��@u��)̻	��T�E����:�kR��{���{C�#��H����J�:1��f�������T��b�Ԝ:E� eD0��~�U�4�.v����_����x\0x��HA�x���g���Lħ�b�H���Hl�B�������{x`M�Ԣ]E�Q�X��&T�>X 	�?׵d�+��O�b��5Z`�.=�mW4i�Sh��%y/�_UZ�~4)?�~����")��c���1�`|CD%oS]S��W���n8Í+i����N����-��J�����k4VP��M�H���E��`�z#6l�],�ݔ�ک_�����Ǹ��7����f3 �.+qvY,�ǵ��
�b���Ķ���K���P���b'��j2�@-ľV��-���AF�:l�U#b���+O���z�j=r\5�a�c�|U���kP�ͧ9�O1!B�.RHw��Y�T���r��.($Vp�t`R�wp�l�'"��6�\r��]�/�4e��3�$;NW��8�k��E�hH��嫆,�*��X���bJ�)T���7�������3C�Č;>դ�a�#>-�~����/�������L�@r�LS�Ѥ3Z���-!E|�Wz]�g^��A�ɭ�k�ѓr|1XG��@����rE��L4���n�bQ�;�Da8�H�Dq`d�,?t#D�2�q���Gy˅��P�B"SU#��ъ-��B�
�'b�vK<����A�~'�Y�x���bLM�"�p���4�/0�����*]�^��M��:��WI��Y�����9�|�7n���v����PlZ�	�E�)�����J�خh�!�.����u��@�Ƨ.BU!�&߃�g�=�؀#�����h��뎪��>���*�L����*g#��w�[~G�!�q _�O�{���y��!�#���(��]t��0�Jޱ8����Dy4�� 9�u v�W�$����/�&�w��k���,���"Ƞ��P'~<��	�9X��H�}ha��yɱX��73:�����x=b� �mF�?�y}��F�
@-��#�_IoC������l��`c�����GAZ���[�J�69<�ħ�����	bM/����=�&�pT��(�ina��=L3ڌtU��nr���XЄ8`�[TCSD�x�i��C���zİR� �*��s�l?��EzH`��4v!�=^����|�-�(8��oi�[�>q9�13��ճ�*ԙ��fe�3���!�� ml�&�ˍ��V�Ux+%%�8r@r	�K.�/���v0D;c?Ym�?��b�O��]�-�)��P�T����=��u%��h<���\k���㊍N�̃n�<��M�r��O�:&s;}�g'�_�ܧ��*�2�
�7���'�!�A��m�/fԫ���$e9���X���}1w%�I���1�О���Ze1�ʉw5��?�\D�,��!���.V���W�x��'���m�=���8��ꨶpi$ztQy�2�b�u�j���	�������n H@���Ć�T����?�A&ʙ������YC���Ƌ��W�[�7Χ��Id�i��H��'����
�Jv�_�+�:_т��s�N�W߄���2���箻?ps;�f��˞�_?�iX�{]���
V_�> ���"�]1RBX��|+��h_���Q좦#�eT���#3�����Wa���{�K��
��Ox�����9M�R�@R�.ު$9�L��ؘ���8��1���RO��1�e{b�`T���DM������-�>B):v������.	��T�~��t����.bR����g:h_���M1����J^����oa=;���7e��U�	�A;I���l����������9�x���mΝOgC�h����/�@��i�t�]T'�3�Yp)�E�ʳ���T��=W��0[ݱ��g߸��W�u6��5�Q�xSG�����W~���s����ݎ��ݼ^[�D����e�L���6�مOo�wk\���հ �H�8PE:M%g���^�V�~��n;�ݬL�*C��n�TNb�wL�~]�ޘ��g.�?�E�D��l��XRD?3E���B+�(3���t�w��y�a�
�[����U�x�g�;����sg-d�����B��W[�
~+^���b��}�I�DYH�p����T�,��f���=�+^̈��ln+�rg���s��S���f�u7�&��PnqX%��\�H�_�	�j�[�u*��i��e����*i,���P�O�7��(r�a����AO���)9�&�'N8t�e�}%z.���HUU#����O���8M���7{�q�.d���?~Ζ�r��ju�wy�E�<�t{��Ā�h���9#�I���]��G�;M2J[����S����)�M������+	e6ӹ7�6�i���T����In���	cnߌ�g����z<K���
v{�y�2��5��~t��!�hF,t��vN���xk���}�� ����A4r��n�ޤ�ӗ�~|o?�w*�H�q=���&�hh&��Pf� f>eD_O#����Ԉ��}����ĉ��w�!������ښ��3Sّz�p�a�q�b�j&~5������-����ə��S��h��%��w��0�����0�
��������I	hD?����,玳�N�-�1>�����S�Nhq��ʏ<�-��77|�9"�AvIi[�Ą��6����"|W��z\ko���W�ig��p`�gN�Ee�JͰnL����[%�I��c���݀��2�v�����^RzN/`C�qF}tq���	1bV�]�ճ�2x�2�<��)8Uʢ��ȼ�l�IXe7��D���Y�b��8��;�V����kR���ӑM��|t��� ��ǹ'�<ث�����5zt�K�E��������;_R�-0�;�iD؉ن�Bu1��8��tiLb12D3�bR��q�dh��Z�-��w����ƺ�:���^1D��eK�J��4�j�i��qـ�B.�����A��Н\+�XJ��}tH����&�ﴜ��D�JM�4�Q�#�A�!�Ik_�������Z�ҟX�k��5#(~��V.�=q6��D�X�aR��7�l<.<s���jeg֗j�H]�a��a��S#e�m�����Giq�{��4�gΛ�|��ȧ�8�5�]6�O�H�aN��ե�F�iF����){<�o����'Z\���8<%��L%ݓ�'��G�)J�(ă�NSN���s�kxs����M��2�_�RǦ>O�̊�3G�JC�5^_������7~^��S|�A�����hj|8kب��N_��i�3x�>^�ӕ�<��W�y�2�a��cՀ>�~;u�ߎ�B11��85w�1%�k���z��-.����q��x�@.�7c�}��P�0�����\t�_J,���g������Φ���~���ZCӭ��3�[�$�f$��ˆm��S�2��
	G��g�he�uk�?�.oz�<e��V��Y�f�}�l����Q�r����Z�9�t�ԥC���:5j~/��Li��7��X14���N�U���8K�l�����a�D��^޶�ja�z����Ϩq�Z'�Q������x�0���,^�{��>W1.O�s�3a�;$z.�L{sB[�O�]����Jn_c��D��F��N�c���dn;�s��i �$�]�D��t�3?IMm�5����'�V���:�C�b��u��޳O:��f6��Zd��C��E�*UD����\e���/ic_��#��������W�w�::n�S86����U=�[�`��M����'nz=��;������Ѭɜ�U[Vt�;+�h8*�W���6C/�O�Y�ki��y�)5z��H:7zK@��~����sgL���)YO�<ҽ�
X�7m3҇x�t5b���g�H�r����x��'&AP��ӎ<����TƁ��%�[��v"xؕSy�uiI=%��/�IQ׭���7U��,]�v�_[&�N[�j����F�&�;��]&���}��T�͋�g�r%�^����mf5g���҅�6������p��(�������2z��_Y�45s�7�iތ7)����`)fܙUV�|v��=j�it��v\�C͏oj}_��v��.���Ok�{L�59k3ئ�ڣof&�x�g��y?�Ꜥ�^��qj��.ѣk%����]u�<�ˣ�݌wО�i��%r���܀���	]<�n��GT�~'�'C�}��௉�Y�NcA��p3���l�^�?�G��Tk��Ӗ����i}u�W_��}ȇ{�K/fS[�^Td�����.��gƤq�i)����6���O�ǔ�jA�v����x`��
�F����w��4�׫�L�Au��Z_�TI�[&��{r;����C
B����i�dٴ����CXu��)f!.;vX�n���u�W�a���T
%�A��0B�mmu��A�|R*L�+�흖g7B�QӔ�'v5	&V$�����ĸ���P|Jې��N�9���47ϭ��B�"82i�:z��q�Ln=1��9>pI�ً��A�ͰS1z������#���Ǜ8�P��>x�X�t��t�Ha�Lh� )���#S\ǈ��2�����^Q"�˞��1߷�޼�����	��}�.�Yn���%�^��d��FI9ھZf�ս?�oݟ��1%�(jk����w�sN��Z~�����HuM�!���X;}BB�Ւw�?LBѹ�xV"q���7�.R_&m]�	�z ��J�HC��f��g_�cB�=}�fH,�Y�;nS���`1Z����
��i��Qk�m������`�X|��c)�8RtM��M�D7����qW�6�ԫ��;����d�ѺO��cv�v*�!X�}�����>m���c|���zeǌ����C�Fx`�@��� �3��Rқ�L���O�T 7�e��@�H���j��,%��O���wN�􄑆�[J��ќ��8_�a�vwS[��r�� P�w��O�n$�G�|P90t8:�y�����׽ 8迪�Ć��!���;?��b�
i)���d�Z_����1�r�T�i�pvӴ���/?�@s�[�'󴴟f@Y��4�G���hJC�N� 8��Qn��jd~����0��gM���!�H�6�ޛ�]w�y��7'�#Q�J㾗~�U+cf�|5`�Dt��nN���0�� ��j������@h	܉>�2��{�ĝO���c�-���k�Pa���� 5w��B���9����ѓxG"����a�~�l����X5�Zp���>�$���'�b�w� �~�5��w�^�72N���r��,�L{g�� �Z��z�%�N;Ih+��M,��5��ZE27�B��͕I�hH/"��9���t}��b��РbJ�y�'�A�ɣ\эJ"em$�'��!+Ox�D�+�x#���m�zQ⸷���i�Lþ���<��~�0��U����P�*q�+M�o���*gAOM<mکA�Fm
�m
GZQ����}���#��=1u/B�x:�L���?��)I��CYA�Z��:�쾮����9.�Ȅ��x��U�iڊ�R	�|�$��:� ���O�6]xo�߸�Ï�|F�SYF}��w&�Į�7�N����XW?�&����-���w�}|�9!:5tLc�˭�4�3:�DY�X�OSs���d�z8�(����@�~Y��HiL2D�j΢%��b��΋�I[$<Ɠ����r f�o���M$����bD���Py�����C�r�x
���ף�� O�~/mJ���E�'����@;����-��jmN�į�B(aH���V�2ӵ�Z �:�a48���c+n���!�d�n���WD�_�E>�-K���S�-�:Ϛ��-�����	��(1��y�S����bP[sZ�}"�Cщ"��wL ��w(�`�0��o�~q�L1~e�z�����i�𴓎"��(n^��%�S'��_�<A����\�Ͻy��?Ag�ヱD�A9�^S�G�:Ju����RPұ=غ/�/L�s�����L��4�CM��� E��ɧ��������K�o���PDhHޠ�'��|��Rb�}�{,8�~s�wG~��g��Vd� �nRp".j�麙�ŷm�L��ks���������o�)_�t�f4Ppx��O�D�=]�f���K�H�1;�b
�y�|@b*����r�Y�w��\��������!)�Qu�PU��Cż��:�K���:k�?a᠂�
Q������m��[�^������oy%^��ﾚ�Šzg�h�_'�����b�-� �y9��,��o�[�͖H����l�·#-A�ߦ7i��9H� KE�hj|��?/�?H�]���x ����{��i�Sa̋��_!����J�R�߄��3�(�/�%�
dI�f��/1h�3���
'�^�b��1���L=��S�C�Z��L�-@]�F�o��݀S��8EmJ��r�nҳ����lZ��B���1y�cXM���A��qn�D6
O�CK���䥶A�]t�;������߇*m�"�lz���ܥ�/)��׋�r
DU�� _|{��?j�7P��+7Cf􀄅�HT�]����4��~�qM�|R���2
�����P�� �-�zu�3�a��х;�y���-z�M����QP}��Eڀ'�������$;G�d�_�X��A�߰V�f���U�Η������2�.P:
*�;�%��I�˨٥i��bZ��X�Vޠz_�r�K��6��1ZY,}�#�H����c��]w�3����	R���/5s���?�Ca���6�b���%^9~^.Jغ���-��K��1*C��r�'��?��d�|O�����G�K)�F�'t�S��ρ#-�ߜ�!{���9��ȇ��(n�)WE9�6d Q��"!�w���ŏ��!�Rɞ�~u��qv�¿�Wr~�^�?n��X�4����Mƙ0�D��Ma��죋���p&5w�Z>^X����.�

P�����Re�j,�;ӘX��`�1\M�l�p�ͥ1ʙ�q��czm��T,]���$z�F�tN�>�η����R�]_���/�1��fw�\xUzTN󕓩4�=��Si�2�>�L�E��  �$j�Z\\d�kpL�S)��5�G��&q��%*Ei*H�<xme��+���vI]����Ћ
��n�D!,���|���X�XX3�vo@s-�׉����s�7������C�D@�H�
[?�G�giP�Y�yq���Przs�������M��:N��2�`�b%p�_�`�1����P����^�.�uH?�����_͍n����Qvs�m����HeJm�<Ԓ���W��y&��*���XH5��x*s�:�v ��u/�� ���BA�f�ț��H>&���"�\�[��6C�4�_:�8�mn���"C�8�V�C鞎�AG����E�dSp�sl$j"�X7p����X�!�u�W4j0���SƋ�C�t�j/pHã/���'P���?~gR/���#(�τKǻY&{���9�C�(7��_W��-NB]f.�X���O�4�ƧF�,�	�#C�	�>���Ρ%5�6ɋ���.�_r��K�6W�6�8*�ӏ�[��c�&��UK�'��y�]H,�� zb��;��b�a}[�ԜG-p�z]��~fڜa7e;�C{q&���s=7�-7�]��ҷ�g\�
ϗ��hR |�0����#��6�A:�Љ��#f��YɊGޝi���>.YB*h�g&�vX���D�
7�3��+�q��)����y'$)�4�{�E����`L�Ʒ���26;����R[��� ��Y��C�ݣ����RB@��v-p��:{*�4���_����ct�K�-q;��Kw�UA�D���ʎ4}�?�� [9)(j�JI�	 !`�.��i4���MJ~
�/-�����e����;`�f}�@|�Jm/{� �]��Y�H?��7��q�  H���־���7�H�R�Q#��.�ɲ���2G�=�z�ͦԽ:�/�@?��\B�~�j[W�Tж�$�3dnKpϦ�RNH2��¥~�TS�q6�>9}g��;9c��浲{u��3�c��l��)�P�s�~>7�J�͜�-O�z����{���\.�&�kw2y�����/��*8�?��>���G��?l���t��G���6�D���N��~H�����<���oKCy�5�9ͶMu9j#&H��6�FU���Q;\���(^�>+�-������i?�B+Ruͧ�I���X�n/�e���\�k9U.�yin{]3��d����D<opl5<-<��/$K���'y
��-��_@|��vU+��-�<,t�v����{��454TO��+��։#�Ɯ ��'���5�C;����(�*�v
	U��_p�/^F�Թqk$��
e����q����/3 eD�9���f���d:vZ��m���;R���}�]^�9դ�^Ȥ�5Ri�r?{�#�jؘgj��X�ˁpT3{5��|z�H��qenZS/�9���$ˁz6M�pL��ܸ���nB�\����N5,q����V�][q�vu%8;{���%d����bi�����^�J����ڋ��~(4Խ�x)�2�J�quLm��v�)Ԉ��`��^>��
�w�;��m�d�t-8S&�~�n�Ƀ5��E�>"? �?���%je�Ԗ��:'�$dHW��Q�N��>�:�O���C_�xb8Y�n,�q/m_Jb4��>1����R��W�n�ժ�N�4���[�p��<_.|���_I1N�zҨ�����-�UW#���Dee;����\�s��`m�B�������yt��qm����6�
YөaW�N8⹌�nj<|�ʧ�M��T�.z���Aw�n٩S��Q����V�G�V0�n��»�����d���T�i{"�;��ߺ�t��b�͌#�i�Ƴ�ۺ̞�H�� Vn洞��R�K&����ǃ���MU
+ٛ�D܃�o� �K"�)�c��4e�<%��p�UUd�Z8b�:�1�%���<c�[#��������G���<c���ItB���E�*�u�����+'\ E��磞�V1���.q0����=x�ў�����og5�yױe����[�:�iI�9�$��)���(�ˍ��~�v�9dB*j��v\S��C�⪇+ﺪj��ƕmn,�$#G�y�� � 4.�m����0�sa�2RvPU�X�k����<�����:G?�p�����<=��<�k�<�87�������ҫ1�@Ч+���v{��ԧJ&�{�y-���[�[�׻^;��%�X��~�s���U������\k(^���O�+)Ó�����J	6�0�EՃ�I]/��o��z�	�4�v��u��~�#Ovq��?�y���j|�S%M�;Ŷ��9uD����1]BjjaV�sB��(y�!G����x�0{��j#�� {�m�O��nt*���B�˼S�5������p���L�WӦ	��"�r6��"4x�����������J=���)��T���Z(2aZP�ٙ�J�Ǟ�bHJY�T�^dO�=��;�w������>��|�����?�Ϲ3w�E����s~��$H?t���b����3p͠[�C|�R�n&����ϗrf����#����֤�Y�'k>�t[	E�i�;k����{o���z̶���LG�zx��3�`3mQP�g���(kFڟPQ��{�=l����E����uLav�����w��=E|�\���0>�V��]��� t�>�i|RQilŸu^��M��� 3��5���H����W�Z$]���#�{:����a�_��.�S�[��'�L��� � �ׅ���t��^7/�P6f��Q����|�Z�	�/-/zn�N�y6�a!���`�%���}N�
��]x0�ňP	���M˛���~����ԭ�bD��|�����/"�#>�[S��7�I7��v��l����l�^�d�?`���J��E��S�Лα#f��y{ 8(��	�_�,�]�B�F�۶B��c��+�ߌ�?����<h���z��
�u��}~�&�nI^���L�٣U���ߚ�����s��RS�I]���{'ނ�K���җ�i�+�A����z��Y�:��C�����	%��w�K��kv����h�0��	T0�K�\ҳ	 ]R���)���ۈ��P82���#\o��Ex�m��2��z��9SajT��_I��m�B��js{��б�[�?�����C@y>?hzlb��g�U8y=]�T�~��<��	���u��B$���\�J��,�gb-�y��0'o�j���O�$�Љ��~�u� X������'՘���|����'�г�b+�XhD�)�ʯ|QZ`�Y�� K딓�6S`���LJ�z4��Lw�8�i�XRC�yQ�Ά�l����K?���c+;#�$��y��A �b��P��0%%����������AI����ATsQR�&A���K�[���
 ��S�EW����l�ተ���:�Az����aM�b�����^Iv�У�t"��&}��X1��o\�Dd׽A~P������QK�xE��G q9�6!�+��V<~����&%�#��S��<�0���a��6�]i �`2��2P.��Y��j{�I%F���Byվ���]���͔8 H��lR@ki�y�y�!󋜚C-��V��t���>�e|VR�yh˹R�x���w#"���<��<�����v��7�$hӍTr>y�_R�t�?hn�iܫ
,�F��5�q�4�V�l�Ƣ.�U&+��Y-AZ�7��F:���6�_��c^1��u*J�x�z���V�<M��
�������!�S����Ψ���/!`\u.,9��`�h_����_�";�K�}D�|��E~XNe�ê&�������T�������a�N�-�P��v_R\N��ܟ���e���
R�r�DHG`&�oJ6u;tTt�=�&��+�Η�@��}μ �g|wV�3��5��x�����*P��¼���2�%)3VC_������+ѹ�AMKa���s���2t��7Yee-��f�և_�bL'~�SB���ڒW~�*�[�`i9�qL����ҍu�b@�;g�j���#��쮈1;(���-lc�8)������\�N�aj0�OJjKYH�\�B_UXL�Á��ϧw��r���N���r�=�(("�u��k(Dm��b�K��N�@m'*m]EY��TUk�\�?^ԕb�?��X�{�R���+�FX�K�Sk 3q]�?D���`��T.l'@Y�dc�q����<4���m]�=]�+�Ʋ��FV	+��\lx��3������l��$~��4�I��@�l����b^N~Ԇ��1,�z�W���1Y�hl�j�Y����E�:�V���y��?��	���-F�y�A�4�<޺3�ﳟ��W	�^5^��;��`�l`�Y�	���?������y��ZE�9c�)-<�f~�c\8]���$|SE$�\�>k��#���PU3����Q�n����������A�S��BcQVh��I~�3^�4��5b|Z�~ �\c! <�e���p���R�������C�O�~�9IM�0_*+��u\���������"�YյH�!u5Ξ6E�|�Fb����"Ҙ��{���%Q7��ձa��VBmL�ɔ��MCT�0U���:�2|m��' ��%1c� ˵+>/���ޛ�eU�1���vv�T8��A^��P:#`���N ^�R�*�$� ��?ő�]���/ރ«��g:�[�u���sm>8 6 �Vt�"��>|
\��&����l���m���� ���U�ٷ��Yl��2��P��J�٥�nE�*��ف���	xRb&�.�@З�/�
qs�cR��H�f��������V��F[f�.m��'�C�1�m}syq����d�*X�y}�n�=v(����ї�	*�+Ũo�,�G���
�U��Q|D>�_�{Q�x�1V�#�Gٰ[R[��]!�����<�o�y���&�y��K��o!tN�=3�W�,�]��G�������|�*�����,]�equ�����WvhK2�8��U������ma���9Kګ��g�m��̍����DWn�J��f���0)��\�S�mR�u�b٢���v��L.�,}�X�`��_T\;�:�`�X���%M@T�Z<^U���5�&~�\���@�F�*{��nK%Fv��7���1EڻO�KP��7QA������4�ڬ��u��>׌�L�BM;c�5��|Y��Ľ���S�F|!�"g���@ꥩP5��3�vn������ro�g��,L�,9�DD��l���>�}�i"��Ce��N���٪�}��VPJ3�A<ѭY���ߩ]�	�����F��l�oG��w�i4���x�*��`�!I�V2��Ï��i&�5�|�g1�t�5]��3v\=�#�c�����@��ύ�E��hV��sޭ̸�g�nWqWūY"3)m�qm}���*�0k[��lB���1��=]i�*)���|)�Fti���Y�����{s����H:�ژ���l���/�3�L�����ըx"�
�?c��V������_��psd�uy$%�׫�W!���)Lm��C�s$%ň��}�q��<z��y�^��(L1zl�r�ӕ�� ���ۏ=%U@�9����m�הּo:��$�Ի�����W��uд�����a�`Dy���,|��8����M��*��cIW�0��.D
��r��"��Ct]n�<ba��cq���8�1m�yܭ7�L<�C��2�d���(�@�ׅ]�In��f7r���V�+v<\�$H'��0�י�[|�_�/�z��78�#���=^�T��ű�aˈ�r���Oa
-\�1��S�=�7Mu�N]$t��M��n�K�]E���̂����C V�o-t-wFg��\ي���I&�c�m���=fl��A�|;���/��ʰx�̈́�+�G(zDZ����Ʈ�!��Kym���G�7��%�"J��lw�����^�,Z(�ME�	���c/]J��I�DX��:p6�p"^}�[��U����a?�����u�[*��.�+��L�/6��ի@q_C���N�`����=J�7�_r�j��j��̎�c�:�������Jj���N���"n���;�����v.F�K���FW|<��K�W���H�}��:���� V�����&����HXGRd��-���m�0_���HXF�)�f�M����kI1�J]��;�w���u��T,ў��n Ԓa*��! ��7��:Y�ԧ>s�-�u Z�+��n�*>nn����v��	 d�%��K�h��ߦ.�l�t��#g�I%���*C�э�f˖��4�y�6��iE�ϡ��w�^	cB��C�V��O�ˋEm�9��� �7��t�>����9�u�����A�Ins}g��������`�С�R�8�&p�҈p��qхhw[?t��io$-�I ��W�JxlB:~�>��oj��~��6� 2T����O}��++�6�����m籟21��U?�Բj a�^ځP�\"�Ah���&�_��*��u�\��f���=�79��b�W�T��֠�S\���_��]h_������b !��8��j�@�Yӷwƺ.qx���;@h�G�Z(X�NcTI�l{\2�@�4t1?��y}��y��@�Dn������N�I[�7�i���h�z���/GPO�cߜÉj��HSI1���,�^�
�ng�E[Q/�ڴ��ϻ]�[����'�Ae!�{������nQ����w��iIc��F6�gj�H%��Hsݐ��ב���> �2 ���!�:�FR�Z��2?����C�Ŗ��� �>�K�G"�G�$�;�����hg��lz�]�d�b�]�6a����c��KK㖋�Αˇ�E�j�[�c�!��߄����Z��ŲZ���FƳ���H�OױE�#F����b����}�_9G;Ń󇾚�Q��ߚ@�IY��mU �2����yhK+�!0�mv*c���e�����A�?���!����Nי-�_2���cCҀ�{w�����+�ed��FI_�B2}ض8�{Bj�)��.OVIB�=W�gO�5�A�L���o�vL��/D��n�c��t2��^Vk�E=I�n��nש(6um�h�/z���>B	2"�@�,Tpr�\c�#��ʰW���$zt*��Qנ�lfatO��7��&���G��gl��|���M����pb�h�Q N2-M^B[��T<��KP���B_?����y,�t@��s����+��	��P�<���j^0��#Bv���_!���ā˂��K�Ϡ{�a�M�Y!g��=�L�ʼ�3_����& �m�}#�6��,&@2��*˘?�����-��2b�Q�HghI � @^V�j���D@���ר�)���_�Z]mD p������ ��sϰ4��µ�����+�s��h�/pr�)zч��1RXɎ�p��KV��^+�"�;���ا0�ǆ�n�p� H��c]r1���i~�T6{�Ģ����☖u�j+#��[H�aç�OH��譢x�\d���Ø�|^����<M����u���s��r�}��~�[ƾ`�E�Cf������k3v�*�z�t�5������J|�#w��b��W�4���>�g�3���w6b���}P�Of�������mOqX]a�^�o	4�`�⤹/J#&���@F��:	Ҧ��Hv]{ꂲ�M�����0�s0�?�ȓ�nX�ex�>�E�j��Ȳ���ai��=���t��/�Q�A.~PY ��i��3�FK����j�a?��r6G�FE�lފ1�����'��n��>�Z�e�LVB��������Fg1\weɶ��RY�6�L=�6��ʖ�D<F��Ff=�  T��Ā�#�@����/z�z���T͏���^�V!g	��̋��d��~�"1�np�x�q2hH���ԩ�_��i�$F*��όD|NWx�<�Ѯ�(�L⃘��F��񣚄��64����r懗�W�
�:	����- ��<2�i��14��[��� ��~^�Mo ���@��O���1�_�|SaO���Q�����n�*HRؤHS��ѕ� �G�[(��]u�E?�컼���:�?z8����.H���הF�ɕ?ڷ%Z�]���d�`�N\&�`�&��ғD�Z�FP��ʵz�����W�t��!/یZJh˯��+cL	�+{-�]9Ni�������!�v�./��
D��T�����a��@h&�ۦ�`j`I��z���%�7f�&z�k�b)���}��| L�H��ň��-�Jl��x�LIf̧��'z*Ǐ�.z�����?1�C�o��>�5�3�4�E|Dq��{�Y�C*��d^����*�F��d�		�%#���\��J�Eñ	G�?R�g=]����%�����ư�L&���!1����spf̷��|�^�m���C���c�^2[F�VF"%{�9#��)'��9#��h���/���PE�vn@��t����_4+�W�sd�)���M���G�	-4�Z��í�;{��l8�щ΀������~ʄcZ�݃\f��c�ܠ�]� �lBtY�^�1���C{�{�2�3�.��j���jYۊ�+=��!�/A;GS*��*��Cdf��he27��yx���2�Z�6���k�G�g�Г��x��Ht:}+u��ؤ�/3��49+�Q��V�ѥ	�� tR1�0?{BF�|~��̮�w/-}_F:�6�����Fڏ�R�=�pD�7�����n��=&X�r��G���B.F�`Y}r��K�v0oy��fgg�FR�;?O��Z,���Z4����e��6��q'��-M�7,�H�?�+�
H����{1Y}�z�o(5�׉��~�XB�Z�j���y��x��2Ԁ��P>Kq]��_ rG���t��xp�_v���d�5t4p���M�[�(+�����]�F?m���6y-����	�R.}�˷����(��6��zKz�� 鮂�<Pu5+�=)�ȱ���X�O�/Ͻ��8؝��67�+�s�`h����ݎ����#�Y�@��3���zt�\Ͽ�3v��_��~��[��%���@U��<%�ީՖ�衡�X���H����	$-+&��1<Z�I1 $��s�m�M"y�L}�����R	7	�_��2���+�yy����	�
8C��h0��b�?� 擲�b(̗Z��
P�YEq�!ꀂ���������G���&������,���XVAb���t�c k���H�5}��c�!�>o��@��Bep���E:��@ɿ����S��>���Q�4 �H�z2蟕�;��V�!�ד߭����B��Ձ�r��ͪ��W�@�|N�y��Xt�#P�y�J��Ϊ����D��\�#4�|t����F_T?Ot��̅�k �ߕ�)���dI���'�V� X_T|���2.@��iڎEר�����a����EK�3 �!ତ4�+�uk�Ľe8���{��֙���#��V0d� d�]�����t${Z��:���^MEU�[�8un���Xs:�Ջ��*.�Ry�"c���}3�����?`Tb�K⟦�!�҅��x's�c�RoH��.jI��,��V����iԭVA�u��n(�=.2k�2�\�:T%<� ����|������q���]�Kn
5���|uR��������!�X�Jg߳��"[�󬚽|���]Z��p#�z�.���ֻ'fe������7~�#I?�*/�0l�$I�s�G*sZ�ж|�/�mz����w�Tۍ��3�@P�*�q���|���f�h�1�_��RCR���d�ze�~��f�̣��y]I9<a�zX�][�gq28�m���FP1��5��>�W\��O����o�߮'ޏ0_Z���e�m�I8=TV�9���|��X��O��=��s�삋'������6vL����w����f�]�Y�P���e�vS�'ob���+4��u7N���uZHɡ]�� ��0XX�Ǡ���,�ʙn5}K�;,��M'|�.ZD7���l>�K��+���45���Ռ�.EU-D��!���ϟ�Ħ������h��u�<km'~��W�g�_b�r(v�uZt��歺��D��!W!Ϲ��*��ے9�W��f���G�q�!��z,�~��~�k�_�o�v�2���*x�^�Un1��\A
<p�Au�O��&�1!��]��!)�̙�s8$1�Z���˗���E!��_A��ӧx:�?,q7R����g�Cٗ�!��5�����{aR�e֢!v ��>'�:窫p\}�6�Y�$�hP���L�/�Q���r�쁬(��i���(�e݀/{[ߧ���6��2-�9�.�@�8��l6t?��TM�.?��|�yb���بݜ�'��:�e+�i���o�O^���(�h�'dP����6?�Yup����l�%�v���<��ݚF�K�}C#����0L��)؊1�ְ��2�t�!��3���n[�Rt��P����x�U���(�-�����F�Žߩ��@�.�DbT�=���R[�(b ����G�g+�� rd�A�6bʿ��#��sd[Y��p����@��^(s�ݰ���';����ӕ7i���Z&]��e����c6�L�!L�7�c.yu|�K�_
�IpO8;H�&w�RR��]u���.i@l|{��^�l�Wb�ǝ �*Jxա�=S�> ��:-�Hd|�A�пX���,���S�n�u��A���uT�"u�(&z(q�?~nz�,��|�`�⠽eXU ����w�,�x�G7������c�`Q8����|���huQ���g��i�8��o��� Ф`�ԋc6[�����&�l>C�����&�\�ͼ<rIg��qK���u���c�=U�]W�θ�������X0.���Wn�t��ݜ��(���z�����c�K��:� �������}��^�q��W�q�$�+ƽ�֨�OkM��i5��F ���g8�޼}�0��9=пZ�Cj���;i��������)-����� �$~�H�)�-tBr+ Y��̟��3��1v�0��i#�Q8���[�7��F���o�V�cA#}�����e�6�.�4E�X�� ?��1�MwD����d�O�]�^[(�����[�+����Zb$�S���q*�˽=j�(A{P۹F�v��Xi�,�c��ҡ c�f�^��ÍP�W8�im$5���2��rԄ��rY�(���A�胚Ex0�=fC�����2��¢�*�@*SD��ǴjE�Z�`��W6pV�N֫�-��~@��,y����i�U��W�4�fg|���E��a7#A�6���3��ǚ�c�u�q(��sh�F ��x����j0���5�9��|�ҵF��o��@z5x7'�� ��߀K7���[8E���S��r�%�cV����UK��s�����/��޼��r{���`��i�s�(�n
OԖןb��-e,��^
Dmp�1��؄r�j��=Ke���r6̨�wXy�%����8�9cQ+M�� a��@�����!����� MB��0�3�n@�� �������\L4���O���	� `�L#j�oO�s������1�X�clP�
�~���j�� v�x�R����oe�{���YQ�{1��-� Ye��N�O�)�F`�O,?�~�����sg�².D� 3���Qmr4p5�!5��dX�Ӥָ�F��N��%b��;��jB�h�;Z_ؽ;J5@���];ʃ�iR�5��@W�X��Z��^��j��W�c�é"j�G��9 ��2Şog�.�J����l���0)�P�r- Q���X���XH櫿?���&��P�V�RV�4fz�>KY[Y�Pbݺ�"�Ŷ��"�|e�8��o��
x2��
~H�4�!3k��ӣ�Ig��c���.̽�-Z
Ar`k����OB��-Ɨ�����c��f�3~�̻���(�墱�k:Q������&
+.:�?���-C�CGD�7�1Q�7]�Ӿ`���m�h�$a���Z*�xr.�d��
�|r�O��̸�tb�������:w�[p~ ��|�	������B�n��R���F��?�,M�حE/���|�h�7��A�e��٭�_�Q�#6�{�+���D�}��l:&�_8M����� ��y�}enڃFY �liU�~q��򩧫O߈;��r������Kο�pC��kL_V���Ő�8�p�3�3a�gZ�g����4����y�:Y�U%�E�7]{�ia�5E�c��y�_Z��D��w�ȳ�@�|�^���Z�M���S^�h�ݥ�|%�����c{E�S�_�[^RC ��(�,h@j8�����5��X�g�' P���qʓ�˞���Q� ��Tw��\�N�%K���~�E�6��c� �.��{������j*�G&ت ج�����d���1S9ț+��9e*�9<�.�,�N�ݥ���+;o��(��e�|r�y�L&v=g�f顆��]�-K(ڂ�*S��SB����}?�1�
`�z���bI��R�!ȑ��8q�HX285�SC;KV8�%`�9���qdl����5���J��+`�M=ʳ��/������=�Fˏ�����%�<	�*2���x���[��b����O*:	�C����m�%�4![�;����-�0Xt��P�iE�4[
H����L�}�{,��~�!n�5(�җ���aO���Г����$�
�!;��U�\��e�N`���Z���'� ���:�,�!�zNw�_��<��>&X�:> �;�4�N��}>��~��Is_���/|t�1��{�<��W��p�*������vtk,t�x���]�c�f�;��y��1O��@�'��-�8���-c����*�oG��4���M
���>FЇ�� �K�h ��a��%���7r,BZ�K}~0 ��z�$0?��q�_ve�94Z��X����+�^�	���3rB��z��;n�V˼���'f�&�&�m�����3K�7�i6�ԝ����������h��,�LY�w��dA���N:Qg?�`2O$�H����M���A��N����0��:���g�P��V-��6��i�u�0�����T.�AǗbHf�{�a&��Џ5��kӋ_z�%: Ё�������}Q違1��˳���d�p&n���(�<3����B����gԯ��՘�Eۣ��O&z�M�4����f�p&c�dcy]�T0Vy��!@i�MF_�Ͱ!�2	*Y���+΃V>�F0����'�5��:Fa����5�7z|v��B0ܩ��7���6�X�=զ���F� `h��o�T�[�(�~m~�L�߳=��;`<�\%E���-@� U�(�O@C��~��S�?�`�B��??6R3��6 �;���$Ւ�߶u>*���W�k���S��ZD�c��:��"*�SUI5��)m���3O ��;��AR��װsz���1 �T���K�C=��9Mb�ƅ���|=�c�;��y�{5�<�~v�/�� ��O������@���n����3� 3�
D�o�}	�0p]@]o}c�1$��Έ	�򠁜gҕ�
���X�j�s�5�H��e�s�Y����`���r1:���m���:��������'p0Oa�ߕw+ ��_���C�#_amZ�6������쵹I��~��اiȶ�
 �\�*o��g�[w�Z�9�,���_XII�B��l�T$���JnLZ��rꡣ8R�d��:�[� ��a���Pf� ձ��_4�$�<`֬:�aC[,cqp?g��p�Ij��}�SC0��Q_����z�� �������>���N�n�/���?���%��W��/��|!VT!VH���½p�s�F W6�����x�/ڋ�����
_��Tg~��,�w�Mx$���3��<��Q�k������8i?$Kʱt^�`�;cM���1� ��P�bS����W�)`�l����1T� W�f]T�1���@�m��x�g�5����U�(T�g z(�/z����X�Z��B=e=ق�D�z����S/�2n�j3��YM �yβn�ڹ�C��t�(z��	ڝ_�mcX~��Ƽ��-�@ka������&���ԇbG�������6��X%i}G�q��D6+I�s��H|�z��H�ʃ
?�_
��	�1� �^�v'wn6Ⱥ�ȯ�����
�� ڳb�AI�Nz�/������?Agx���40�UI�d�z���Q�XzȨL��X�:����=�Ҩ� pe�t���� �{���`����<��4��:�[7�)�����9�XhcWYQ8L�l ~�K�������$u����6���A�o>�K�� j��7(X�*�7�cUy�pz$ik�~��h�U_��T����~B����{D2 ��+ޛj��= �lNwmv�J���9��Qu�Q��e�	�eDjw����w�-�;6�+�Yk�u�0"<�I�D>`����rF~M���C)u��,���]u���<��[
����R2�L�U_��j�i�~gbp�e|��Y�]�֝`6|K6��/��A�TT��y��,n��
���|� P�.)α����/��Oy��l��`#�`#cP��׏�5t#�`τ^��p�_4m���[^f�Μ�i�i{�wC�>����&&�u�gI��?�J#���nݸmn�%T�@��s������H����Ot{w���<�OO �������&H!�=�˸}e��g.f�æ{4�����>��(�B�D}�����[��9�P7d�X y���/���
+��~냖� ��I����A�e����]̝����0���s�[�3u��У�B_n�]_d����R�l��,D��A�1zQ�9�\\7��cqN�<�O�ap�o�����_�ǻ���g*.�,Ԉ;Ŋ�| �𾈑�^�P��)]��g������Z��6su2.����i���DocK
�(��}��.�� �����@���^+e�o{G^��WaVfC�e^��i
-L!Hhv2lp��r�@>+��(2�I����!����-�!ӡ�I˩��L�Za������h��\�}�sW),֪A��Ș��-<�bR���U�)v�G�hw=s�]��Wt�T������A�~��Tť5���%�Hk��-�<���D��p�
2#�C�l@�5�J}v�z\�@�íY���kP>�����W�����}�v��3z������	0�"�<�"���i&R���ޔ��[&5RAeZ����;�9u	7��9�GF�[�P>+>A�-��sR�5"�_���PuO®Wo[�+]��;e��J�%!ƭ����ҵ�4�����"_���H	�������*�OL����^��&��x�<o�1u�/��}6��9����Ow��52�?���[��jc\<g�c��T )VG�J�B��~i+�ֻ3��{z��3�,��� �(u�Y�-�����F�wN�K�l�Q�m���H��ڂ���
���`���B�+O�Z�y��M��5�(c�D&���5S�t��CX�ӵz�þ�L���\���Y�26�S+M���uܰn�m�'��Xt{�����7��V6���:�Ţ���neo�����,��/j���ک}���>c[�ݴ�}�mE7v��'V��E��߹��*]8s�yI���]8����LsFS`zN� ��mWĐ��4|u�u�J�;�����-r�I�����CF<Y�qqN:���`��Q&~�)��-�k��h؄���I���yv��aL��T#�wh��ja������fY��C�>�)�XL�u���{A���:SA��ݖ��敜�=�;o{¯d�ߒs�]�kF~>������Mm��L'�3����,�:^�ZvU�5���-����PE
F9�-��|H���i�]���.��A�$�*�ete_EEt[<D�Yi
#]��}�	���T��}|LS�V3�ON�O�e9)˂���3��=hv';G�}J�imΝ\�<8J��]�~7��Ott��ʉ`W���I���g��Ԛ3v���ݳ��=F����AyH�ͺJ���_�tPqw���[��x%FȌ��aWG����:��?|{���ǉKrI0�����?��Xfv��
ל�K����v��<&�9�c2�0��M�17��	q�5o��$ i����x(���V�X��TS�1�퀟-��y�鋖��^��PI4C_�]���S�����Y���I�ia�gn�5%R��{�Xf~>�	�g74�~LMy��ven����V��� S%_4���)O�j�r
�Wv3�H��c-�����Z~D�{x������N"�6��OM�`��l��I�e��">���I|�՜�}_�y����s�f�nc-iTQ�w�T��U@�2l7m~��U�SA��5l��=��7x̬���Ύ�	c��G_Alș����A,{������Э:���|�Q�K׹C�]	���X ������ph�J�= ����Y�'�7��`�A���L�>Sģaj�����d*()y��Y�X�ucn��|�־��9���K|���N��.���{��4!lm�')��K�r��4�.�j�oi�!/����}G��Z��IG�q�_�x�M�*�/�#@��R��M��ח8��_(_f鎛���#Տ��4ݰӁ�@�*<-�+9z&�N�D0�0[=���ЁCY��s�oMenb݀䜓.����Ǻ%Q�ĥM��$���H�:J@(a-��D�ʺ�� ����ݢp�z��dVs�bhO�{���x��r;����z��}n��Y��ݕ���霫��b:��k����&���8og�������~���z6d�?,!��t�� 5�*���*��X�=$�a��c��O?����)��W� Nz��|���[*�kf��ao]wAڟ����hW�w��4G��ץ����������Mi��x�4t��Ȫ��a�Ks)�����ebG'�:U�_�ퟗ�*_���n?��u1��Y����[s��=��d��e��GG
�뺃2ޒ>�l�M/WE�����q ��uͷbt�<񝉉2�^w�V٩��I�E����'��S��� �M�x���_v=<�EK�����_�O��P���_#�|�=}k���]C�7���ux�S��g����S�M�x8x>ms�%4��F���k*��Y4�}��H�AP�v��O��v��~F0�(��3�{e��7��m��f��wW��'ؑ�`�!Jn�gzI���2� �Ybcz��W�|A�х�4��=�����
cH�.�?X�n���!��ۻ���Y�tٺxж38W�C�R�uKhI����x��uKe����o+�z&�3��� �+HďI]��D^�PR��[�� oP���٦^�0I���<-�]��������-8�3�`��� g2��Ot���/�#�(����x�Ľ_F\�wFʳ\����Nl�1N�s%������V�"�r�n=V�{���{�Xw0��X��T�b*������|��EN�_�A�D�?녰|]Qz*>����'?���]�:G@����7y��6C�����a=4Cv��Tj�?k��y41�?;܋���m��<�ޱ��}zc�Q+g���{�Y������|�����B����W���a��@�Y#�_¢����0�r�dAh��i�����C��Hr$�~��DHJ��S����	qA�	�Y�8Wc��Q�,|��y٠Ox�7	�����:vnB��s73J��7��pZ2JM
ċ����3��*��NH�2?ϵwZ�³묓��!XE�7c��1���\{X��,�'QC���8&ޮk�;�z4 x.3fw�&vK��4����86�0�Yҥ�)�0�	������_��ڋa��ǟx�1&��G��	�\��0k���#nq������׵�ʵ�գS4��˗���g�'[7k��8�XF�B�7��G������i/�P�ƪ7zE�j�X�7�_ �d�[=�����&��J�^P�(k6'������ņv+A�OH�Z��C����i��<"g��R��v�SO�WRQ���&6�.t֞��I<5�O�X3<��h�-���Pǉ��4���;K�Ӻ��U�����cSk~e9�����H���AI�B�E��]$�VU��[���������Uż����y1�)=�m�����ݳm�j<��<5�2M�?<�� ���7�ߢFrϓ[����(�'�җ�q�ߦ �A�뺆jQ(pΈު*{8q;��H�^��$�:�q>���8v�sJL���
ZxW��?�[��H��@��f?���NB�T��+ƛdP�
 �d@�����{G��P�)؞�f�z�u��?_k��t��o��6x��P �v��,��ފԇC=�����)��RB�r��P��G�.��Kś吞��{è
��ph�v�f�O�\����@�*�g��c���`�4 ���]+�3pi\�#TW�[�w&_�� �5��H��؇x�=�H��;DiM%Ep��l�b��4�3u���w؍�j�سН~�]/:��:�t�ǒ&u�>Φ�NR��T���c{�\�?��	f>�D������jΚ����CB*��D��M����|Q|���.�'��'��ӤQ�m�)q�����G��l��'�UJΗ՜4�tu�h(^b{�����|�J�@��B�j����ZW�oZ �<J��O�z�<#����;����;
b�CI4�F@��t/O`��ˣ<]�Pah��r%�t�qA��Drz_0LP7.����u�ۺ����ӣl�@{ʚHmw�6m�����yS\��:��:3��v��b���}i�dѯ8��)7T�3�v�!y:j��"voZ�l>��^3�?�W��c�J�^$�D\[�{�ך��t���Ї��d��8m�ݳ�J�mn��1���%�����w|]y:EN��Hn�p�W�������4'��?rO��vCW��ݕ��E�8T���g����T�3����y5�?7�94��iݘ���L��*׮��x9x�ux��S�9��R��F��(����CD}
��2J(��*��,��Qq9�,���&�a��G�|*%N�+�P��s��;��EŗD��L�IW������"��o`�u��U��!p<�zn[
 ��
�~�I1�\*�?�f	��H�f-�`��ܞ\��i��T<>w����c~��hK�q(�Q�BS��_���5`��z�,��~�]`��%c�,M>��:lb�y�X!����V��@��r;�V3)� ��&����?�����ުM��� �5pRԡ �X|��B%�e6�]�d^�'9=�R7_ޜ��ѫ��y,�OY�\4]s*���] ���ksR:�k��e�b[v=7��)K�$)(؎,�;ׂ��+JA�P|wZcg/4b����T:?z��O;ֳ#̊N��S7{t�zrm��Ә1q��tu,a#��VPܑz���C>�zn��@���} Y��˛��f��R�J2�yֵzXc���7�
�c("�A��p������ƽ��<<4�LXq~5��j-� �g�)5�m��8���L��k�C��x5�K
�'�C� T�v�=c�^>�����=��`}=7�%�a-�#,��bR�epJ�%�^�-_K�����
'#�v�������_�Òk4Yб�t�ܒSCJ$!��u�mAA�������(��r/��k=EA,dWg+��Ȱ��8�wv��s��-�#�a��ypw��O�>}�74��$���5���j�!�Ҕ 7�'�����Z���w���l��t���������U�qQ97� O���(n���𶒢WP��{��"膔��9���8��5��y}~5�W�ihB%�����G4��@u�j�0���z�r_�lѫ+��ܗ"�����m�8�����<;^���E!~�f/���^�z5�:a�IA�����-\\�IH�X�{h�_���z�h����[a�PU!�|/�3[�̝��oN��27��c��qx}}����2�B�7%�ޞ؀�$�t,C����]��q��n�5Յ6�,��������F�2��ſ�^͢�`%�_�B�����),���L�S�~]N����(p�t�^l ��k�B�R]�9�Q�ڇ�kk�_����q��ރ���駰�D�ŏ�ɜ���C5����o@0�$����z�X�4����cn!��R�lrjj�R��E=�Sq�$g��\��5\�Ƴ���7$�~1I~'\k{#A�kA�?�z�9S���#{{��4��p�vYq�A�w�1dQ��oN~�����a���\�>K���+)�����F;�>ˏ�joX��A�T>F����ܙn����2sTP��)¥�7��x�Gd��'){{�qb5���DD+��s�g3ܩ�\�j4�����~�삷���VZV步����_��]�����Є�C�3�J:�ZXוb/�'�B�i��t�ae�]w��l,�? �԰��J���4�Hl����[?�%.P�uy��G����9�s����y��*�a��:��){{�I��{RF,]ȷ/`�Fս �oC7�B�{�X]�sR���m��nt���Q(.QI�*+��g�]�nW��_�kء����50�����B\����7@�:���U'��1/��Ć4U�p'	`'{��f�,
pw}�p"T��[W�Ռ�_��
e�u��dv��\�.,�q�R\��u�j
'��!�:�R�4Z�ȁd��xp�I���p�s��咏�[���^��C�+����Ce�U��/E5��۟�B%�q���i�_*Ƌ�`�2�������#�T��Ri8"g=�ק{��FjO]k���J�{�-�o
�YY�)Ӻ�M���!���uh	�Yw�w�R�
�%ǋ���z��0���$B�V�{��������P�I��
������3C#��(J4�L �~��E��S\l'��t5E���݃a���p��h.Lu����M����P�7�^uDI��؟�Ǩ�� ]��l�6��.,l*���<�R[��*Q��FC�����=�"��m�;�.�#x ���P� s�۫�~U/��d�sZ�@�9b������Ъ\Be!�/�E�j��@F�Y
bG�G U���6�Oſ�Z�z#�я�La��S���e5���Ԓ��!?x��g���-�1��9�dhC��9�G(˥[6WS�<<�PO�ԲC�P�_�Ws<�G���/������D$B	Ov
YK�Ȟ��eߗ�����IO��I�o)����!4c�:�|�{���������>���y�׹���w��[����������;A��$h�B4����tsB�߲�̧�gZ]�h��������<��d)���Mh����;� ��k�>�����L����oϛ�m@�Ʈ��À5 F ���Է���S�4oR��D�����s�����&3?_�~�<i�Zd�d����&�%�E�b�n���2iD޷x��. ���k��q���۷N��%��ѭ��ss̓�z��Ɓ��<��,�v����o�k��5�ZPj+�IZ�r%�����ٿ���n(<r���G0���B$����x�ld���4�r��%�����������Y-����m��M@#�m}}�g��G��bmu���Z(({������k0_�HCn���C�g�5�&�>qk�S�����vv�2��\wr����ٜ�2��uX^��]����U�����x�����j���	h	��__��?;�I2ˈ�ό虔h���A/�n�ĭ�'�mssA��,B��G����x�m��E� 3x'w��D�5��וLb���`��c�D��� �;
��p�ϟĽ�k�]s͗#@����{�qS�G>�~f�σ�"�3a��io؁R4n�3q�x��N ���O�{������iw��s���t�͟S�t������rD��ȱ錄�����Ԍ,�W?��Z2� 朏8>1��۬���r�_��>V�k�3d*�k�'��߶m�)7�e���%���#�Ǻ>Ǟ�y����I���'��tR���	ٔ��R3����B3v�Ԝ $Q�	NNW�У���[�-/-5S��U�6��)s������תƺ6h�Q"hɺ	�6����Fo�\����	�5�:Oh�04R��8⬉3)߷>�D��\��c��)0���W�-�>8�zY{���Ұ|=ߺ�����_��V�=�����Z��UHA2�q̀���(��3�v�'o���6�=�R�V�d����Fp�eGh�F0b����%j~ V�B9��{^�@�*��"�vj��K�G}V��Au�(m��G5.��}���/��!#��.Tj�P�EeJ
�KG�<ƯDd�G�]Cb\7 ֕�,JHX�K`����9ڈ|C{����ÐO�;Mc�'Ҷ����\��i+ȣ���q�Abx>-b�Ǘ�d�70#C�`��	Bs[�O�yxd$0�41����F�/�4���n-��]A�	��X�WD�,�� {<�9�FH��.��-d�<��H�i| �s܁&tS^�&���H��cQ�	�?(�	��RoT�</W�XJc�"���M�H��&��Pu�;����WA5��	��oej3P�E&�^��0{�[�U�N�K�'a��nGD� �% <I���?��_b��p2jl��^/��K����sZڑ;��I@_o����x1�h�ޞ��FO0Ϫ��--�o'�
�����'�+D�pqb�Т�..
4�
��MH�T0�V�^�K��?KK��*���lM��,�%�`b%�=���ڍZ5(7���m�О9��P�ƍv�#f!������g���N���%���l���p���FM��0��>� ����o�t`�y�߫{�>��*{��m��@��� `�U"�{D����-<��n���3�Zg�h��8��f��J7p���<�n��Jɛ7���-�@����_�M��-P���px�����#	�@�d��11-��G@��|��Ex5���@+Aˡ{i�0����(�8F̗����˜kk����2ww�\��	5Dہ���������%�f�`�� �jڠ��ۢ��F_tzz�2�a�:�C-Ƌ��O�>]�f7��?Uu�_.4��d��E�Z�SPY`�N�^��I��Y��
�����Wϭ�[]�Ե��!�D�S~��e��֕��&/��T�P7�U���t7�+�ra���P��4�5�8O�u��hnֽ&��\p��>��76���y3[��||����n9SN�����✮� �������s"���X
PZ�e�0�o >�3�^UWU���%ޑ��\V�)�6�t�UNx��QPd)=c����~��k#���}��p���o��_��<x7$+�$�m߇��x��Xҡ��ru�f���H�oB����˪�+A�=�ba������P��	�$���9W-> ?��2=�`4���>5�HEZ�������W�LY�+��j~�RX}z�b�X�F	��0-��L�d�HIPQ	:/�&w39�\���q��wL�@�hyʌ@Ӭ�V�I)u�ַ��(� �����U2��fܖ.yg[�7�8�̸Z�r`I��xUU^To�铓z6	��##��3wuL���a7���Р(4�G��Z3�J���b>����c�nqC�P/�Ƅ"3��*�b(��6X���D��ꅃ��JΊ��d^�e�U[�6�L�l$c�L�w��b���i�T���������xU����C�UU��Y8�%�[�x9+骫�+g������H
����x��*e2�`c] 7a��gh�n?'��]�>��ы �A]1r��s�#������ã�%c�e���L�]�\�k��	�A\_W�-� 9��`e�{6�,���ήO-;5$Ԝ�b��j���:}��3�?�6pE*��c�%hȤq��t@d�"}[��8���=�6�w���a%�s�������{^y�ME��G$IV�63���X�����]�Lrs��IB�≸���g�4�]�W9969`0/Y};؋���\i�%�QA
�����p�dL�ߧܼ�,���Y�Ò~��x^E}����������DW
#EO'�����<-���>1����w�I�j36X3Q)C�rӁ<]����1�}�v.U�L���J���DO��oo���
��(�W��"$f�	Wu�z�uH�1 /3�r��� �@[Q�l?�����I/�[ f�c�>�d�Z�����mb h-}�g�P��`�&�H��EZil�\�A$�hvY�3�<�t�b�}����A;�Ryv���ev�ç�����C���.�F�T�)�9%�=���N\��8��W��:C��Dw��tv����_��(�]v�V�
5.�p�+���r9V;�����:�} �OI���W!ݝ{o��f�����5���B�8��@�ي���遣|Y���J���qA,6�6j��틛��OA�$��j_p|$Ş�,���F����r����j�X�|��K|�S�,�6����w�M�����R��>�� ��w5��*!�!N���M=���l��|p����+���􆧾�E��,Y�@�����YBi]�3QI����~9�G2g�`�4ꕠt�@�KDu��\��������h��$2U\@��c���CH0��E��3�#"r�@j<�!3_Y��q{&��]��"�g���"�б�a�\���$)�	��e'����I��J��~{==ZU`N5+4t�K���_�� 9�Ԟd�~����	��"u]Z��& ���ڔ�j���I�$�1����EP�m��c�Յ�:��-; R�V��K^��t*gln��}��>�Xv�x�����_�b�AV���������N������u��fK��>��ur�EA���&葠(�q���ҋqzVm'��!i�i5A+��;8�N�W�g��ۯA!7���sx�O�>Z�:��Hۡy���q�_���u��{Ig ןIT�}H��qA�?b<E��P����U�~&������gh��9����2O�xA`t�i��=�t.�An2Uu�5�t���:�R==��} r���P��"�b����H'N��Z��4BF��̋]��K��C�f"(B(���%5�ײ����2l~�~�u�L����ϻ����-��B5�m@����������J��ttQ�8v�!aq��
��Р����s�)���t�v|�/�Iz�%�!��.a�W�gJ��:�t ����N�T�J�(XY�83��I�wM�[3���9<�xI��\�)�x@jv$�����=C�k!-ш]�6;�?�(�oh���\O��Q�ǎ��lsS��?��A%�Y�z�
 hј�Ls�)$!� ��M����mon��1^6��,�Bv�|����/���q�(������ɿ��+�I}Bx��۬uH .�D?,��#4Ck 6Ed��x�G�:/��$=&���cQ���jS�R��j��]�b� �.]���(@�뢥.]�[{�6S8&��˽n�p�#�h���R2org'�����G}�m��6Ӗ���*\����?3S�<�� �91����܅��j	��E"	���ym�����=bm��+����V�L�}�*����R

rmU<��\|p�Z����"ĺ��'�1�`�*Xҡ4��i���VQ,}-���fހE�c�c����iy@�L�oԈ���̂�D	�d�Ds����P�}!x#�+�?pn���~�\��ut/�h�ǾM��/"�� ���5�e�v��t!G�@���^B�+����.�@\a�����>�MԐ�qCC���OU&�3Yh1Ȍ�?1�sمf�p<�_�x���D��!Ŭ+q i��]�m�'W�鍘!�?�Ek6�MAT���~�8���~��A��ö��np(Aզ�?778VE��7����f�DCf�ۘ�i�2_�%c0q�R�Ǳ-�lN�<A�8A�0󢢢��� u�'���u�s�<Y��B⨈ӄ)�I[ZM�����>�숑K�d�=�,�;4_��F ?���L�9����[���=TG�6e+�@����WS�It6�����Az�\:�^��Q��Y�ʀ��>i;:Un���:r�у*+!�S����(�|HE����
�+�������������H/��pq���ez����(� fm.�������~U�̌��e��A�6c����$�}�{����r5��}���ˊ���t�>%W�����@p+7��Ƭp�밑Y�^��$�=Ӂ�)��� �3��{����v�b��FD�SdD���;/
y���<
7�����~H��T�B������T����{kOD t�~p�A����Ac;t�쟓{�뚗��I�Vk��E�*�"+�g{y��1uS%��Ǆ� �@�= ��Vh�>�����!��|�q�f�1i7,�t�.gi1�����3j�x����;�O�;=�{kޞe	���*y��M_}��(^���.�*7*�F���a�3H��q�(7P�5rD�/�n뾊Q�����ҭ���,]e��#8�ə����R�{F���V̯��׍@�!Z�_v�2p�=��0�+bϵ���P�V�P���S$���'а�Z�pe�g|�Mm>_�Y�!jHN��`2Y�/E��~�SRO^���>��
לMm�Z�I|a�-j������n�2��݃�Au/�؇	��j� v�Ji����QM�G���q�����F�T'TF�����w����}��xDO~ϫ?Ad|���jD]@�l���ܯ��,i�F�`�a(�-�F����G�gi�uKs�� g<s:�χz���M�T ʆBc����ڙV������2+��X�:������2�`���4���B̤�5������}[�=��M��$���4�(�(��Ie�D�HȆ`�nƹ��[6��b���Y�t䚂O}�?AAr�C9}���<r�N{�^�KT��4�d��u�&�Q+�'�n�+mq���TF>��N2l׬b$9��E�1�~W�l�ڭ%���^M~�:��	U�P�������@|�^�z�*��&���tv83M�+u֯�~F8��k
j�g��RV/���xس����ՖP���)M�g����_&u��u6}֢�@c��0P�c��d!1��>7K�<cJ�*��?=6�Ԃ�M��w�D1t~����".+{;1�@G"> Vn��&4���%�(�!�!�i��=�	{�a�6�y���p�J�肐��>��q���f�����X�+z�Lm�+��(�,���v��5��x('!���quT�8����r���?-�&�����#��&�GԞ\�-qJ�<h�9E}� |T�S��è3|����]¸�t	����h�~�j"�-v^I��F�¬CX=z,��^a��-ѣ��eNG�&��p�n�()�iԈ��#�Ñ>Y����3	��ۛ���IK�嗇2�!����'nfiΩ셌T�%�'�P��.>mo^c��ߎ,�����o����Ȭ������ ��};�[莪*ī]{�rI�u� �����}i��XH^$�*y���g����G��7ծ��j"ʞ�s;��zy��s�Trl�7MF��2�>*
�m�b%�u�T"���U�U��G�����3�� ��?f�]��*g��X+�,�*%���}^)���j�H�鞮�,�|6A��:fF�������|�KR߈cY�xDV\�?�P�A%�k�t$3c��2�އ:{�g;^�����⵷;-K9EC"�P��Q��-%��m
'<d�|G3'� -S�U���ڝ��Po�C���04f�'4�\��s���h�Q����Pm�a��`9�?.*���XW�N/�|(I�hKϵ()�B��Ó$�nT_��S^������Ae�����f���d^t�[��옝��ᜡA� v̬��������j�CL|'>%�ToiBz3U䏴����~�B�9'��ʝXy�p�B͎�O���}jQ��[�vLIQ�T�<�qz`��bZe1�h##�ݾT�L;��p5wrr�M�Ǜ��������$+'%ER_Ŧ>�՝-*������Jݵ+M�"dz!/�52��vWf���C{�C
�n��=�G~]�~��>�`W�T)HkU���o�5�wX�7��;�o!�#������u2����P����k��bRH'��f ��q�x��.���/�B�ն��WK�AnAi��/]�2�w��|�77G��
��'(�|�z�G��ج�k��76�s�{���l)��ɬ���hA�J��Nn#H�\�k����F�O\7��8d�L0s��$�*��� ��\f��^��?v¦2[-��(~�Og�)�tO������X�\�~�"�dD��&8����
P? ���b|�� ��=I֝V��y�l�v�3�鶷ہxq�BII_hp��JM�n��b%A����� ��I�x�	���2�K0�\�	�QTW�H�����\KUU�"V7n'mϭ�=7M���J�κ��e�QudTF��-�	%W��9�*(��֧�O���&1��f_	d��/���d��"��W���,;8��Û	�C�a	M�b3b�+8�$2�9��0�^��-W�
�	�s��t�́�\��#�^��Z
.�.Nc�An�A�L�g���,�n?�!�3�4��H���������Q�ǝ�D9�uKjk�]�M����+f0R���i�#��
H�SQ�~�uA��ghe�t
�3�j�s��g��Ig�l��S�:/T�tu��^sy#	5
3y�x�
q�ix3�ٌ�\IKgܹ�,��ʀ/(5n*���=����jo+���.
>S)l�`�)�WD��W����͜Ø�:C�W�#�M�W����rF�M�=}�ࡔ���-����[�Rf'�d%�$����M�F~[e
v���,~��#�y@NoU&7�J
�?Օ�>�9��䝮p;�y�k�I" R�ab��:E#C��}���q��
���!����ʻ�;��V��<h?ݍL���t8��:Dam jO�?��eekv�Q��å��yͲQ�}'�pJ�p����lX}������j쾿ˈ>:�h���"P�?t=Aj��p�[�]+3�k'�iWa��3<'��^̓?w�	����2 z4�K� 	#��sm��s�s�Z���nV=:�?L6�ܹK�3�l��'(����m�G^�$����C9NLЂ�]�yx����|��+�Ꙥ����{�٤O�:ҧ����U˻0�qf@n�$��OC���)�8(�O\`	��݂oF�V FI����P�㱁I����cGlA튔 (�b�E�p�8���Lyc��P�i[
yk_��$�@�ޤX�:����� �`�Z���J���.���:f&��?_��8�����W��g��b<=���Y�a_�djR�{㷪I4��abYC^�����;9�$£\�q*yok�6�r����_���ҷg]��5.���C���߃U�-�>�-m@��8�$:%��ep�!�*>3<�k_5�VB���C�J��|f��{⹫7$�v.�ٙ ���>��_~��#q���=H������,R����Y+��0�:c%%�kR���"��q&����R��V�ww]�5�K��,KD�LH�[切�e�{��&��`�ݣ5�G��|X
'P����Ư�{���@��Hd���C�R��l�HE��(�F����^��cs3��]�������E�]
Ww*�eS��r^�T������X��~��F(����>7�!���w�����Ak��O{���	����:jc9ˌ2��o��ǡU��O�9�c󺐡�k�	]���'�^^�3c��L}sL?����}v����ڙ�w��ׁ����B��<�����Vh�(�t#�	h�9�.���i���,mjT����������������e�0�����s�`^�6�u��k��.P&Z挄o(]��Xբ��h�:A��v#��v��k�h8�h��7a\y�g$!��Z~��6,R��3_N��;f;�XyGH%�
<����/��ݴ�)C�v��J3aJ�Lh�&�2�k}1SpvD�|>DJ߉X��P|���R��D��V�F���%��	ʨ�A�Y��{H::Yr��L�=��[/9�iv�ۛ0������yr���ӏd� ���K�
8: �(�.�D���z�#�J��@膦�v��}v�=9�����9�"-P�E%������<��V�$�;��ߍ -y@�.�d���XHXH������ѥ/cv����_�h_F,�B(I���Î�Z�I��,~�u�#'p�kХ�����$&�,G���cT��GB�3Kmnp�z:���<7���_]��&��'T(^M�/��k����#����u*�9�PE�����GI�F��`gCCA�ngZ� ���S?j�|��Q�K�.�Qv���g���[�g��Fu5_c걫�t""b�\Ei�:�t�킵�g9����ܐ�[t�8��}��U�>���RR�w�JO��9�x��.�EV��l�xR��m0�a��9ӵ��.z�N)@�w�cJ3���eR��<+l�:�Y�z�2�]�l)Л?�u8>��.#��g���zU3��>�MQ3r�nRi� I��W&�RgHڴf�J�� Z�������OW��Y�H
�����^���?U�	rz�U�Mq4�^M ���l>A����֛ޙv�����O��X-*���kY���Ŗ&uz��6�yA{�)wj�O3�k�!�ÍTң�>��� ����X��םi˰њ��K��Y'zJ��%� ~����o�ƛs�������r�~��t������ � �Ł���/(T\TB ��iuY�۳�����$1΁�_�F���B���L���JU�����	pHx�ZM�޽Xn�<���^��m��4�7i�/k°�� IR�1f�Y��0�?AE���������~���7fU��ɳ�-W9��7=�Q6���8	F�;��xڤ_L���&��`J��������ԓ�F_��Mv���F�S[�U��bi�T�E��0��h�A�aYQOd���@(���H+���Gg��2��5��uYY��,��˃ڒ�dj戴���b��\^�ܽN�����+?��Qk��F&ޓ�\�ذ}��"��an����(�:�O���������/xZC@"�t'V7�NqEE<-�E��O�hu^���ִ��%�z����:�]���󾑹ц�s�r�d��q7�w�DYAO��Y*~��͑l����D6D��5�՟q��M��y�p'�?�2$g�-.贅�(��=��Ͼ�z�	ݹn% 
D�g��]�����T��`�yR��R:��n�m}�_��@��!�B��Y�d��O�����L }�U%��i�)<�a�e��P��l�IՆ~��ڪH�cý�ӳ��js���H���uW���J�s�fSih�����d�'�'V�6�O:=�sѴ��Vn�gOH���S.]Q���ŵc"��\E2�!���P�D
1>T��J�	�7\QQ�tGyz�h�ط�x���IHx����D��<�8�Y;.���m��jY���o�[���Th�NF"��cSg��5� usS�ڛ:&th�cLG����$�-$ޅ��n)fҾ�1�}W�nx���u��oa3�����&Jؼ����qz���q���q��3kNNN�T���pu�ίB�>�'�$��t�zh�G���R�:�X� ����Zm�ԝI�ߢ��t�9�87����m-��CC�=Q��' �W�<c�8v�wC�-����C��]i=�!+{�E���G��PgC"���Y9k����ኃ����[1��Wĺw�����5`���Au+�����@o��UU�ɛ�roS]gZ3��(�p%:'^(yCG2;A�kT�W]���1���v��g"�ZZ��M��4G���u���O����gĭ��Bѥ�{�p����|T닢�4�'����i6�a:El�N6Vإ�~4�/b�\��}*(��朚��r�'���^�}T:;m���u�Y'�dF���Շ�A�K�k�%1zz���:����B�H�6	j�.u�8�g�/B6���<�_�	Ci�]�	yVp5y	1��$_V6Ԫ����.#-�{�r����p����b��*�7޳�)f��[������.Ǫ�t ����vA�Y=0y/OZ��YR�/q�M�u��;�ݧ�ٴ�#=c� �
(�Z�d*w���"�6}��Ɔ8���y�V���B�f]��S�jlj7J��!�c��kލ�b-B1=��(��@�t��p���n�R�´�9)Պ�����K�V������!���̀5ǰ�m�i�g7D\"���L���{��B�-����[^�����ٕ%B.�xS	�fݚg�;/K��K��6��&ZZ��A�2����&I��c�6ixkP��z��MW��2<D�E����r?���e2gj���� sQ��`J?��	�������==��G�a�'�d�1
����g�	���XHz���,�6��!LK��{��=&��3�{g~]��n���ր��޹��_��"w���hWE\��V����o�:�Zh������l8|��@
�J��P�	$�S����p�TTe.�.s�34;�Q}����-%"�����K���XB���fF���V�a5���r�lN}]4�R��5��gE�!�'�%C/͌:&g��_��x�{B�DE��5<eWh�$�-�6%��u'��V�E˝�i�ˎ_���W�j�3]K0s����D-o{��'�bz�>�N�@j\��ZB&J'��D���g�G�~���FY8j�<�)ФT�`+j�R��"ٝ9�����Ǧ=��[I6{3��;������I�l���Xj9ȝ s���ތf4�T>���?���c��I��^x�|��q:�
���� (	�W&l@3������h�,���mE��Le��K<�!?wN JL�@����t�Zg+���'p �*4c�<��-c>��O��"�[<�9��%`��h��Vn4�0Q=A�Y2����$�-_W:X���յ�{\4K���/֨.�M9$�g�G�gK�a��I���<4j{�m���a&�l�����C���p���~]q����|;i��ى&ݹ�\�i��M#�x�����~t*~<aI�B�s��5K��A���o<�%LL��%�����W�4�wD����E5��)Y�i�j��������vHl�>f��=��b\G�<�Q�e`�Emy�r{{��@妫W��G�G���"�@G�:��h�Y�"�&F�Cw�fI˥�վ��c�؃�
�;���Ƥ��M�����u�%�nyU�YA'X¦_R=�Q�E˩[5��g�b��5[�[�F?�h���=�X6�y7SR�;���I"�M����7�Ӎ����M'�xjgO,r.��s_�[cS�z݊�c�������E>V_��X����`Ե"w��c@=�loV���Pxv�خ�Ţ��-�n���	���^V���/�䓿ہ}�󳵍XD��T��ms��2�n���
���✖�If��uta��^f����`��?�^xTq����y2ZT�ΰ@��qѕ^����/�E��]�g�,�3�Y�vCٮ�Y���t�=�y�Y�qt�Iٯ�g'��&��9o����l��_T��)V�RhJ��4���n���H�L-�G)27s�ǳ:I��Y��I5?�YR�X�F��\v���;�S�m���k˽�����;9�C���7i�]���8歕)�w
	����]u�V5z��`���	BB��}j��Rô��+f�~@j���a�0�!�N�g�4Zv̤
�B1]���$,���f�����e����ە��XD@��]?�e����綪H���3x���q�/�.��)_m����͎-��yx���,�(��1s�Ǎ:+�C���K�O�Z�W$�F�*/�y�.�b�)Ø�2��f����Sa:����F?���q�G~��D��9>�t�M4�v���{���#r�	�U똩�c�ʫht�g�u1�x/����es�h4��L�?T�{tnt���v��W�%Q,��vo�N/Ifv���{f��;L��fVE���G�/��#�.����"�[b��'Zj��?R�\��_�c���U�* yKmj�|^h���L���U��I�&P��̊�}�7z!)i����Ì(���s�Z�z���7��uUڽ�o�3+ҿ�&�o��j�|×��b����V�u��#�������&D��nX���(����_�����v��jm/����LN�n�m[p�bnqzǏca�! ޅ鑹��%���������h�5��E�������$�Zw�Cَ�/�uh�qU����w�2�p�Xտ�����k�Ӳ>���3ή�t��IО����W�wwcS�,ރa`��dㅫ�j8������[˅�鞆0�R2r���Jע�x� ���x���s�+|�����a
�M��/�.z�ݢr�G�
:ť_Z��jǡ�eǼD���%k�WR�XL��f���)��e?��v�aXN�mM����-4'gM�L.���f���m�4"x�z������
�g<���vy.��E&v���{�X�o�"�
���0�SJ�]f�:3�8�[��%�6k&�9�Qa�|��kc�VK%�� M�_�0�y-7��CW�Y��)�M��w�����#*X)1���x(t�dЈlʉ�~��]���)y���Һ�3���wʷA���v��=g��[A���abڌL�F-k:��-~�Vqyy�9V05�Z>�:l�oG��Ȯ�f��h�O��=�n��S��R\���?e�;n�&>K���v��(�`IE���_���i�=��'*j��9��d�p�
��Y��.�ԯ��+�Soe�)�S����.A�>�:�p�Z�����5웳�ޡ"���έ�'-��蕷�rI U�O�{�*�������e�������+����\�v5Z[Ӟ=�My+�E�se����4ߵ$�?eEభ�1��
KI6��;C�睎��YF�=ȜBjZ�� ���~��
 �Ȫ��#̱�/�E��r8k��`G$Ѵ^(���:���TI0���F$�pa��b��]&GDd�$�x�����<�OMnw���{�^���z�sjΟ58y39�>�!22s����W`�+��b)��v?����X�a������e�������|�zVs��A���!�s�o��v\L�g�	������2 �,ƃ�l���š�����;��	����t���۞c��7Y� 'v��ΕK�R�7Qҷ�w��Z�I�<O�mɰT�M={WW��Ee��a�[�K_��b�>��y��DAH�<e��y�:�&=#��K�2��OJ��s>M�ϙ�.�x���9��P���s�#�; q�1,����KP���㷦إ�,�Ym� ��+ ����M`*6}N����԰{N�[2��;¹jtQ�f�-����}�B�[2F��V�h���2At���gl��;׍~m�Yu�+�2�	���K!W`H�[_6��EVk�Yb!���D������g��;�[��.����q9�n���(�H����B��A^�����I��=l/�D��^��h�cQM(�_ZcbQ�;���CٌOm׻�5N�'J�lm#��]�B��f	������4�`"@�#��o��8j����}�x������Y�W����,y���|�66��J{h��Y$���$�����5�� i���G�e�J�}�l�uk�4W̻�~����O�.�	�n��Aײ���F5[�z~�wo���+"8,t��e�7�_��)������}4�1�ކ�F�A<pP�,.?G�ï��?�8$z0��,u|{�|¾m�OR�^�pFb��(�G���<LM�.������L@� ��?^|d]����n�Կ�����J��1�(��B�o���QN��f����e��T���h�ҳ��E�]�0FP��Da��i	V-J��u�»�k��P�ɛcyN�Yx<Sb2�K@Y�M:�w�n�"!sse?z���l��L�0#�'��n`�� ��G�&����<�������߶&���4�h�<�̊�m��20T95��i��?OH�	�'������}C� ��h�'�s-(��p9(��gM�_@��30N2��͗F?�65GȮ�,��r��3Nb�(�V��7Zs���*�Q�U�F���ICޛs�����c*E�d�$iD�f�A��߭k��N`Ys�X��
�r(`�H)�F��Z�Z������X^^ŝ�&W�sa]Ե�p��T`�I��f�+��v6/��aR���O;bG�%�h�����`K��X��d���h?u�|���4�"�u��+yC�س,��Mx��o̝�}�Ǖ����&�0�)�$���^�ɳv�u�K���.M�D���5}�������gM���[+$��v[/���"�I��h��w]�}g���N]�w2$��@�Zu��P.:�wf3��b}@������D1	���k(QS��s{uOx���p��Դ>{�ë�n\.�����#�"3�#,Z|�i@���x`m�LJ�M�B����kتӳs���m��0X�A��l@0�aD�Į�0�~��0�[��7����Á�2S�i�&:�vmo�i�?3��(��ϹAf]��B�|��-=�dc,�� G��+�*���TJ�53M��Z�9�&B�V'�r$<��ڐo��JRe���M�F���E?O��/fћ!5��fW�������9nP*e�U��"����6;��Ђ�2U`V�Z{�i ��4��g��У�/^� �� �{J��M�y8���^��͗;�B�L��}P�5ڊ�� Ņ.�e�T�2�5ຜ��YJ� 9l��L�de=h�]�����rt��g(4�@���.���4|��ϻb
�ax !�Y]����T؞)K������K_�g6�^�G����4W�6����wA�(��#�)[���g������z�a�M���U�*ӵ�?���Q�AP��|��|�P,�m�s�Ű���'�Vj�l4� �x懟T,#��+F��L��O����^�!1,������ɲ9"Iw�O�����9����Ui��t��@���m���S��k:sOTc7*8��}��v���u�����zi����Q"o9�=4>T蕬b{V���?�ԠP�����q�O��\n2��?w��f���+�-�=����p׭ �~���
/�k��A��ݱ���2�r�ǟp^ԨK{�Sô��8�
D��fX>x�>;{��0b�r2ܡ��`\���5I+莾��������֟4=���L�E[�E'w?�V/�"}�$H�V�؊�O���l~.�a��2VӍ�s����ኗ
E KG�v݆Fge!�n̿,d�,�y��o���ꑋY��k�]S��8����&�xg�W��WCG�v�42�Z��SC�����	
ڱ�d��u�uiN^�]��L�)������ኙ1̠��u�- ��9����,̸M��bb���ݭ��[�ڹ�p�^���������rٿ"JO?�^u�!����|��G�;���.~.7�r��OR�X.*���c[��*�	���?�,�M���wB�g5���Tf���z���sv�����Vπ���H����_����.�gF\f2�.�0pz˨.�|� �z�^:f��Z (��i�E�j����!G-3x��c��9Q[���kz�<�9�Ӿ�З����,'�Gtq=J�S��c|]�����Y ���;��?|�����$��p�cL�ԅ}8Y����I�B�^@S�:(ߥ��E �k��$�۽�{�E>����B��\P��ڑ�D���g�	踄X��%�!�h�2+� ��%��s�� �X�4��ZaUl {ST�,��C����br%[��z�nG�O �[Ԧj�.<B%:�����%�t�ѭ�5K��Ǘ<3�К���,����fE�ui�����"..<9e��[c�4��u^;�ȅ�+{�[7�KH>�QLt�l��lV�+�@/@����+�F�JA����9P��Ũ�֢9�k��d�(����)��i�G�� ��G�9`�Wt~�͓Z�E���H�\��!����~�Y��*�`$���ʡLY��2��[3�u�X�,П+B&<�VG�����O�s�?�����z��1��۳g�f����wb}G�eM���kқy^X�>��Ӣf��(�\{�sy,��6vT+���v?��*)�,?W�h�^�8ُ���$ ��o��-6�2�g��%*�jo��63;Vcv�����w#h),���ؗN��Ɖ���������`�{�9��2�
������OW6H�;N�\ u�tZ�Y������)��j�%��D��u��7,�_S[@ݪ9�`�.g=��=�H��U��k��B�/̊�K���"!���@�M�� �ޛE��-�ܭvl��Z_\HcP Q��R���~�S�-�r�_��Ujm=�.n�/��'����#т��/���������nra�=��z����b�h�@7��ܕG�.Ztb.lV�\��J����܎��~$�l�b�yV�ʎ�Zb:<��~��z!���K���B��y��	��7m:Xس>Oڒw+�ж��J��w��C��E	[SS:�<T-�U�����a��>�X�G�v
�h1�����쇊�"�!k�N�g��N�>RYX�'�W���|;��`>fӯ�p�W!��R��r3���$_��Ix*�X�ey���㉢xV�ݝ��%RO�~��"�&�w��<��gV��=�D��W�/R�:��������vB�|��3���~Pn휋/�a�g�O�a�LN���m�F�)��`Y*�R�ߝ�0�:���{��#��d:*,I���_�uP�n�'�}��f��Cy���+��no+~�'r�z���1ܫ�|$q5�$D}�U���)]��;���:!H��?�^7:e�tV�9�ś&>�$�\��&�2u�4	�R���K����v�7~�ڐ�����6~o�����$�Fp�aU�q���V�i{��;S������*���!u{��[��s;��j�c�d	��f��V�&[5���:� -���ocF��,��
�����}4�K�(X�f���-(�����W��V����57+|��~�U�|3�(��q3F�Ĵ���m[�G�0A�æ�x�����p��rč��;��_:3��t��p_�tj��?�x�+1i�7G��ޔ(��եy՘��?T��#��,i���l�!A#������8��B�o���?Җ_y���X�U�����p}�?��:,��{DAE�E@�AJRQ��.II��4�G�����Jb���$�`�y��<����xyy1g���}��^k�9@�}y7;Q4%��3�\d��{��_N�^���H�B���}YeX���A[�]峐'�|�`�Q�t� ~Om��.wP~���?��אv�T� ��;dږ,rDe���>�CN�A+?�y���si�,��%��n{<�9����%� �z��|�]s4�����ǝE>��a'4�w����@�b����H/�X����w�		��w��G��-�O�CK��9������8�8f��P��G͞���y��8�o����N\���C8!p)�XZ�f�r};��w�$������z�w�R�|�~����)Hv�����"��~[GGg8�pe�G�bz6h��_��q+�mY� �HA���?{�,
nE����;.�U�yrs��9D��U��>���T�Ĥ �,,��֨炵ۺU�}c��	��[<����FW;F��Eo��k�V�����՝��J���B �q��y�|�|S�D$ dθ��^���ɣFw�ݧ#�n�ē`�.����_ 	DO���K`�ɾQ�n�U��.$�|�:>B�d'bE�y��6���� ���m�W��v8���8/��D��]�`�Z�v�ی�:�f�?�6C��Z�YN�����
Џ�s0��s�Ah��}�� ʅ�ȩڋx2�4���홓x���ס"((�����Y����KST���(�� ���)������$��'�}�-�j爇�W�8pؗ�q��FvM�ģ, +�?�"�Lz{����%�漨�]���!Ga���^�D	�WeO��Ou{a��"���*��98t��!HV�exwP�k1�޿�y�~�N��YKE�D�����{b����E0C��r.wb�;�_�z=��o+�����J D�����R��r�
ѯ�Kɔ���,Ѐ�M�,��Fx5d�O��ѯ�zH��������l����R|<�V��+x�����Q�ӧ�������..[K���	��G�Y�@cQ7��2nm�+��ϧ���c��&v�:�����{��9.-�,SM����ҫW��h-�:�N�$;�3(k�������e��*�?�j��WZ7��(uHT�^��P����)�i������э�*=���K��/�rfڢ*���`uwO��)�7q�svW�'w�"'�9�DbwP��5Qk*���%*�$V��l��)f;��9{Jٳb��N�c&���,���I7�+��4s��p�b�cwm��E������)R�YςkJ��w���R�0��Ώֈ�xy]�C�@Z{ըw4n�7�����{����>���xS P8�}/"��wB6=ȇ�2�� )9��e:<����n�?C��\a�)w��� b�x��X���+���C��}��.����h����dw�;̡�F�����v��c��>��Κ�+��T��2�_5Y�:jE������Zj;�Alnr)�^x������[2{}r^e�[���1y��^�%�D#1��p���'�4��o��NI),�I����iHx�̸����6H���2�"���>���c��=S�����j��eW����e��0K.���"�:Wٓ�M���J,���1V�8�l��:�<4�@S`���s7���ZNlPKK��5�3;��!����g��ޗ_l-W�	��e�-�Dॖ�N6,��o|{���d�<�"���k��@r�����ƁCbخ��|�T1&��UN�7T%�Zak��VX�BBO�1��3�x��'����Y b\�@3�()鮑e�����N�Q��Z
��(��jCYWp�R�Oi�����;u�[�	[��$�K����$px:SH^��
U�Jt��{ �@2�Z�Y��3k�~JH��H�_h*#��xm��)���&�7���f����V$�U�
xl��y���WM��+=C��+�����ѸO��cw%��0GNw݀`�w|���|quS��`�'5�E���]vW��ĩ�	�K��̉IT���e��w,O`��,cG�����xKH;�x�W~]����P�}8����p����C�~o^�vnع���5
��2�Z�=ѵ��v����>��}v�1�L����q����sj�!.mΫM���/�S�J�����{U��0Z��g2ҙ�$jf%P/�%VP���O��8+��w��L�MX���8��w�A����aQ������5�C}�wJ����CTbי( �m�����Y�%��e��r���;��F3�$��EA�-�/�E7N@���&�]M(�C�E�"j�X�#��_Q�׆�x�"73Q>�%	���Z9�����sG���Y�1�9�wx�-���w<���-XOXVơa?�w�
1�e��+VA�49O{�#~�J�b�	��>�1��ןg*�������@��g]_�����L`��֔N���(�(�*�'�i<�3?�<�bp�EII��.>I��3���l5S��	œތQ���[fD}U�f��x/|Z�<ۢH�쇈�v�����\WU�2���qy'_Ֆ�Q�O#ݼTf�h;��a&A�x��Z�е�_�W<��h��]�7��&,�o�-�.��g]AA���ݼ��),�m��9c2�9������lP�f�I�y�w+�d�zr����0㗞������=�����Ft$��R�/�DC����Ą���7��jj;�����~g����xcj�7,��r>Np���9ahdc9 k���^xچb{n�c�O䔂N��	�p�ݨ�:bG�MA�bR&�B︗�[�5:�/�)�\�d*Y�'�{`�:F?8��S�P�e��V��V��\/�]#Ǣ�>����/���_��-�bf�����7�"R�I;]����Q
~c2��;���)�t��J�B��]bV��.�(|��<e��2fw�T8b/39� g�Aby��E�a�u\�2v9}8�8�����~��FY5�h�0�w Ȩ��+�A���51���J��ϓt�Z�;p�P_��b"��j���?�1���/��2����:9u����U�?]5��YTFu�mq���x�[��~^Z���X�����J�M�Z��]A��ԲL��5F4���Y��W5�!cq�,rq^�>�������3K�A�χ�jČO�u�\f����t�ݘ�Z�����>���QSY��W���N��գ�Cp!���dC��� *M
�X�P���XeKdP?Z��1P��CQ\�zG�lN���
~�ʯ˧�&�-��=)�m��%� �An=��������˲�w8Me	�����Hs+�o�V��*´�486ۀ70v}��g;fџq�Ӱ����f�)Gwj�`�խz��8R�gh>}S�KC�g�</d�
;S�����䯏��e+��'"��R�����,�e�bK�v�-PU���:�I���V�i���i��n� ���J��K�}�����\O��9�Y�^8l=`|&���_%�]��j��v�\�o�s�F#&�����0�g��@�����}=��w`�R�S�p��� ����?b��Io�])���Z�N�׊���`���sr��}
'yg�;�ٸ�\ʅ�.�
{W�Ϫx�H��07�v��%G�w����]��@"�R���+6�S4���\�<X��<PռB��N�TV�Jp�$�$=�P_?�q�9mɷ�N��}�����q$`.����un�}UG$�sGSՠ7O��A$y+^�K���\�~�|K��_��9��>M�:{���͂Ad��M��2O����Y\�������5�$��АW�/K���w�J��3��{�l��*4A{�|����^fS\��ɳuȬD��&���0��^����Y���M�	�Zf�������,g
Ҹid�;u,��'M~�p\a���D��v�!��k�X�9j'����D||Ӎ��x���Sq\�1G4�尠�Gʘq�mX�q�Cx�+�s֨�^lR�<3��Ь�<Eqݝ���҆�~U
g��]k$+�#p�o��=ӼW�&�R5va�!/򉰌C&�↯������B�~�ă��;�`0����GyEu�
��6�`Wt�2���Ts�6�v'��=����ә@�"c�w��쌺Ys*%�)A�L���!�7�0b�z��-�-2x���W���Xe�0ԉ�Ɉc�}��z?���G}w%%
{��/R�A��9� %:��j�����M��g��Q\)R�Mb�ų�]�aY�qT!��Ƅ�2<"W
q����%�WM����8��j�8��UvÛ�DA���*/���	�XA�홣h�z��Ԟ5n����ƔI��ry��<�i .μ�|���}֫0 ��I(���!b�<s����J��`���(�ӿ>U}a<j+1�s$$��#��Ӻ,4��߅}�[аע}��f�`��s}�6��;��M�3��$<�Б >�OQ_�y�Zԏl{��{�z�����
��9}9v��%+M$���p���E/����N��N��kL�C��H�Гn<cX�\���/�L�����O�Y8�pA�X�wp��~H-���\����pض,q�/'A�:�����V��5��:O�u�vG��8b�綦6{����R���w5I��<����l�j�ɧg�R��P~8����V����/e��t���w3p5u�@�g�ӡ�9�@,{��>.�I�����;{����"�Z�?��/s��@('���K�h �8w�K��)�-�`�uw8���"^	e[%~�W���q�(��\i�	�J�L}O�34�oPk{�;oࢴ��zN���We-����Т��S���%�¡�{)΅�ӧ�45�֩�҇�@��'�����]0�{-f}���>�:��}y��5i3�<O����a���rx:0���w׏��D���I��<�o��-��ځ*�lo��0����� ijz}��(�R�ng��d����$f�(���浑gf���;ļ��	+1�_=X��8Jb~���/Sf+Z��-z%�(�~,��ܓ�n��V��y��N�:�"���K����vW�C86#ޜ�a����`d��f�o̵��X34�g�JM��<�=1:��<��'"��jC��.����6�;[kyu���A5T�&�f��3K�$�:�<���~ؓ�a����F0�v�����)��~K�SV]k��@��s�: �'��qB�L��R�)�eII���נ�vKbȏ3!Rqhqw��sU��^����ZyI�\�k��,w���s}�v��5^ޛ+�Z}��q$
l�FL�U������
�sP�5w� �@ �fd��Uc��0O�/���Yh`�1����b'�n���=Ą�_2ߎ.�ogbFy���k��k����F�p+U��qy��m��m5v�=[S.U�%w���g�4��㋪v�P���}V����A��l��y��q|�}� �~����)fq�&)��?bbV��H�)*�v�	$Qp�yRC�k>,��q�ȴ�CnH�t�D�袡-�ӫ�Wi=�3U��$<}�'�J7dO��s:����T��j��� ����>81+����i��S\O6�;�BBE���3��g�C��ߒ����։<�{M%���*�@���O�6�E��|�Xp�z�i��4��x^��T���43ZZs1�}lD�>�K��~#��)�%v)�W�j�㇘`�
�TX���1�c����G���}wR��wܷ���ǄF�ϷX����r	l�8Ծ���78`�A�柚�i\�,wAW�vKH��M���͐��B}�.v�c�ԙ��7�+_����s��@�=	n=�d ����.y�V$�ׯ:�S�L���=6�N+Z�A�󘔔%���%[ِ��ND�,�(��f^���bgC�}|��W�<<$@>>�sU�Z�A�z���F��c-9�9d��m~g�^������Ξ���e6�s��}��0��EF�Y%�a*�� Y̛�{�rE-sn�{J+EI���k�AH��&�F(8�Dr�I�YX��ry��h_��k|5�ס����ָv�_��9̲̔?ix��]w��Ꮾ��K�^�A�ё�l���b�ui�'}�c�ʲ�������,y��A��������w`\�<`ld�G���NJA���7B�5^����Cc��([�޷�458}����:)-k��`��qGb]8�ɻ�2�6�5��
u��]�|�-T9M�w�m����^mT�ij�L.w��W}=��(3�@�X&k�hZ�Ϳk�og��4))(�(>`�&�z��Vj>C�x��~؛�5�a��\�d=/
2=�ʳ��ۆu9gS��\��R�z<�3ē0:{K����R��X�e�$
��>��Ii��b��X�_�0���Jӛ��{25##ug��4=�?:�XgG|�Av�kp�Khjn)�/�/������D��*Z��F��H3+��6�^��]�ޢ��%{u�%�l�%myM��c��K�h����w�C�����^�m��r�I|q��f�7�
�r�~F���;wB)|6z��-`KfS��õ��ʒy�n+s�����.^QZd��춓E�Y��WT��G�h��r\z��h�_1
@A-��އSW�\/ }������	2_�e�Tfi����n2���v�b)�Îu;u��.����r��v���Aibۻ�=�t�}�P���ۯU�K'�|m�)�:n�q�ʬi��Q�P3��R�I�7o����E��a��-���2VG�������q�)3��$��F�b���J��5̐��UTvTV8�Ȟ�:8���П��7��=�|�C�տK�,���X�k%��5�X\Y�y��;uqN۞��Sx&�+p��o��Lo�0lMLJ�` �ԘvǑ����`H�_�ў�f(ΰ���#��x�ksV>$d�ͽ㞰��JQV��#Z6�C_T_�|�  �T:H'mpl�m�]��u���Qѕ���C=�g�6����}�3i߻Uֽ� ��^�w�d��B����$��x\^���v4��26��_;qfk1��ˇ�7��W��t���,�gZ���ΕTf$�r�V8�ĔHoo@�/�-]�FS$1���#��.�a�/N-t���ר�_gnn����`1�{XB�{�H��cԡɤ6��
z�e`Э�bt���4|�#>��&��M��ZR���#�$5��Z���YB���A���b�7d!��^P����pe�`��m`o���ߊ��;Il��N���Գ�����ڗ���öRQ
�^x*���fb=���Ԝd@JT��	��#A��c�as�X��QzWG��v%���z��d��U�ڟh�H�|��h�M:�L[V������_珗{�o}+���BL�YS�_�̙��.�F�!S����N\���@,FD��K��{e%�&+�be�q�[��2mS��Qx:�)��Y"�@�D��k���-[�|�"�C����4��C�AC�)�[��<Ej���������	�,22[n|�
���)��[*/ {��O��MA�pm�e-��q[b1w�z��P��k����!�y�^[JZ�&e�l84`$�@����|z�~N�IH���.�w:�Ƃ
�;��JA'��ꩃ\���)���"g��<�ge�x�&�ֽ��&�D&�./��o�6��E^������gM�8���hA*��Q���͑r.�G�6b*	�
�X�$b�RC�<��#��B�W�]��N .T����xM��fߦ�c��J�:V���:띞���M��(�$�m�C�^�{Bi�I���>��q���7oj��*�;�vwo��^�h���6���v�Pt:��x��1��W���AQ�b�@�[n�C�^M���Ҿjj�4��d����^u�6:�8�E4+�����N��Ó/G�1�gUC�bbp?�e8��R��~�J����#�T�sv���Af�Hsy�{�>��Z���������}���o�[O�{�Bng�@��ᔡ߅q����?ȉY�+��B{3�����7J2?ɚz�����M�>r���׫̭���U���RD��kl�˭��'�XU�UWΫv+x|~$)�VOl9��R��Sw[��]�S �Z��XϥãI��n���"�;�U�P{�
'' ��M$��7_`�(�Փ��M/�;3%�eq�c����}x��j�A��p��ҏ��X���م�R0����P��.y��w!ZL�\�9IM�#M٫�7y���\�����N��YZpK\�����4%Z��>"�DrI�|yW�� �i�a�ŶNV��;:���է�
�a8Vi'b�QY�^Y���(I���lLW�9z�X�Ծ��r�ۣ��3xѴBP���JK��+f���5]�c�v�ݑ�]���W�F����R�X�%�0"�M:)vv�����#"�6��*vm���N�����ط�x|x�>�W��싦����/���9�+�����g<e�8ȂG��,��	����X!l������� �e�ݜ.a��NQe��s�����6&e�u� ;����A�{>�� H�=�֧������K�A��-#b0\';}��g�8<������p�*�;��O_��kW�K� ���7=r}N�EM��51��L��NYD�<+�|�.� ��V�J���>��0�:���R��1��ۓle��X���hkda�b|T��[�Pw�M�?�������xqj� B�cH�/ՠR��ZsߌYR�g,�斖�������ɑ�#����J.��҅w��
�����֞nJW�u��\׽�(A���½pF=G$#��D�����.Wt)[�aW
w�~��(ߜx����{T_iڮT؎�_�y���J�F�����|C����Q+}��
�ز}v��<��[�KK1�4}rvI���cC{��O�dq�C�>�h������V�xEݘ�|������#���('�P%�`WEUo2�p��Q�䴍U�/N:Npb�@�
sԻʭ���4��	��&/ ������ߋ��������t7��$��(G���W7��yH��x#�q"pKe"�%��'j5_��ks�'���D<6	}L�:.`�GP��5��.JJy@C��ᖤ�O����� �<5#�ظ�k�Z��5��Z���2[���d�DWyW�U���;�;QR���x��^�`�(�l��^��d�ڟ%���Y�@��რ˴��@Ա�Y�ch�tJ�x�R�R7zrjs������u���K��q�N�\i۱nq�S�(a�d�i]���4��Cv�?ޮY��bd8�L
Q����Ȃ�Ȯ������_%�ϝ�/�Q�\f��{�
�U��՞*y��f��a�6�@F%������U�D1os�+���R��E=��{�G9���+�lA5�z�ѱ�D���)Xtl�+xCQ�h|؝̹>f�Ha�O`��(/��Zg�66GZ%�&���~��
M`
Bed�b����MΔ�a����`qA �g+*�-�ndx�_~�����.3e���;o�������k2����p�	��>�2P�9V)�����-	��O,������Sz��i}�P|���ze��[wY4��mg7�C(�J���{�3�- C(a@qʫg�����;���3�V�N�*����Z���_tn�^e��'��~�����@ӥ"����ROv���Mi�g��#�����
jNO�����l�����b���7" AB����m����P0�(1|ېK��Rc{���a?�kܙ��t�_7�_5.�'���"�1!>>Z�N��"����G���+�<�[v���
��.����ևd]����+���	�Y~Xz�F|��S�Y���;�k�]45�qC�O��a3Ϗxy����dd��t��Ź�����L������ԅ|Gu����B'6W��.��j���t��h�i��a�U�����r��McuMs
u- jt����Ԍ�x@�y_'��;��YM0OO.������Q1c���E�V�>�? Қ3{8�"�8����L�ݿ0�J� ����HF�D�}�A�"�L��,������bQx�NO5m��?��q��x��ho]�;������ ���`����i�f�GwK��O�uV����ڲ}^ъZ�>2��W��Hu�`j����?�������uU&u���u�cBB	v�	��s�^ɜ*��!�y��b����#�ü5��ޠ����W}49j�It>��$ޟ�4����	Go�\��t����~���P���0n�|�n�*����Qp�٭�Ƒ˺��=�1�&Y��{�	k-�X�����H�o�-�e���diHAD�9^�8;O��һ�W�3y��*Pc9��iN�&NN^��.�'쾉�Xp�r�yK�'�S�_�n�:L��P!��#�(%w4�)jf����҉����Lz�d%Έ�6KT����y��I��A�௓]��NF��?T�)���o��bwM�	eXc3D�v?kc��������	�xpQ�||�� k�4H��h���{���I��Pcr��C��tֶV��n�=�W.��8,H@O�;�z�#�F��'}��@�dM{֧O 8�ө}��GB��|��*5�iI�u�B+K�ЦW��T�֐��d��)�i@��u����ǽ{�%���XL��;V}���OuI4#|f�b���G�T�7<���`������+��#�N�x)�������1�B����".����Zy�6�/Ga8�؟�f���f
�-�E�0�o�<R�w��ɝ��u����C������S%BUmJ`ؼs�X/Ǹ�<�verw�9��-H�P�|Ҋ��M�/@�S�{|�(@~�I�m�QI�M���Hy2�¨n���ʠ���(����E����'�*$����c�"�G�tw����e6C�%v)�oޔqj=���>p3����hJ�B�T�qH�� �����w2QX0~B�ˋ���j(�LJ�&��xE�i1OE)�;XG�i��C�_�H���5���%7߅�|D&� �jʜ�s�V�s1.2��#�O��l��:Y��#)X�ۏ����^�l�7 ܵ�����	�ZKsL��("��+|�t���e7�=^������L��z>��<���&����+��Nzk.;�e�:�^=�^I�˩5� >��4(O��{5���7��{%r�<EP��U��3o3��~��+��h.+�r
"��e	5�|
��5*҉��O;�Y�,ߓ��z�o���|Vjd�����o_�пc�^��,O��75��"`n��gz[�N��Q.{�@Z�Ίԍ=,b2��2��9CD�m�s���ط�˙���Ͻ��{��뵡���O��"�j�?����|F���Z�]�Vj|G8}�C�?�y�~0�����urpȣ�<��=Gz�Ma�r��ɚ� �4.a��&�C�_e���e/󱐌�_��,*�ɷ��Fx�F�J6bP,`��c���Uu T�(�[)V ��e�^����&�9�Up���7
��&JJr�9���Mp;�=G����Uq�v��eR�e771��b����i��
[��W�߫�?��i�6<lh��"��߻���w��a����h�	M[a�� q`��L6�ɯ�T)�����$c��$�X��#�`rR	���n
���G��ϓ�{�j����������񝇊�o�k��~�tY�*�	t�h&/;;4;Oz	R�,J�Jk����*3]LM��[iC#��}�F���`�aќ�����l�-�;�r\�bY�mn���b�w�H�*�b��f���VE~�6�s��R3T����PA{q��䪤�.�6���ꋶ+��M*�A$�=� %��#T�r[1�>ة��A��������ڍW�%��b�Q5�ggζ��[GT��%���M���h��q	�]��;PZfX�b�J[G	aW�Ԗ�A���6K��u	T���^��K����HI��!9�Ւ	�2Ȱ8U�}��jzdԢ���*.��nu���:���b�Ǯ��s�H�sn���#A����1"��wG~�7[i�2��p�]\��q�����e��wQ�R"��<�.�Y7��i� &�Z=��cz�a�$�J�n��f4�jCb#�ʽ���J{<'?��ԙ�D��#��Cu@��
c���5�� 6L]}�
��ǹqQ���|Pp���O Z�d�z0�����Vv�dem�q�+�Z�v-)V'Q��\g!?}��L�Z�t���~ ֽ���y�H''÷�k>�,T
��B�Y�MIR�����x����gAzca �����h{ �k�mR�H�IL�>�>�03�NɃ@B$�Zr!u�|�oJ��ϲ�z���Z�O֪�ZQ���=������SW��EObi�0bin�DD���'�x�+~Xӻ���{�'	�M>��b��"�����r���o�.����� ����7�V-F��,l�1����}g�6i;/�!ˍ�B�7�#Q_Qђ9�Ŀ��bN�Q����P׽�^�vo5p^�� ����M�������@p�"�)�߮7�=UO��*/a,z#muRu�5ϝ>��?Sb���ls�<�W��g
�(!W>N�R������3�u$-l_�:�D�F�p|dļ�e�7 <��B`��C�7�և7�'�駝���c������N~�<n���T��)nv"*��q��`�p����1�� 
A�E�X�Fj�E/�;�X���>c�)�e�h�nfθ,�gH�-��@�UyVY��� �����z�njKݡ��� [����q�~M^^]�7��/�<�㒖��&����
X�A��
% �a�#"6Y�����|[����7r�gβ��V?��F���ǥ�5MG��/��7��%����'%���|�EE�����v�� ��x��S2�ps�O�&�n�����;Q+�ݪ����r�؂�z�\����)9�d�|�kd��[���o���M5�y��hZ(mU�{���"���Vod%����`t�E��'eH�J��v����G�h�E3y�$Z��i�N
b��n�.;��̟>���PU�k&�ل�	�+���c�}??�˗��?�t�1鍾"�mm�������;�P ������
ğ��j���(C�:����J	�0��$P�\��t����ԙXV�q��뫂l���t�̿�v�tm�<���u�ģ�/)�����l�C��d�s�؀Q�mhi	�,h[+"�}��ң='�[��-���u��#���K���dL����j|X����� o�
'�7ߑq�o���<���A��\�aaDS+Z��=n)W��������J�b���U]��fH������~Csj�_�Z�nɯ�̓�}�HFG��h�'�n��w�DZSg�̈́�I��3�s�D���D��Y�v_r-���ȍ_��@�F�xn|h2���f�)Ĕ�k���S�m�ҬFIR��2�Kj�	$�CL�Y,��M(Ɇ���q�Op>��QH$'%大�����������KH{�l�i�����dm���M�t����b�*�u`�o���(��N�L+�O��u�A9X�9�B�11�d�1ƞ�ᰬ�
9�� �B�0��қ����X�X9�������Ⴙ؏�ۻ��b#�&VVb'�8gS�Ft[�x̾a�H������Jg辱o3ԁZ�_��%^n���N 2��j0�}�G����Q��]�u�Ժ��X�?�?�>&iFAäG��[�B`*d�i�����DKγy	ʎ��.�2����(*�ԧ_��aa���%>��/٩�8}RL�HK$dBY�!Q�j�1�:o[G�X\o௬��k�{������_5[����xB�	���]�T�#uQ��7��
9Z����QRǲϒ!T�7��Q�&6�o@w���(�z_�����=�Y/k��U����h{&(�^�;qI)c��܀��_T�p*R���`�����3yu�BuW��CBy� �'�eO�>$$�1�:�]�C[��_^�t�~�6�O�*�rT�F����ńA���
���5̈��6�w���A�>��RD�(W'x����IxS�x�-J�HҾ��)C����)��닉�k{�T=&>7��`��N�)��O��9(�VW�>�>�O���7s�h��I�l-^D��=뉨�(�~:\_�z	2�����6`��oQ�>�����rH���tKȿċ+��&���ƍ>��=���[��S�W�@�7�et������wΊ�p���>a!�0 5Z~�޷�Y'�$��`J��K/�����}n�R��6.��q�<|гU&�d���� �f�Ρ�F	p&��j��e�*��t'�d��_[��嗻C��H��"̃3T�u;���i�M8�B,��:��ji@�qn��b-�bq4F�Gl�kD����&'5tR�й�?T����9P1���܎���	ed��V4(5�[8��U�s�t�&��Y5�������@3]���;��U�V��zw��@��!Q\Y���q�?��޹/(�
4�<Mn��:1��0�oϳ���Q؆�������M{�F	ѣ �����ɣ`[d��.�ڂ0�l	)��ި�s���ūu&������a���r�I$�q����'�h5~��&��¨.8>�Jc���a�'�oE2#j�����"#S�ܜ�4JW���y�a�j����2eU����1<.J�8q�]�~����YS������q3F��A(L'���:��Wb����kFt����=b~�#��C�%(VĻ���q��g�4^O!A��\(�}+�X� �c�m�-)�uY���l������t��g��9���'.S�b*����M2!��d�G=��x����)�[��� wj��=	T(sֆ��6�ͻ�2S��MS�~Kym�������5{|�hv�n����c��~el�kt���[���U2!JX����}�k\��B/�B;:�%fr����E����+E|��~}"��V89���yN�W�㢹q��p��i���Zf�O��J<㹤Iy�c ����t'/�7J�GQ������~�k�1���;�·�0�ww�JkIΉژ/��X�3��ߛi��F-͙!�>�����I�O�t�,"��i�2�?J&����y��.��_7
����Z��#*tǯ�n���d�+(.�>��W�ϱ�#��x����/x(5��e��N�L�؃Z�*��yTQF�^���+��d��c���t!?�؆!�����.��R��q3#c(�A�P}T���8�YÙ㭝}���u7�vw��X�OF֗D˯zRU]�J2�����	.�k�����7��d,܄��]B �7��q�4{<ݬ�X$>�9Ua�:�N�`N�K�Nx�_���&Į�f7nP.M��p���B����pJ��@���!M�� 	��9������d�h��`}p�xr�P�ռw����y��^�-D%q}����QRH�ӈ��z��C(�b�B/� �����p�r�=���g}f�M�{�9jp�R%'FW9h�@�DF>>��˽Pu������H���li��L�b3���*/�,=�{c'�ؽD-ë,"�cS]��^F�ֱ�|�+Ц��Ih2m�����y�����h���,�� �w^��(��r��B�fz�\�X��3�N�B^��dH�����!F��k��z�l�Ǆ��R�ﴌ��"��ja���U�_��}�Z0��͖0���Mc��˙^{o�j(��۵��А�GJ�6b��������*Q���E� &.��'u%���7���c؏�vv/�ɔ/�/�|�O��ws ��6갇x���՛�����d*�[��%�D�]u�]nnb�U���I���a���hz��D?���4�eܨ�YyɃ����OdˋriΪ ~��~�{��I�B4� �wE.�40�/����m���kܿ��S&Xw�F-��hKM�a<p��W"Ȧ^���"�}����1�ReT�B
�w��]h'>}������io�����"\�W���M��[�n�˅�l}��r�`�]��߹;�	,E��E�O<����\���Q�sC�ĺ"������_�l�fA�Un�qj��Uf��In�Q�� �U��WP0a��^�}<�p,s�V�	��QN�:��f1C�DV6̫W-����(+�,�������*��>s�W:ȉ���?\�I�� �j���NA�D��¼_���٨�-�TJ� 7w�L��jWey�Ue�D�g�d
~c�=M��8H�J`��o9����XF&Y�x�x'�he�㴾�;��"-��z����|R(}=JY�<O%�0�ׅ��m�V�� Z2Oy��^�ӸnZ����vQ�j���ǳ��=ߍ��p��?��r�t���ӝH��/::�7��6U�) �5�t0�fD4�p�{�N��h�P����Um���vV�0���}������])���5T��<.��XRL�wZ�l��^�ܻl�\<uu��hX�J@��aV&���9�ql���O�	\�:�vMM͚��@���䆸�t4xW��~5�{^��\Y�����X��l�LH�R�ꂡK�07_��$2��N�|��J��N�l0�t�Ib#��p�۵�o7��8Ml�y͟�b��z��VT�:�k!:q%��خr^��4q/�17�f����v�WB��#)&�ݡWj�/P|Ȫ�E�E�]��0���I������ʢ�0�_�h
<A����]�`�S��K!�V8uB?@^�����\Mڶy�m~^IHi��J
�����r�(�|fHt�5HR�,�	��Y'ʖ�$��ՓhS��9�ݹ�6��C�ψ��М�5���.��4#Z�L1��e�`�l5�r���C'��yB;�>׫�م*�s5~sH8N�b�W{�O(�ƿ��jD0����ݚ�c��׊e���t�k�������8��Q/�z��vRkk]�����7ߍ�/�&����Q�HY�x��J�g�Y
h���b��Y��s�5q_��7g� r��������(t5�|�@\/ �Y�o'�7e�s4h�'y�Fߛ��as]RXK����>o��B��k�"���2T�� ����/��t����P؎d��{IHx)�H��mYm�p��c���[ګ�sj���dnwP0�M���M
��<��¨�c���6�H���dm�Od�����kA.c�T�7o��x�p��E6N�Ş�)V�'x�E�p�����-����1l�a�t�.kS�ܦ���^�~�!��� d��L@�ߏm�c�R��^[�#����|�;֕�G˚Y�Ϗ��	�vP�GG��F�����O`���Ӕ�]�͓��NMO7����i-.�s��cǒ��^�@��{
!N����-)as��Ň� \ ���M�u����O0CF�)i�>_�Ul^ao�����Kl�*l�艤/�۶W����&�LT��O���n��Sx��YYw�{������7{�g�:\]��Qk�;L��=K!4�����5�[[����1�z�_��3K}S����Žá;��	�g��8Ǆ��_��/2�����ꨨ���CRJJ�")�-�(�݈t���3��"-!)� 9�    �� 9� C|g���~k}���z]�9{��y��y�~�9>�B�PE�/��~����B��z6=��[������YcAHZFPE+���m�3_���}/N��ɮ��G%FUY����͎Q̡��̈����GS
�7s�&Q�p�Є{�ڢ;p:�d�J����� ��U������>�V��ރ�eȢ����_fF`⧵����}�o�7&W�RF�s���8UJ"�e��yw�׳b�����i@�WL}�P�0���;��(2�8q"I�hR{��y��-t��P<m����BWUi���W$�����s_��-�}�<��jb�����Ź���\�h�OO
D�t���S�T���^S�W�eˁ��7jxnV�z�r������ؿ�m�k
%�=`�u@2���F~����aBʞ��7I�Nc���pP^�|F	����C�~���R[SWr|��3d�rN�.�J05�67w���R ��X����n���`����q���F���@�C��<�1Uk��?�|�ϓX1 ���M�7�=��k�\�o��>��r������M ��wk�0�����%��f=�pA_H#wO�p#����ވ�+k�(X�,O%%�p,��R_�c���׮vq�Q�Sc���*���x�x^��.�P%��41W�SE3���ƪ� �|V�|6�=��E&j$.����j�`a���z~�
��t��0l��))���x�Dk�T����k� M�ب�|{��<�	�%��J���&�~�H~u�{T�6�@F���u�c;Rgɮ�:i���Ղ���Ћ߼�pY��9o�o� ��Iɚn�UEg��Ǌ`�������f�����!I��T ��oë��bT0��b�Z�ݪ�}ӎ����s9�#klbB	w���d��y�'Qm�&)���/D훹�/���;*���k��w�0�����Վ\�.�k��.ڴ������ݥ*RB�<�@y�|`�����pa"�v��r��Y��������-X��I��z��m\�� �zgY9gJո#{�eE����*zi�G���:b����j�'!,i�p�K�8st)���.����H�-��E�� ?�9���r��x[ٺ���g>�l�k��t�u��O��l>�%|�W�j���lN�6�E�������i�i������K���c  ɞ��"�.�"{�Ȗ;�[���
����K8�/�����0ֶ��4j4<�M{;��)��# �Mb���~4�����`fe�nQZ�B�;�����:8�}^Q�[+b\.E��qN��k
��B����冣�\����-P��衽��r����B�:z.L�N����t���H�d���������#UN:>u����ą�=e]H����5�?7�p��Wa��`�r���R�Q�
;�x�L�SO��0BO��W�'�XXb��q~��#�~����`~Fێ�:m�.��T�*C�t
?��t6.�S��	���=��+#�q��F��`^�w��;�cj�s�;�`ȷj���֔��������oQ���o.椒��ZS���tL�9%u���_
�������<$�t&��)з ��yƯ�E��#7�j�0N#�sr�p��c�+����=*�Q��>��Rn�G���)�N��g�HY6S�Q��66lB��D�m�Kd&6)��'���YcaG\�~��A8�����9pu�5;��F.��j����w1�=L"��C���&cB��@��ZQ������-��$
"��y4��]�T`Y�����Zh��ځ�g�ô�LBɢ؄D��VY��r����y��w".�5x�1FUo�T|8�tLLrr|�zst`��1��SI��i���;��$^\^��� )R�C�%z��1U�&T&*�=�BW���6���k|T�l�Fn��
N�L�zg+��'�*ѝ���$<eB|�2�O����bK!�:Ĩ�WnOm=�����nɊ��5j�B~������v}ĈOt�vg�p�颫��iCa������0�3Ά���g	�џ��5~ĳ���7����t�"ID/M6��a$N�p�.��|��
Bl$���\1t$�L�!����	I�� b�{Z�>��ό�eX-�U��H���L����&8������	�<y����˅�S⻨����oڧ�t�� ����vt��#m}R���oB"�I�����{����JJc�ՁgV����|�O�%9m�q���8�k]f��Y"�
j>˰�ֲ�W$TV�*��^��)����I��b#��ސ�~�����Ol+���O���n~�L�74U���$�����ʫ���O�����|�*�[D��i�z��q�o�3���,c��#"O����/������vʖ+@�
bIket�������qZǙ���J��j8�j�-gF�Vl^(���ߗKJ)�t���]X؊�WJ, -��WѾwo�+��3s[lJL�z<>1n�1������gCw�tf�̆W�@����~I��t�_�nn��.辵� ���q�cĞ
�h�TQN��~�^4��x�}��S{�q��U����Q�U|ٱ��Wh��g}F�Zh�-����ܒv�Q��0�m|?�����g�Ʉ=9�͢��Nl���eˑ@�}����J;�~l�6qˋvdf� &4��J�+zä�S��ۻë��|���l��������u�$��%�����2����[����s��JDH�p�����Wǁ�ǧ�g2�)���% ����w�`*�5��j�*-����k����ӊ�?�lH��lU���ϐ����O�T�%����n}Ya�"a�#+�C�T�嫇�-`�،y��/�	g��X�1 "�,ʼPP����J����u�1�zd&u��]����95���Q�,�w��7/f��~'ݎ���b�a^���͒�.�>l^�n��Ȭ�fnO�E�z�A��2/<�	p���{EA蹌)Ɉ�c ɨ����O����k����/�*!�+XRĴ�'�NOFn�E=ÞbtC����ǘ���J�ts�5K�*�����CeR����XJEt(mgm��u}q�����Ug��
�;z�8N�9���{{Ka���>�ۺ��7|����d0D��HI�o�PM�N�M���]�L�o����Ѽ�nt�@{\I�'�Y�/�a��w�_E��Ȟ����_�B�5]�b���xf�h�;���Y��a���5ܴ�g��v5�'8���w�#��E-Y�	��WU�{��h�M���UQa��#5�F[����A�n�N���	F '����:����&�y��.\��0Hlr>�il^֮o�Wݒj��Lm�pf��n��A�U��d��שDad�2����Z�Jg��{ڣ���As0�;�zy�_���:�6���ɦ�5r|�B��#�<��$�m��&����K^�rYЌ�#�!y���f�Nɝ�tT�A\s�uּ�z	K����ȸ��ۉX�>�ӏLJ?�aS�P�j�&��^s�/��*�N��D6�w�v�]$��YŮ'G�����J�T^��)l�X�=2ʢ�u����*���VDm�	�{��gi���#+I�B���UE1���l�r�A���#w:['�ϼ�K�޾&��d������ϳ'������$��.{���/�}�9�C�S{�ZB�;g"�\�y��*����r1r�lC�@6��y�gX�����f�\)�q��ʹO�]%F�}|jW��1��ڒD�дZjY�`j���5����S�T}����ԀAU8�����?����΁3�=���w��W�j��sd)�7]��qT��b��HLJ�EE��}��I|�pÑ]'�b�_���.����PH�_�u{j׫"k}<��k8\})�'��U<p��������r�����(*��N�#�/�����th�*4n`���y	&,6��bVEa���$�u���w��N����ﯺT�2����w` a1"����������_ճ�,�=�t�1ޡr�=8��H�����t��Pj�N`�4�$��ǧү2�1�k���uS?cr�sw�ϫ�?�x��w��
"����~������z�Ycj��2/��)&2�'�
�'�L�Ʀ�����R�y��Z���3~��ձ��؈0�E[���8�֟���
����M��L�ݰ"s.�Ha�?̢�R/uNW�y�� ����Ͽd���t�n��6!�oRa�vR����\�Q�����9�n%�]w�Q�����M�Q�1m�
�1�-��5���ȿ�b�A���l_�F�ܵ���Q:u��n��o�Uc2�o�@Z�J�NB�����A�*��8���{8<�>��&�В�M��c��.?�B,g|߄�8,eN�}�X��X�?j������Ak~�o��a��"�X�{ ���`�������з���K_a�B��Rj�����f�yO$��; 
)VJy�C1�n��u���Rs� � ��ox���sb�u��E�b���ZC�O��N�{���22�)��,����(�~f��{Bʨ�M]6/Ɗ/�H쫐1��=�'K,��=���tv�q^���r�\, (�gIs�Ѩ�zF�eE���(B�ʖoV��P��HP��\w���-�r�6!�;8%���\Yg�g5:;���*��QD�$Dd ��@�,��l��[!����EIgf��ԝږMޝa,�0�/�в`V⊪ǽ��4�Yسb�z�+O�F��q���J�c�S.W�6���ΟL(�v��{ojwS�&m���F}{a���O�Ur$Ȟ�����E���1������%yr��1�����N�bN8�W^L$o�ǘT�����	�G�c�^Y��!!H3�Ca� �qz�|�W��o�+�;�U�:���w� l����͠{�����
 q�N{�q:����t�k��cf
"D依Ea��VU��z�	\ȑ�h1��1�ۻ�pnCja�_1�囱gO�G�L�<T���0q2�+�/9�V���$�$3�χ[]�7/y_�:F�FF�c�}d!/���z��r3}��vGg��z�ZA;r�Ǻ����[W�K5+^��zPT;鸬k��0������j��Y��l�c||�ar�:a�r����� VW���zaj��U2�̱
�=��|Ӭȼ�hb"�@�^�Fm�0��"��!��QR�bE�Mof�� ��l�5orB�W���6����I;�G�����zДx��
�{p�M���Xr��
�"u1C�]|Z��|9A�2�v���`�)1�-P.���	g�%K����g:X�ь�>,TU-˔������M�4[̭*�*,@2����ah�U�qؕc���ی�7&z�KiK��M<��8ڞE�t�=5H�E�|��d�0��y�-�W��s��{�6!�|��ˣ��� �p$����1 f�✦ �@J���J�����;*w�t�0T�=�wB�_�wڤ�I��7�R�z|>���� ǹ/���|�}�E�'t&5���l׏�������^^�x͇u�+l��U�y811��}�r
=��1���w�t-0TG<�7�9Ѓ���ic�`���>���S��`ⱖ$���u�Ԫ�0�xo��M��M*����^p�KH��;���{�L?�*���&q���h_)�V@�bǏ�2e�۸lc��K�Լk�[>[�>;m����9i0�r<j�K{U�6ѻ���bγ5�5�G�l5���ܤ��$� ��vh]��d��/��둪�� ��RXׇ읈��.��s�7�[��?��
M�ȍ���g��Aw�u�#�4�~g��Tk����>E�Ct�g�8G;�����c��x);�ɘ�������x��xV2Q�9�$u>(:��
��U� Y�NT�t~�r���F����@����H�@�^�_:���n9�;����L������ڈ�_��4�!o���KQ��|��しoUf!o�S����ӺeG�n����ӯH���t�����R;��QD�}��|��ba����/��#amȧ~�6�f���ӓq1ku��M��/�<MJ���:�.�Z��\s���͉��e�bַ���v�����H�g��n��ϲ��υk3J��#��`?������pw��.{XeTe1�zz�R��̢�@P�Jg��z�իN�\�b2Z��,�8�1_l�^�ϛ���wRBe�d�%��ѷRR�L���Ժ~�čǘ��x��kG��Q
�����+� ���8ʐ?/�M=)g���,<��@�Y��B��������r���ݶ�B&�Ю��WY��5ϳ�k�@-Կ�� r�N��bd�UN�Օ�c9e��>�U�S�M�G*�I�Ŏ����P/��k�䰟~8'$�:1��wRΫ���\\|���#�NkLo��������?;Sܬ�I)\ّ��Y����n��%����}�庡`
Z����S/��Qi��F_�z!�-�<�A˴wI�����s�S������l�6j�s����>��p&&
J3�W:M�$u�2�k-�cn�bO` �,���Sz�3�;�W-_�\�'6�i� ���x�s�F#�1�e3��:���y�s\1&M�`�Z�w|�n���m|{��ԗ�����P1O��N3��3�GR�Ľ���@�����1����ˏ���� <��AI�\m���b�}�K.�b�T�S��g���(;b�~~��>�;�����F��߶�����ep�MH����<j�l+5EI��{w�i�A�e���Qz���,�|(2_�0q��ycڌ'E[���+�U������{~��V_�u~L��(�]�+�����w�d����%���q'm��`�+^!q\���Գ�+��%*� ��Ə��/�N�Ο��i�=@gG9Gu� ��p]�5(�Z��Uߟ��©��é9�M��&i��g��3Ry/��w�f�v���[u�������A
����>	�]��+��g�|t#G�Tk�2�p��NQ5�_{��r8�H���=eװ��NՁ�23��q
�J���K�/�\=T[�!���T���tA��S6�bK$gr������J�y�b��F��k]�gj�
�o�d�#��HCcq�>��U��Ԑ�M��	
�������x��-m�|���^���kz�A�k�t��d���b
Bk��*������g���2~L%L��\����j����$�����H��!A�T�m�ϡ\[�z$L��J���\Tz�:Rc�����LƳ�+�lK�J ���3z�R(�>�,i�+\�SF��o�yD�\���=IZ�M)A�"V4�`~d�e=�Q�ŗ).�%������T_��Z�~�Z��d��"2�J��N�L�ю(��k����S� rașTy��R��z�l����Y*2AJd���tZ�(<[䓰G�i%�����N�N3�-p������]�@fD��l�ʣO|��v���� ܇����v�d��6����� �k��)���"��ba	�3�gr�Qҥ���1+���7�'�1z"YT$˾^
�ޗ�C��ֈ�77�%n;'���LHX�0�5����փ�#\��?2F��Ea�`�E<EE��8'���g�t���������|j�UCra�6�kNV���.S;/�#��'�������:���;�L����s�^h�b��ՕX���G����eϳ++�]Q�A��4@��	�:�ʟ)o���|H"�>m��A�I���,�^˖�[/���j8
�T"���/�|�$��͹��2ڏ�Y��Z?�;e��Qg��4�nT0�_%���w� Ỹ��u�Nc�%�^�r&Ϲ���i�|+�n^�G�)�&��b6�gԌ���Կ�7������9X~Ƌ�1�3ry�Mm��m��K��8O.�#�;n�4�tȇ]�:3.Nmߞ+x���� x�<��v&<�:����v�z�߁ؖk	��9�^]7�l�J\O;m��3�t7�;���vw�4�ţw�g[��7p�+���^�
<Co7ST�lix���$0Ya�(�F��X�D,<�S_��Uf�vA��i�B3�Po��H�/Z�����ŕ��-w��	,`��ԋ�J>.yfO3O�Y;y�zI��[0}گ�GU���^�80i*��[>*�/���+\� ����1P�l���ӥ������i��p���"ے6�П.����L�5]�t�� �6�<$n�)m�/c��)���G_���X�ߏ�w�:�=�m�d�'�.���������着D"��)h�<"�%���N��hh�Kq\.�ё��o�(�Z����䋞��mww�I�p��xֿw$`b'ӛ�6�o����4��t�Cb_5�j�F���N8A%=�h_p���5��-[V!��-Al3�ٍ+)��߆�gk�Qawvs�Bg~��'m��Mt������}�>�1�[0Zb@:00޸��p��d��ϲe� ������k?a9S��/��e&�����.>�)"�B�h{U�`e���k ��V��kk!��-�� M�Љ�cr �>%�z���o��j�����u��,��x��ͥ
�4J���n}v�v6/�ʎOw��,�u&� ��T�rd�;�	1�-������>��o$(��y�Vڨ@ޓϲ?����F��w\	r�{ LgMv0^��o5@ެ�\�����!*R��9�g�	��?LM	_3#�ƑKǧ#b�mz��y��ʀb�o�p�	=*�@����5/�c���ۓͥlS�	3�K.�7XS�ү�9���tTAhu,��lNԟR������n�;=Z���ÿ����R?��۫D�@�?bm� 966bB���aP���)E��_�!��f?[�X��{�S��e�u=7kB\��*�H�_%6�M����0���eS*�C@4�J�R����Q��B�1�9a��x ��i�
�ߡ�} MQ65E ���h��/��a��;����{�^"����΋�/㍅s��e9$	A�&�AM�UU����-|*<ch/��T~��K-����BoPT;D3'��O/vbq!��F�����M�BN/��Oo�O5��BG39v^Z<���������{<0��Lb �S���D�2��4NP�R��F�!$�j6%���R����<D�a����)5�Haӧ���?pvsT�M1�ФF=1U��B�5����ݣ����3(��HU��p
S�l�(�;o㎫�|�-�N��(��.����smT�NN����YK$[H�o>�m$��4A�C@+$��r��ﷀ80��44t$�wS&�����M7���Sl͔�k@��'�[�*O��0����6�G$D}�B���Ћ�^�����Ɲp�D�����4��$2z�W&��ZK����iX�G2<����%�!��m��@f�4����Ab�q?��6^��ז6 W��Hm�d�B�}�W{,�U�  W
�)�ץ��F���	�)H����C���DN�)���g~�
�n�r������K�zğ{V(�E�J+��[S$�;>�2ܤV�!��|�n�ǯu�20`��йR%�7O�J�<��vT������iEʷ[����gk�{
��<�{~�Ϯ�;�n���_]}��ߝ`L�W!ߧ����x� �L��yT��x�����w��n`�d]�U�r.���)k�tv��n��c�2ڏV� ��?�"5�6��:hŵ���q!��ԛQpp��
��[c�V9��G��cO���ߏ�ʎ0��[�ޫ�c}R�ȫ��Y_� F ���Ϫ���NA^�Թ��`�BtXA^�B�h����B��%����y�J�=��)쒱�r��"�[�9��1xt�r�wJ<�й��h�:���iW�p�9���YU�A����t��ªc�����?����p�Y�w���S�e��i��t���3�>�q��f�-8/q�����S�zl�.��"7�jEF��K��#��+��}�>ݜ9��t�6R�J�ݷ{�����Rqg�'w���@K�{.�@h��sr^�`aBf�&N~+(�[����P�����c�\��{12�H
��@�j7�������i_RO�)�̆y�=
��)��Y`��[{sO�(�O�X�%#F�6��آڟ.C@B��
��cMZ
��#3s|P���	8M���VXOʐ��^�;\�Ь�$�8�ͷ�"uʮh���z�>5�/��ه\~�e~_�q_����z���?��<PDۈ-��EvR'���\8}@���,n�_X���ߪ7`���m��v��/���n�ߴ�d)u�_�EU_D�����Y=��ˑ�X�c�u�}s��H�t<72�p��V�X�u���p9����9hu���� �M&�p|iȝ)o���`�Zտ�DR��`��Z8́v	�mkj+=r�q0�Y�<P��h��Ňp�m	��d,Q'�[SΈ�s�"��}I�����%�d����D��S�>�.F!ї�����'�\���@��p�̥�&A�GV�kkA�Ʒ�o����&$�I�H5^oo�ET��K4��q�7�nKmѓ-�n�p��8X9�k6��yi��h7w��?�i�ЙKy���Kr	��[Q�-��m�_�B��Fz}#������� ۫���A������ܕ��>�_RJhb�iȏ������VP{6J�+0/�__�O��f��Y������&���"��cw��I�>o��HШ�ۋ���Eɕ��H�j)��6*哤&ѵ�`/��1���):�y�yW�p9�����e6�z��GM��y��S�ͨ���,J�(7���[���ۿ�-�iͺ��V�BrU�G�VΝz ʴ�w+y�CZ}ՏQ�W��+��O�ߌ����CPQ1���D�3�aX�ۤΌ�Y���زd;ܠ$�(%
�92&n�e �OHv�tNT����r��h͐�ԓ��x�`_��P�Ḕ�1����*����` A�)>[z�#�g�#c	��^-+Z jd�,�� j5���L�H=A��]�'k@l[���a� roW�����н���i4"��Ƽ�g0.�w�&r��) �E#%��69o2��u�画0��-H4!}Ɯ[��L`��/���[p�ap�,�L�lX��b8#c����ZV�I��x��Q��Ol��Hl-�%$�_`�}���ܬ�X�y������硔ܾ��~W���c����'5��ӭXV��}���$�^��~��>�-$�=I�2.�Oy�^$ KE:OF��'ٵc �5��2�@܉ޏ�Ы�fm;�����T�mH$u�S�y�ү�S�|�Q!|-^�`Cb@.�O�~օQ�΅��\n�ն�!��� ~ H�����G_Z�/�,�^��M�3���#�g:S�WЋ�#�#gp���1)2��������`�Y�L!�����;��ͮv�ՙѮ��4���!�cD��Cy�h��/�E�a�L��b 9H�c!��=���n���e�юq��l)��5���������􏩃Ǻ���b3�@_���?i�������Z�xR�����R�w�>�c"���(�U.��푒&��.ZA�1qD��;
h-8�V�$�6!;�f��O[-�<-:�ͫ��\�g�ƒ�a�<]7	&X:����^<��{����{tBfq�eM0Ú땄f&*�TW�u�?� ��R��8�F���mL[�67t=�n��cN�����D����� �-yQ"8w+�y ��H7��^GN/�@&��emS�	r���J��mU��x�o������ ��o�s�W���	���qaP�c�� -Fn2��ꍚR;����ށޔ<j�W�4OL�HLZ
�������b�j�b�ni~ΰ�3���2�\l��l���[�J���۪C����H];�;��  ���AWװvWڗ����%�]|�3�����^�][T�v��7���_j�Q'�g.�3p����9��v ��;5��'����oIo���ؔ@�14��ǿ;B��i-O��ׯ����X���3��z�Й����]��p������$��3�^�{"|����j�[i�3?g��;���o*��"�م����U%%R������6�nc`x����IÌH�ו﷈wHpo%�O�@��Ҕ�� D�;V�.d�C�%��� ���dŗ���Q���f��7�<�6���ʣ��-�5��]P�jgD�K(�7�r*ͥ���z�}��zc�׌�����R����p�x�!AD�=���Y��r�Z�ٶ� ��г���"�32ğ���Y�j����)#� ����'��ک�#�G�x���~�!��]Q>�7L���̣J�`����:*�'��OM���-��çV�.8�#Y�Kϟ��[��_'m0�V&`���?j�,����ro�f3t�]��?dz�o�aO���Y�V±r��h�	�;�1p9�֜��%��&�()�e��?����.��j�+�"D����X���P�8|A�0%娆 ��#c5��%W�v�%���&gZ�+�H�q�� �e�[5��%I!������P>2gĜ-d6��1��C�;K�JsK4:��Oho_x�m����q��afv�#X�O�ٟ��m���U��)�I����Q�/��`o^e��y����5�\�������; �������P�E���Ku�ׂ�nхsa�t����0�ސJ>5f���.n�N�֐$ :��셈�*\��x���L8�Z`Ϛׇ��9��2ľ[{��<܇��2��07�:%��T��Y�G�fR��.��ES\���B�Qh툉��EI�痧���»���m!r0���R��iu�ϛ��q�@7�pd�q�ФQ@`&�j
!|��*j������Ǯ�����u�V����r̲<<��Hۚ8�O`��{t�#�85��/��ǉ�8��A����=_���1/׳pj�:O�� |s��o�d�.�^���77��&+Z���SJ�ƴ���J���N�W�R��z����''�O�X��P'A���n�۩�Z7��<^a��I���lU�����k:���*��Ȟ����P��=����Nj��GZ�A��cՀH8�=ݍ�QBb�Ao��L��cp�X��EY�.��=Ø�g>��O8���L��l�`�	���${BW�����Kw}D�kZ��<+]�Nυ���;]!["�Ϡ��B@��:�|聘xE���+)NA�r(�s�=58��1-[!�Ng���1 H�'��|)�M�����?�b����YSN�����1�vEx�sP.��sPZ��x������ssm�l����`������xr�o-8�<l�ɦ�}{W��LX�X�l,(9突:�o�6����#��kF�R�����q��"�r��2��	�h)!5�!�" Of�&y�� ���\���V����kd^z��h������A�OK&�B�x�k�A�%)���C�N:[���A�1}H)MG���z��X#K(<o�c�����ж������0qՉB�?�[^����@rYT��Gc)u�-3_η[%�F$=�����s7߹��զ�]��n���q�:�u��E&X��|ď�k��*��B��>8#[ջ�1&$$�;6�"�.a	���
2���kO��ft"��fe�~4MS�S{9j��;�����bn�J�M`9����r�}��#�+i.]�����>��KJ%4�ZJ�?C�1���QT��@��>�l3�~��!XO�o`
r���������Q������|d�2�x�����(�6��V��n?���
y9�F��"g����΁-x�q'�B�}��烳��C��HA�������F�z VAΥ[�4�#)�����at��@YT���������c����f�G��vD�b�����xI�`�[�4�i|��x�{�;����U������kC�Ho��FNj�������6@*�"y\��U�;��4��Z����i�g�N�oJ4	H5�"m�,MG/��^����^����v8��~4�s�tL\^ϔE@O=./p ��67����=���p!Gߞ�ҹ�z�N��Np�i�R�5��)�5���#�fC����uǅ4��ʈ;y��]��s�0\�n�܅Dbp�u
a����Op�9c�P�����@����p���⁹�K�Ƭ'NꍷF�����V��,i���X��`\��rj�;3�W]vU��*? ^=�����T�����F"�ޒv�z_����DrX?�>V�����5o���~�&p�����Aߺ�'R��p�"gL��gB�.o(��_i�<bM���F���B����]�]Ӯ���o�X1᫸�LD�V�+������R�__�wq�U]�I�2BB)+�{R�<�Μ��]�x]�H�nBm]�����{�ɮr�h����X��H��ľgƀ��<��,Ϛ���R!��+X��Y�d�9|eG���s�K>!ê��8
N�k��-�� Ζ�󭬞�����Q��1g	.�R�l�*��Z�U»��� ��a�&Xv_Y
���|��&Vĩ0O�Bg��Gf����GD�像�Boj8��8単4�J�͋��L��)����3�=��,Kd���=����_�m�Ʉ������H�_�"��:�p�y������c��{Gk:tՊ_ޞ�"�#��)����M�{V~HZ��׋X�Az,Hl��1c�߱���If�G�3C�t.Ժ�U$�7���͖(��ԈI���8��$��8f��ԗ��_�(��|~����e�OG�Eo$�e�A�̼�hs�&0f��pF\\k gq��t+	��J������0+wA��@�]��h�s/F��0a�8�2�R�-j�e�X����x�ѽ�	TnՐ��z��D���w.��rR��L-����@�ĳA�͆����o��]E�Y)��1��".�t%���c��4�b��0����4��8��"�rpvt$��'%��`������_�:��#�J��V.�nY�������N�q�?��L�7�P-I�`B`�N�:~l�,�F伡.����#�͠ �Ws�|``5幰�])��f��Ø���t�&u`�4S ���U�����}6�7��Ō����*�G���Ƿ�rᓭ)~V�'3 �"�F�0����Չ���@
70���~ȞJZ���j�${f/2V�xﲨX��j~d~��_�5ԭ��΃�@�;�^�#��|��bs����/�����B_r����;.h��v�����7�\��T�$Y��I�Ĳk�[����D;����2�N��ͳ� �u�՘gAg?R��t�̲?�/H����_}-�U郎�\���S���*��.�w�K�հ��쨣�ѷY� ���Nɱ��4}�b���~i-/�d�^�Qͣ�(uv��39E� �����5�6`�y�\���P���+�i����??	'�IP�M�����涚�eּ��,P��ޫ���?c����;�T������z�v� ����D�pך���x˙sy����mb��O�<��i��>j�	&�y�^�N�بgk���$�t��7r��J���\��\�յ��KK�
M�{33MPT�<>^���@�ۯp� ����%�vf[�)偝Ebb��o�ž�Vb��̏��W�\}�B&�'+�Bx�a���Ow�Ծ��o,�������M����G4���
ڝ�������_0G�����"��<�Q�w}g�Py��?�ž�h�sM�z� )\��<!l��B�װl>�z��PJ;\*r�ߋRk:?�����3��	Zm
{�7�1?����̱ٙ�ة�LtM��[?I�/h�W�jI���@�u�;�5Ew�z
�^�� ��S.}%M�6�)9�w��}��$����o΍F���LW�� �L�zń^z���P�q�⺵ԕ�+H�Ry���@�[>��Gv�L[�(�g��;q����?R�G
X�-zE!^>�K�������{�k�q����%e�1�4�Q��h�k�;��A�:�pb��l�8�8dH+UM�O{���8(��sb�G;b�N]�o�l���>�?]�[���]�I�(��Em ��i��G�\���uc#����U�F}�����b�i�Q�>	H҈ɅA����
*�O.<|�f����������8WZ����2s�^��ptzt��xؒ��/'cY��z�$���x��\�����嶐�G=u�A��)�����A���oȵ��5����]�7�
�.a!��X�N�I�{��t?�K�;;x�hg7}��2ᐺǸ��ׯ&�]�oG�Q7�v]�ŴG�%�U�i�{Vjp������xD��u�ErvR�Y�� `?AHid�,�� R�~�I]5� wEu)����^�u^I��V���RHFM��r�R_j_�-jyOW��U�k��W��+��5�=���X�l@����ۏ�1�J�C�o������a��l��d���l`�B�{-V+;�
��L��5��C�3愴����Q�W" L5EŽݘ��U��w�/�%�4_Y1��s%7ކ�R���0�I��^V�L�Cu{*�v� �g�+��w����3� !�� �c�n�r��
e�ـ]m��m�Kx�ir��Ŀ����%��`�#�@,�G�!��tEvYd�p'_2yh8�q�q�����HA�P�����tF]@zgΦ���g��&,��ס������2�i�t�L������mt���x��$n"CsO�e��!x��CWdU���C�Ψu+���u��%.��8�7m�i�4ҿ�g��<�)����l�o$�����K��a ]�����P��t�X��2��q���*S+��]���m7����S�&�'��8^��Q/��x�1<,S<�>T�5�^>�&J�k|̻�ru2����m<�2{�ǃ����mR�-���Gq�{ܼ�������z�޽�%4=[�[98�h��W4�����'����f���U�.O�%�6�4�56tL�}�n%� �̶����m�%2��筰3�uX=�$����k��iJ��H��ۏ����V�z������:�3)y���$^9��g�x���Q �3�;�3�#F��΍�f�4^�;5G��;k9%&�> y�#�h\����B��W�}N=tx��
ĩ�Dj���
qa��&���D�����aM�]�p\��Ea]�""J�^�G���ґ�Kh��(u�5�D@@@zOP�K�:��BK��L�}�x��}?���t23gN��}��Mfr��2�Tl��zΉ}^�S�j6�u2alr�2�X˕#��������L���'�t�@�n�ʀ���iq���@>Z9N@�3���6��h?'�Ӯ&a��H�O	����a|gO��\E����ʇ�q8X�9���*�R������ӐC�1ev�)����4�X�o�9�K	���!
+�WoO�l~"|:?p�s��Y�ȫJ�{�4��yz2+��^WA�
eQg���K�wE�V�Q7����sH�._-'��/ �^\�5�󹾯r��v�yN�>{��M����Ҍ1?Y��X��"2}[�~�ҭ=��t��f�D`a���՜��l.��-s\QY$�KJF�٢�ܲ7j�Y�����8���*��]��zz�.�yM����=����tqV�����v-���x�{6Z��ʗ�̝V}�A:�OfV��>yf�c��5Bz]jm:��ܹ��|k�Z㽫�n�� $>}"u����m�����pFf&�;6p�����Ȍ�{%�2�&8��!���a>������R�c�Jv6Jv�dg��Hֵ��d����3[U�`(�gȔ�����������fz�� Y�E���N<CS����=0���s��~���q��ʵ��Y?\i�u�w�*�8`溯8��`�K�M��ޭqT��᪡/�u&]l_A�X���e|Y_=i2Ns��i�������Hc<�n�t]��K�Z�3��9�;6��ǳ�'>��:χ�,+��ȶ0�~"2�8��:.��R-�2�Z�#��|��ҋ���+�o��6��l�>/�Ђ�w��,��}�A�@�!�xb���c0+$��:�8�Y���~����1�=-�V	���w����%u Yx{M<�2�j%W}�{:�1���d9��$ĕ�X#��²��:+��I���B�</8��Ռ����ȸ���y� r�O1��d��؜�L���fzg�~W��,݁>&�~z���#^�5G֐�[���#6{7]^N� ���w�Vp3�X��Tr�Oʫ����z�Z#95kē
0�镃�	?�78P�==��W��3us7�I�ە�Z��?qM�"_��H�O�e{�0f�t�bf�`f�����pn�����/E��?�e��z�I�f���wŗ�@:��N�r�H#�2�TJG�|X��R�O��!��@l�h8`�BL��e�vC��Yi�/޺y*n��)t-��₨G@�1�1r�������~�ͣ�1��n[��Vz��T&7 M�o�2fr2f��4O?��҃<��*k�j�D�Ʒ�_)�?�E����B�?m����z�x�TNn��i�N+p��%��m��X�>��B��`oq��T��l��F�nL�6��N�ʗ{�Én���_WۡBPg�����6i堾e�s��#e�Yj������E|�*m���4G��ϫ-��;�$�;p¯[����ٗT%���c�%��P"�"cNwbp��K�����(���E=��]8O\�������������嶟��K��b���.�7�����n�j޽k��Ok����������S��oz��jߛ6x��X@?���t��E9b�3��Ҏ�������S����� 4�}�]�7��B��A��6+�&�О�[��] 4��；��c�T���ESx�
��
{����Ș�Y�l�3�Uos���w:�^@";S�k�q�쾮@�X^dK�OAt�����]7�(Μ:����C
B��ʧM���)�a�����Y� ��
b�5�j�8�	�	�SW��C���� ��Z��^�b���•�L˽��S�N��'/ĝ8s{j�	�25z�O� ��3VR�������G���@J��:ޯ/g0Z�'�4��*܍)�`�EY�`��?3��-'�k7N�66�)�z�uQqϯ��"���2���ϳ.�}�d��e**EV��	� ��t* C�W�$a7R_<�#!Z��w��l\]I�g�	a����o�@J�X�vXLt��R~����n-k�_?w��K5X�_����c��>dx!�R/�qt���%��ޢ9crc��r��������ڧ�/Zj��|��"U�g����"�m�%Wֶ?�nw���x�v_��.@T��J�?�ܟC��:����3�ţ�|�Ej�F��#d[�孏�|N1���,�v���gw�l��!�<ǀA�[�=�9m3��Q;ϙ�G�f���u���A�|m���;=wý����3`�5��`#�qO6���_r7��}()��cOm'��NO|���?���U�滥fvZ��%�1���� �Al@�  J�����t�5o��V� �˕6p:���Ѽ���!��O!V]�jN9m�� 4m5S�FE���J�/�*���̖����n?���Q.��kk̛�~ԝ�H�Z�����b_N2�^엻�"#)Ȟ��p�˷��F��>�x��	�ష����u���R�(6O?��7��+�����L��Ypv��*/gcO�O�kU'�UY�����U���2ڂG�����K
�S�b��r ~��Y��u\l�~A(5]�퐡�[]n}Z�qʒ?��
i��`RN������_��i���,��yO��.�����=Y'��9ؕ53�n+sU�^�;��p2(���Ĺ��8�q�sF@����'W�d7;�#dw;U�r��i�Ͻ�erxa>$���9@���yOy>���ߡ�݆S��h^�hx@U����dV�R��H僘V}�t���ⱖ�8Ks���E^��Ԕ,r�7�0���|�W����2��F�������|8o��*��덻"�F���I�Ĺ�P�l�,/��:��S܈z	�̒t�×���\����9�d�5z����Լ;�q3��sť ۵�����8���ŝe��D6,�������|�Pw[��T��o56���khRGr�H4�m>`nJ��G)��`����:�M�;М/lʏ(�RQʻv�@{}�4Gs�9P菇�2:�I�ͨl	㙯G(��4����z��J�j��7X��{h(gF�[C?��8���������Y���![a�%sU�Y*���ʷZvf�oL�c���m����%6]��Ļ�d_ҟ1A����l�x��
'�p��V�KŴI҂#�-�u=���'��f��R�͜�]��6�2��.�;���w��
hFH���5�2����g<}���~x��#v��t[�K���~gR~�U�}/��/>+�}W�4�Y�u�y���5��*�@?�3��P�ZcՙW�`� v#@dn٦����ZԢ���.2�:yq4D�c���2Ax����Q��7P�ag=�Χyu~.�7�a�Q��Ө�]x{S��M�۩� 1�q�+ot?�Y��c��t'-�#������k�]S��
�ͶȬ�N��Mv��s��t�n��R��p<\@^\P��
��������a��������Vk�&��ai�]�H�5���[�f����L�$�� �xb��;���B6? C�r���L�~�hG
�"PZ�<���fo�Q��2�c8�2��D�)��X�����=I��vo^����S(K�[Ăm;09�M�Tr�<*�*�T{�� �|f���&��j^_w�|HY�c�j��Z�l"$t�D���j|@��~� ���'=��r4�b�.A�!��#x��1縦�\3.�#�R"]�����?(g`F�l�w�k��+e�c���olb2�B2	��"�שB��g���B�����$�Yce��|@������,)�\��G�w�zw�X�T��8����'¾8�H�}ac��o���cL^�)��F���|檝Y��r��G�V���ņ�[W-W]kO�.u��:y|<K-7���ty�Tw����`ݟV'ơ2<v=�w��PX��������(�^��q�ޚ�Y�����lRl>s:����Hb�g]3�bsn ��p#��f\zO�N�O�eo�0SH����;H.� �z �ƎeS�E1s"��2�~��e,qi���̞7z�����9/�����W���<,b��4g�	���R��Y7������3~�ц�h?Z�%��b|�m���$�� �����B�d���Dws��ak)�p[1�Mz|�J�Xi��=F\Z��^�.�!.͇��(��gԷ7������̾+8/^�k�q�(����]�U�TZ�S�l���PK����mȼ�$h�'�g����=�`��q*^����N��d����	}�;!���A�U�8ǘ6ǰ�:SY�W�=cf�{�]8i����@ePl*&ȇ��n`�J.vC
2�m0��(�hbcc;����2�?v�%J�i�'Ԏ����Vz��x�3VVl��f��Jn;�[��w�5BQQ���Ѹ�:�t,�~Oz��}
��͘����̀}�sY@�4�Q���$ �ݣ���-�!�1��i�J0bR�^�Ɩu�!u� ��=,s yI��49�"(Ή�ZtU�뫦��"�k�������� İ�A�W���D��_���mݜ0�z�{�9�G���� ������j��gj2�����l�j(�۵��� �P����̹[�܇F[W�.ܻ
��{-]�� .��MO&2D>�5��Z_-��>ӂ�vE���	/��|��"堬�Ƈ�v3��F)E��Q�L���F� dkvr��1A_�) �������'����X��@��p��'Ov���;/�1At=�-U,tk�� p��+��.l���`�"�2Z2֥�h��$�Ǿ%�����=���=�~y�?�̙��������%Ģ��@S���ӛ���>�J̚Ԛ�{f :Y������+�DiP���W���?���AAt���̲��4�C~��C�"�湛���ư����[͉�3�t�_-����ô��~��H�_�$��l�h���20K�A�&n nV%S�{��}6�t����SPTf��<���Z��I����@t�G�H�y��DC�GȬq�jď8���*t��D3�/gfg�i%�n�,��ک�w3G%�n���|([�f���^��9K6�[)����&�F!���\�N���V~x]cq%"3� �ڦ+�H�Ո�x�:#w���B��E,�,PW`��R�����^�᭍�l�X`��S[��'0>=�����f�I�����RĆ���u_Azgٞ��$����{i�[s�7{��17?�|��"����wF�!�������8���
M�W����:So�7Dǫ_�M�&<���eC�˳��lp���X��S~������Ia
�404��|7�1�KXR��TDD����0&�"��(/�X�qQ�Wm��u�!�0�;��
�2	�h8�\�� �lm��0�ww�S08�1XL=�a}U�;�S�뇭��9+���K��+��F^�����˗�{=�:�Lj�
����oЎ��N��z�����$ō�j�;�Vi\�qJdF��"�[����
�� {���EԚ|�[�ž[�	Ӿ.�G��n��KKp��,	~% t]�Ҹ}9i��L��b$��b���m�2|�@fв�v���5ZfJ�}����T�X���u���B.�fl��5�c�3�=\êӃ$!�Ǽ:
�;��T2z�W�~��RZ���{Q���C+��HhUV�jʲ�݄h�s��׋L��W���bh}FC�V2]�I��&�؋�nĨ�o�qpP�Ɋv��%��b��P�mu��Oܙp)�IrKr��SFG�q�[>���t��������0 ��9�����e�J��[�4^�\��0�c.�Q)�hoʥ�?661t����
"���4W���?��3�z�Cxnжp��܍��Q-��_u]����4s��w���10�v��՝<����@y�e�#LW�QgΪ�u����z�J5 )�g�޹���g�*S���I>�Q�N��C_z�3t�5��8}�|f��ጧTVM��=H� [�R�\w�g��_���Bޔ���G=_ג8�E�RZ�@0~�W���&�����~��d�I"<�su��_(sų�Ӿ��w��K��`�b�H$[�N�l*T��f9�͚=K{����
:ss�5�|��8K�r9#:�Z�����y_H�H���Տ��z��6�W��QJ��/`�Aν3F�B6/��� Wj��u�'��t��
���� r�S��MB�+�J������MJ�R��d� ؓȸ�\;{V-B$L�ӳW;?�EQ1s����	~�<Qq2�lrs�����3��3�[���q�,
(�����2Kog�����e�-�ǹ���k������u����;`�ǻ[�(5�c
���D�C���]ͣ$&��
k�8�v��3�u�ϰZ;h_������t{��W��	��H��Sb��q�ga0z?^��A�s8�w�03�ڎ2���ہ1�T�*���*kP��P�
�z�48��.ј���t��*aO��[��H��-�9X4����;aЭ���,�:*�,����T�>��bY�У�GYl�����&�%�ǰ����{c��XU�ږv�9;�9���ip!.�')�֛��s]c7����8g�QU��{7㙆.i�
4q.�P�4JBWV��| S��l����Ϥ�`\��M&�n���i��%MW�7�������>�3{#<��\]�c��M�@�/z}�OҢeg��A�1z�,6�57�V?��C����q�?6��6L�+��N�'VGA�oWj!��Z*HP��S	�$b�2��o|��s�DV=f�9 wBe���8� ��ۜ�í�4&%���~������y���#�>@qډ��Πǲ@XfU�u�ស����YOAR�'å.�11�>��L���0��H�q��U�C'h/���AN��OSO��������dxM����(!�q�I3���2�F����}��=54�[y���{�j�z��C(T���B��~����w��Wed�Ӫ���e"(YA
r�U�]@���xV����6�E��i݂�P���P��B�"�@��Gg`���� .hR��� �a��{�n�|�߂�z�ޑ����◲�;��l]0�=�T(8O���$�u|��J�� .�B��,�[����W*�
�}/ۘVPQ�fmf�8��(b�=�=��I�����\����s��F[P�# z���S6����p�B���������|����dN�x�v�݌eX��J̉�C3�ě79�GG��pm;��e"�����'��[�U8U6�o�;�t=#�}������ �Q�};g4T+N��c4O_��/�:ّD0����/�-��˯6��1<���d)#���[�ck�|����"FJ���
e�3�qͳf����+�VY�Ӆ%GH��g��`�
Q�9�X�ҹ��L&w�"�;�6�P�k�M���P"�{�߽ �0W�	zٝI�|Og?ݍ��h�1��F�>p�@O�5���V�;}:��0o&������){˞�"�.�{���bj�Xe��9/���1w?B�Ez@�NЉ
6^��:�w�!YR
�ߜTf�R�e�+sSVT|3���S�1ʺ�`�nzO_?`<��΃���m6��?�E�}�5�Oz}�{z�-uW���hImV�_]�샇ȝ��ll}O��E5�9�8�g(��G~~A����	�-�(�V)`p����g�JF��{�|�q��|�������� �YUP����yj�޹��4���^�=�u��{���ի�t�[*�^����� #��eru�p����ڞ��\�B?ZY&��e�〤ܧ�t��j�v���Z�$��_��Rq�WO��ߒ �*�����0��*E�K��!��WC{Q	��HO�-hlk]�5T�2���6���x��-��zl:KvkKü&}��c���D��s���C	��F�x��GU"C��P�M�t��8�Ҋ�N0oz���C:��7�?Aw��(qp �R*�8�
��=��{��:�r� ~���n��-�N�5��B	:N5Z�n�O�x���>����
��r�V/����б/�k_�G=N�`�"	��4,>��H��)���pg�K�ᲆ�����nx�@O~��>oί�_\#q�L>{|��kWA�����J>�䅘�V=���r�۵�+8���G��H����.�D;��cJ��i�&
S��>99���WA+��a�cn�ﾢe2��3�BX��&���Ҡ��L�ׯt8��w����� n��.��oh�=ǫӘ�F�$h0V-��+���������(�B��`qYgSh�}�<�����Bۭ%z"���bX=��������d�rL�%��);++fC��������PYM0�g���Ԛ+}����U=c7|IHH`��U-�wUȄGX�>=�8/qm���p��`�����&?U��[�oH?ϝ�h�Kx����uXP�ݛ��fu�f0���/%6��a&1 �C�ۆ��wmb����=��b�۳g�XAg_>h�dP�)W���e<�@�������܇G��S�s�����l���|��ys��f�%��mu [b�^�ŉ:~��i�?�ljk%bz�
j�,�֧�o	�:�֤�O���� 3a��Q��$\M�S$�D��[iXC��7><=����Y1ݭw�hi����Ʋ-ʷ*`�A��;�?xɶ�����8�3�7� K�B��+g�b�҅n6vK�!�<Py�Er��.Z�tg=�u��l�p��(cF479�ea�i��g�|B�<�����������I8<�B ����99�2��5��]�e��.�2��~���r^2BKӨ!��9��g�}|�8_����+]Q� ��9M��"�7���<Ck��t��FS3�j�ߔ������/$��30��x`����D
���<B�Z������V��Ʀ�{N�dC~�x���lgĄ���]P¯���u�E��Z�o�
�
�9��F{.�X��3V�1�׮d��v�eDr����1Ň�Pv�*����߽|T|u6E�_�gS�T�:��bz�(N������ɻ{S����7��-
�0f��y�l\-j��#wE�{�:�G+��;e��E �+Es>����_�䉗�ǿ(P�l	� �j�*�/=7`����o��z�R��S.:�r��Ux���_��`����%�����K	�)0W�w��W�g		GJ�}L��L�I��N� ��<��sf�� �[�R����qʅy�2e�劄F&��Om���eݮEQ���u�@����O���Q_�l�)
�g_����|MDv�to/�8�_�<�A��%8OM6���� i�k{y-��o���@��Z��n�?>;t�yFA4)���;㿛�5�~fa��ipgcj��:2�R?�B�(�Q ����������<=E��6=�B���)'�/ zSS_��e���oy�L6��A��3��Mn6���xD`Jny�'��Q�/g�d)��o���\��+����b�ws�y��H?`��AS.|n0#�NL<���bF��.��U��0��KY�Y�d����&�n���;2�!�r�����0[+4�*t�
+�W���\5�?� �c@+G	�e"�@z�XS}���1bڑ�7��<�-彺<t�9[S��$HyjQo�ɗ�.�x���K�.�>�@�0�����ou�0  �VlQplՙj=X-v.s12SW�Z��!9�!dj����o-@$�����A�=���ܞ���C����nM���p�m��Vg��/ˉ�_��Lp�����!R;Y#�ts�&� ,��m��JluT��AR�]�X�����3���/�	��ζ�P�3H��PeJ�uζ�ӧ�� k�,��	T�@zeL����%�B�Fg�[}"���)5���E���ȵd�� ��tY{�������MO�{(��)��H���C�f@�>���#�/�"�
�h?���"풠�5(,4;��b���Q���?�uI0�9LI�	����rGc��Z�$ ���%�E�S��bM��������=���>2���"45A�J�#J��Z6�\c+�Z�|��^��a6�7�9�Z��߀�zh�]��W�@�O�}����e`x��N�E�,���Hn`�:��.>�ɏm��UY�[7�.e��S&�U�a
l˘q�?b~�{���5�wiy�)��Z��'6���bbM;��^�?��m�{��C��o��K`{�t���$��q���'�o�y�E�Qgi�i���>�a�b7����5_EEf<>�Sлn�=��c�xmԠs�_��xn�Bg�����m��9��Tw����d�t�#����L���o3�(���SHTKds����s��o��n2�N(t4a���y�Rg���(�DAuOϦ��ԯ�l�J(]�@�zYII�T��O�f�"���^:���'H�� �����ҟ:O)W�%��0��J�+���/�"��ᩆ?y����U�(N�L���䤵��]�Ԁ��B�Ϋ�2�QU���N�n����
�CM1�nh�yʯ@LK*%:��w�J?+>8r8;]6��+̉���
],D�+~U�aץ��Tq'(}�2��sΗ��V�����E&�/%���HQ$0��3�2�0E����Z��߹�� Χ?>=���	G�� �^9����@A��T*���<�����[i��N}�ME��������ڋ�H�+����Yq9+�������Qg��7�rP/@B��WP� �K`"�D8��}��j2�'������cx�?G(s�%]��uF�m�߁��CPV�5(���F��4����y�w��Ґ���=�%i�^�Қ?��˨��aa�u��;#�����ө�6l��k_~b��o:���N��2��Kh�8;]!.��kW���<��&K����d��ol��Y������L��ZSb�'��F�2�h�����33)c�����|C��L
�o ]}V�q��M7l�����yk���o�yV�,M��Y�M�\X�4ppĭ;����]��� �m�!��*0����Q_G���a��E"��֕�}wm�����ė�f�X�oF����u�_g.��HLJ�P� 9n&��Omy��RJB�̳��Q����A���Sg{�C��#��A}Ǚ�>M��J(�e]��{�����;N��l�\c$�]��b��c�(��?դd��
��nݣ_?�1y{M)�F�^,��ʂ��K5~Ʀ�	�!���Q��$[+�E�e��x���*��n�	��T}iiJ-A����fg��o���/�N`>Gg�=���ӳ��g,Єfn�ZO~��o�}����? ���z�Зb�+N��Zx��`6ByIYR�?�p�� �h�P�4�/g�m�EJ%�.���<S03f�k�D�OG�q��򱎈���CS��/��xa�]���s"/�;<�<��6���fe�j��#1 �S�II�+�2�9A��z@�X��/yi��4j�p����NB�\��S�D��k��*� l[�߰���Ï`�e<ut�d��{g:<� ��UX;������'.[�I�K˿`���Vg'�ԖWQ�az�=�[\L���3��ou9�n�J��}`�_[vdH�7*���qw��k_�P����IM�{#��L���B�4ہ�˓NLe%^����W�-5������:vw�r�i�yA��.���{7�M�N���~�w�o�
p]������K��P_��|���6=�����s6?,����,ޚӰd����*-c���(rFZ���U���N�����ላP�)���0��!��rCX����1�(%G���g{D�����f�fF� ���F5rbH/Y}{��fcX��j(��x9�03�\��oL�?�g�ȭ��ѹ�ա�*���>����x�ԪE %�sfֲ��|c|�Է�&����HyӈN���>�ۖ㘺Øz��i�~�b"b[@p:3k�K+ ��JT�����wQ-2m�"���g�����9��g��F�G�����V<\�;�ʊ���H����Ր��'9-&\!���8�[�Ft�U0��D�}2�I�bc_�?�%w��7������%�W��!te�����Ý�`�}Tv��@�Kee"讞-�pn���F�q�Ag*��%���T��ѻ�%�z@�nq	%-����'r+�îO����8�X��Z44��7Xc`��ŉl��\��N�{ދ]�w2>1��wW �9����&&��Cx�!*����~�m.��=R `��=\�W*�j�}�c	��22����#&	���")�Fݵ7��� �0D+�������A(�)��"�������t���E���m�9�w,��$�:���#��M��i�y�4g�� �)�x���ra=� .\n���H�brr�]��:U���^.BMr�={��LD�'���֏��~��>���ںH�=�%^?C��U羺�J�J�4��X-o���&�-a�S^�qyG�r� o��U8(9ygz����t��A�<^�o+���~ �h� )�nV�����{z
WcҲI$@\>��&P�r�ZLlxF�w�30� Nr�E0@�Q��8/��3ߨ�_U�6�P}�ʊPO�'�c�$EEl[R�IG�Ԟ��\�G �	�M�0g~������tĒ��	3�4~�]��%T\�\[[BC�SQ�<� ]K��n�)/�
���5l�hT`m�?T�@ ��>�O����q���b'� ��Zv�#n�̌_F6E�H˪�~*x��߽a
�76|����� ���ٙ��+E��0��{==�w�J���B��6uc	o�;~��Y�蓰�ܜPK�nc=eO.8�n㮝��� �j�	�g��61q���S�Q�M޴q��Mx���*�W���. q���V���,��?����xy+�#Cԭ� R�3���ƹ�&'6c����a��Ҡz9َF��,-�����[��6������3u�Q~��Ri��:آL����a�3�D`�w���-���/�es�Os.F�YM�_��`�ژVJjjʮ�;�KX���U�X�y�EYVߨ��ӧ���`��~xϷ�"NGd��r��V;V��eώyf�,?�r�����jθgE�4��60h�ihX�˟Ů�<k��QSC%6P��ڴy����T{;�#�y���J�ӧm@�L�
�P%��h#GU���@C���^���(�+��x3��x F(�|g�D�&�;4�����Ol@�ژY, ���?����3{D�����+�!!F���Cz�m�L�8R�X3�ﱈ�_�'r�K�6N�q)<�efU༢�K��Oҙ P^�˜k����N��g� q�-��7of��Q^��{1���3����huqqs{r'R��T����5Wx��Bs�[8 J	��M������ǁ��Ύ�%���gϘ�n�L���VP~���W�+���U]�;�}=fqW��Q��Z��&���(-���-��"�#d�:[Բ�PR�J��l-?�VOF����t[�"��V�qY݀��D"'s��T۳A�>q}SS8� Gd�o���a�zS��c�D��NSS�Q-QSK��M54H����h(�e����햔:�QK��[�Y���.��Iʞ�rS��HK(-.ݨ���5� +��1eG%&����IK�{:��\]�+�?{uIw)X0��$�|Vt5/osK���+M��sdFq���sע� ��e9����d5��F霼��Rū#T��U����hb�ײӦ�aiU\\���s��C���q?ƿ8���1���-����)滛"=YY��2j��y��"��j�%ݜ.�3�'�4r��� ۝<DG++��gL��\]Ӑ�{��?�x�7�A� Ô��Êv�t�;;\H]��[�^_�������\�w7�ݽ;����I�y�($�8�ˠ��ǎ���Ϙ�q>�+���&�l�:u*W�ԁɅ)�XZ�Gӊ���hb�Y��zcs0�P���G";���8;�Vդ�[��Xpw���:���"]W�9����:a��yOC[Gf 0I�p��3�ᳳ."2ȧ�:Q@���x �'����H��+��&��1W���3L�'`�J�]*jmhx��7K\m���8��ZZ&����XYv�!�g��:�,]D�������C	�\��V��('�:zD��bz�l��j\VցD�DyR-6�jxT��zd�`��,�lm}��^dhh$�k?C�Smh����S���w����/7T�YE�r{*�? �a��:������i�.��z�N�LaF�P�Hg��?XGq����mxex:��%���33��x,�{u�<�R2]qeM�r��z����Q��E�`����"Q�V��4�/_�~��?���
����g�05��o=��ػ|p~ߺj�<�`L�����a_��z��Ƶ�f,��E<�%׿&����>�_$44(ܢ��1�T)��$�Dk4�X�.x$��Еb'|98��4�L'+��ϟ�%&�����$#������#� ϒC�ߟ�Խ(�0�s�r�h��W}�I�3�R{Ȯ��j���OK<b��	�'Z1�.�n�E3������!������|aAƊZ\xCOIT�p}UC?R������o��H����(T��#�m��}�T���i�W��1Pkt�"XMc��~���ʽE_{�*du��T؇��Fk7T׊1�ǖ�L�0}�ç�~��3��b�%{��!�,��yr�$�1����Su�u�U%��v����Y�o���}������*@�!<�jP��R�=���!�;!y���`F�o��նr�f�~=]��>�Y�c%�Q�bK��K�>���.��RD�t9�k�\��{�M4ΞF��<�H~�P鏉��h��k��Ϝ�z^���U���q:*Z\yچ�z�gzh{�C�[����޺�램��� ���i��y��**�����P�Oc�!��q)�{P}��>~��q�ܢ�U	�|��C����Đ&jB����w����.M�0�I|�9��b�[� [�gOk�/N8��p�v���`"�$D���҈�X�П[�Rƌ�ש #�?mja��]�j����@%]���߭�yP�g�3|�]+c�MA�A�ꡖ����iS����`��\�ę=�w�y��؏�*�T�u�Z�����U�ɑ���k��W�=����J��[���󈐀-���m�(�2�Z�x,�r���渹K
3����7�O�s�b�'-E�Yn(��|��_�ǵ�Ja��n��ǵH�i0��kt�JM�����
s����'��8�?[���k��v^��v������;������;������;�_������5	|�a�
���;��؏�[?�~l���E��ߏ���'�~l�����c��֏�[?�~l�����c��֏��/�.{,�����+�n���h�N\=�W�	׋1�1�
��xo&P�\���<TQ&Y�q"Ź/��ގMH��R�;iy��������˿~������N��O�Z�����1fj�]�4�-�+�k���L�a��I��]���n�B��������^�+���m���BߏS��������){]З�U�|�Y����7zz��꼨��Y��=�)�Yk��?}M�jk�a��S)B����s���������tA��*
}%���t�@õ�9�񋰽�,4):3B�*J`���B��e6�A��o6�o����k�.	��D���q}�������>���o��M����.n��+��8r�[�����.�yM���|�C�?<��}�qrq ��7��/�m
}�:n���̌��o�µ���T� C���IP�١\*4�ۥ��4�b���Ŧ�h�>��p�FA�����;ڧ�//]����tH.n����Q�O���E��[4:>�/�}ʇ�����@8��M�Pl��� �4�$������U�]�y�A߬p�ɑ����B�{JEK.�߾������LE	�7%lV7'����τKF�u�߰�y�;�d���z�ף㟣�V*q��/)��I��Z$��צ����C�B�����C���!�_@5���(W��(���v�Y���\��k��Y�i%�hx�r�?���e-V��S�8lv�\^t�W֣���|�.Q���#���@Ay�?v�e���VrBo�	�������YJ����Q~ڠz+Ep���;u%����;ڿI?��B�9q�M�+��4�O�(��ۂ�d�v71�g`�9H\Rcww��t����971��ndd$�C�o��7(+)q��⳱o�I��#��!VI��v%� ��1@����=�"**� d��e��"�ww=�+�]O��@�K�8��^�.P��f9tO�f�7�:W_,j�����C*����q����PY�}ee�%���;��u��e��OPS��0�L��6t�2�!�Ԋ�	�J�eqǑj�`��������M��	fbb�8)@P�p'��\�kI�G�D�8M]��4W�7�u-���� _[��g&*�nD�Z �С�Y��X��ᒀ��9o~$@K��S�FPj�7Pm��_�H��C��\X5�+�{�5�!ǵ1ƸlA`�����̲\TM��h�m�"�g ��`%��*����b��am)Z��ԑU��h;8�-类;��B��uG�T�J�`��1�a���v(��t|���V�'wwu%�(2QQ�	8x��M�]!��G��X�!��̃�ammmVV���Co~���  ��'Z���kӔp�ySllk?ӆ�?U�#᜸�?�`�M�---=�d���eg�/FO��srh�A'�?:�0=M�*��P�]�"� �ꈟ%09���T�R��M$w�|��&����C�$p��E�V�"�˰�K�vF�Z}O(V��ZN�е_ @z��J��<���~<�팘�~wR0d|G��ˍ�I���\�X�w��f`�SR�H�4�ae6iu� `���LNFX�p)B�q��8me�������ɷ}�`àOܭ�Oc����u�;ݎ^P�+{�1r�4����x��R�e=Dˮ��~@� R�;�ӑ�Km���ߎ�y�ǓQs�+�oBrr:2c���gԔ�$=�����-�.� *��/��P��Cm�8�����B���?c3����I��$��B���� T�6k
��Xv�@�P�^M�:m-.*�HPv��}�\Hs�A�ǀR��yH�� ;� ��"PR�R;:/�z�j�#��`o��	L�MR��?��p���S,����.F�r�p "�r�ɣc�b��b��N�-�'��GZ�w�h\T:�Z-�vy���G�V@E����)�wtv2�.1�j=�zn�)�/]����W�ĸ���v/{��2�̓71�����UU���j���l&EEyD�$�=B��� Q���#ge�+P2�1���=�	���Afi�8( �p��0P��%�Rڱt�g&���Ƶ�}TO���B郻��I�'��E8 ����mc8P�:7A��^��n~��ys�m�)Z�|R�yX��sH���K �� �')U:�<L��y��0��yj �C�2����b  K�{3)rEE��9!^8�r���k
gAX���J���f{ĕ_�컀�C}F����&��*�*�Y-�l�*�hY~mHNN>��Zh���#��azT��V`*ճS�h �E��������Ǭ�0Y��� y��׸pv@���U��tP��g:�JKcc#[F����815W]�CՏ��*F��h)����g�T�$��
���Gb�:v0�p`̗��!`�\>�.@����L���[���� <fa�<OL��֦X�q�[@�ٌ��1�Ud������Gd�����Ǘ�&
8n[����EnJ��{v�6���	ǌ2T���A��3ZUV��0>��z���<� .aąs��93:
A��:�D�޻�	�7T,��Mb�\\!vh�|��)��������J�j���R�`�TY�(Dl��\��@Ԋ"�첷V��P5
B ���,.,���1(����Md�fNr/���?��9sf��yfι7�l�w������..uW�Ӛ�Q/Q�����u
�4���yw����:��r&�OS�B�:K ZG�3	LC�c��(A%#�M�T�pG�a߻�fӰ�e{$�~[J$��эw34��'��\2�/�d�OԾޢ;]UXs�x7�j'��-�8a�!�w�}�V�ߕ���?e<;D^a�\汳��> ��j��3��O��`)��}�١�|9
j`��N��)���7��9@�f���`^yY����WhlM�&P��'C�jzw�H}9����w���9(�Jm�#>��&�߹��G�-	�-n�6֖���4=Id8��f�~��c� �u�x�<sΉ<mA�:K��[?ɉV������i�R,��5&���$�DSe�YIKe��1��`��u0�qǿÔ��2�!�q~u1����n�A�xa]�%�Yi���D(3uJ(���_��16�i^,�6��v!8�'�el��$?�)�QHXN"U���DW�#��Í(S0��[wz�����ˣE��d�4��Ӣ
=���O�}R��*�}q��I�o��(T���zZ��)�7���95������w�/ 
||�c�k�J�3���b3���p������R�c�w˥�͡��wi��T�cPo�|���`�zT��vH����x�wO.��n��2�ǒ������\qy���3�W!�m� �Rh����@�]~2eTT����0_*5���nB��[˲;��(p���~� ��c�_W �E*��E��2e�W���ڰ�
)��z�ѥ��̢i����
K&�<���v���nkg�%���\�%~i���B�&&��A�y�D��TŹ��սc�"CD��[�0
B�)O��o*�}U�ݺ������2)4*J��x,&L�qGam��/8�Z�6D�oPk�=��!���<y�$(f� f*z+D�����HR.g\����m� ��<�,0hEzMލ�ք�d��x�rf��4.Z�F~�K�+��H׼�81��]a�oE�v��G6����'L����e�T��>���N&�i�5����6*���h�y��w��#�^����.q6E�Zq�_ډY�݊�y����5�&[�����`-���_Q���k���E��]�Zρj��]��={��5$�S6�d9�o8�ϝ�s��z�m�?��pn%�ХH3뚛�k�<=,��>��R�c�����
=?��DD�{�מ���2p����)��@=^�y-��>ҁ��{��3(�����
[�M��y/�K��j�;P@�"������Ԯ�\�Ө^ZX5�t��"7���V�e�ye�l���?*T`�l�D�3���.R�� '�.T�3������_PK�C�{�Z5�{�H��gKK�W�P=�/�۸�8^������%zz��I�Ĩ��]�($_���8�Z�L�$��c���J����T�[ePA�W�-n����i���m�YMt��I_�@�h荨b��҇p~�ܨS��䘥�U6l����DS��!//��I��d�T�*�z�Qcwp�p'm,���-�I	�5�F�k;���v�Ռ�u�?�ZRS6t@��+��%}K̻��3�+"㙪�S���Kz� uv����A�l2�q�בV��<��dk��z9L�Z�
'�n�R���b�4�w� 1)��rp����gz=�?IzO�f�]o޼9XS]=C�`��=���C�1��B1M���׹��5\���'_w�b]o���I~5j�t׫��P��u�\ۼM��(USv�p��p��P:���{E�w�׉�r,�78<�y���i
����Q�\��&��+��`�IB�u�hx+���_�����eb9���'�QķG��wqr?cD��Hz>%:5�`�0���ҝ{�t}U�D~��7����	�gɦf*ԸK��Hw� ������_�>gK���^3a�u3v�,p�h'�x��J�H��aN���s���������lIp����)֥�pmF�E�����$4_Y�Xߒ���Ιk�Ԗ^?�e��`5[m�$��)ƊL�"�Ҁ�����89�e�y���X`kY
_>s�����'�Η�c��}6�}b� iU"�Rm¥�Ӈ7�Z��N��}�.ni�E.����[�,;�ߍ��]��<�c9�!�Y)��8�Y����$�h������H��K�4}iU�Y��@�tॏ��Y�9/�8l�x�m2�]���Q'0��V��?�1μ�>�A�;�dȰ,��H�i�ĸ�E��^l��
d����o=^��-�x��	n�O"�������M�F�6v籃�mR����(����!�W�T-f�3㵼��bK����))����E��%دcc	Z<uh5��"��\��s�=	<.��J�������C��į�Q�L���c�!���B��jL�w�<L������X�$��5+It*�����'��LU��� �P�4�P��T�"��������q��I��h�8ހ��c�C?Ț8P�
�$b�2���<�V��S:8z�'�u�H�l�_X�o_�4���?Y���{��s��7�gXֿ�b���{YE���߮NO[Z}��__��u��k�������W�t��/�}~�r=�.�L�c�qo+?�*è�Vm�ќ"���Qmc���_+@V���]O�
7��}���i��ɓ'�$�i�:EfO�BG�y5'�[���wg�tΘ8~�b�=.ەi�~X�g
�K�a<��d���p����P��WۮA��3���jhd[�#t��-;������{�"��[_<��\~��օ*eKa>�$�$"�G�)NH(8<?M�H>����4�./��H=���7���t�yc�#!hU�i�����[�N4?�w��؅n'zӷ��v�-;Ў�AP�w=7�KGy�)�����x����H.WhAƪ�(~����F	b�ɅB��O�#J^Ң�$���P��A�nQ�-�����"��ϧ۴���~���7�\S�Qk���ؒ��F[H�O�[�`w��fO��zG{ޥa�)�l|��Q�l5�竅D4�"
�{��ʤ��?p��W�,Y�`�<��1����\nQc�!ˍ�z57��-Mt�_O|w��rc�Н����"�kɳ8��������(T�⤶ƢQ?O�٤1[�}1��9b������L�|����������}~V���Jr��+[����-Q�J�vg%:i�#1cTQw1F����0��� gWȒ�---}iJB�_�mHN6fv>���gXT�co�=٩BgM�=�Bg������Z��l�AvM�y�ۤVG��p�� 2��w�L)'�b!q��J9�� /�]�h �y��
�z˥�ÞQg�ImO�Ԭ*QC��}:O�(A�+0��������M�J�f.�!L����O�0�ߝ�ȑ����*<����AuuujP�9X�^ÞQ�Gb=���h4����>cSJoa�S�2���B�z˪"�������lkW���6(�V��0�w�z�č|�ԙ�o�O':��)b6���8�F���-8L$��6ZV��SF��@Ss؇;d�>|�pgHȈ^�*��3��*���ǎ��Jf�������J���s">��(l�Bh��_�t���C��)$x�Q/�^7٤��m{�YfW����:v�<��==B؈���|�Z��|�L��,-3�B�p]DP.*�kw;���s �MzxyQ7�Т�Q(�F^�d�����k&�=�e���\[�����k���]ޕP��N��W�������G�[����j��A���+E��|���~X�@��8���L7�����ۥ0b�
��w����"Cm�w7T�I|~I��gݻ�Oij�Dyo�E��?�5�)�h>��kd2�������i�iɻ�H�xy�����s��
GmqQ�o@ na��� �L���_��u\xO��ΓJ,���y�u_����5f:��5nٝ�b��'!B�Pa4Al[CA [�s�l��GfĮR>j��(�0S�]͊E��ڥ >1-
�יe
�?5�w�fGp�ߨgv�It�%�,Up�����B#-�<t��s��?>o�w2g�H��82�/��v�^�E�Hff��$uá�D!O�R
٨�#���dN�	�yCh���a�}����F��J�1�F���y��Z�p��I�����W��[���۲��݇��B2�<#P�w���O���ų^!�v5F	��)�1���ʸĜ��ڀ��;�Mir�Z<1����������s��c����ξ��J���<(z�B��)M�1d�k��u��������I�tY��޼��?��#�>&�`^��"�����+dwhF��{�5(�-���P��{ o�II�ƶb� n�N�-�R7�����N�vVjʶ3P��L�(�Rw7B�@��G,�R��J��T�vR^ug���ѣ� ٜ��Go�Ȣ�޻w�Y�;��MwJ��4�b���No-O�wk�S�G�9����9�L�:/
s!���w�.�~Se�hNg~�)>�ȂL|�Ν;��z�6
�)��%��f5OA�S'7>��QFB�E���4.��aN�?q��?7��tM=� ����V/�	z��"~n~Zk
E0���@��R��F�w(Jk�����J�MP������)%S���i_�Oi#�`��	�2<��n��^���0ϙK_î/��zK�WG�2)
��C�ū#oƐ2G���3�����������\!�+A��S�%'��L).�ް�s[��nS:2<8:[�3�Lff �0�ܲ�����F�w83�u ܘ�%����Bn��u���Nl�
6Q*�I�n�r�װ��ԝ^�P��bD�R��?��s����� �`��@8|�[���(�LE֯3CGG��sFW��8��fܺ�Z1��}�@]� bX���G�{	s����2����K�9�(��F���{z��$x9�A�6�T��+n^�}���g4��9�k���Z	6�:���DR����{�i�&�,�Ǯ������|f�)�������J��k���v������hcJ/� ����:@ �qM6��" (Fg�X�{x=�ŏX�v9��
�b?S��� �L���H6�a2A@�,�&�b#��
)kZ���!r:�9���l^���j����H�#�Ϗ��n*�P�u�'��J&gj�������^	[C]��X ��|��<U&����D\s6���~M�dB���#�}ɑ%eն���4�6%Z��0џ)MR�?/��[E�*��O@/�k|�%��s)LW&)�Zka�ZY��j(�] �;qK�?G�l�k�!cѫ_���5���<�q5�)s���d�\��=��-�1��]MԼ��Q��\}�5x����P�&�υ�VO|�_N.��_'1�'?���X��iS~Dx�tt�b>� ����Eɕ-C��1JO}ww���aP�5Bé.]��z��l;;b��n`샱�7�֧��G=#�����A�Uٙ�oĝ��G�'&֢L|����Os��*�W��v[�:S[?���N݁����v54\�)T��ׄ)�������BC�@�����b�0����=SA��h/D��Ľ��Ə+�M�i���9����[&v��}x�#ۈ�ϙ/4�(hx!� GK�^�,��m��0�.��OtvvN�b�/�8%����]��,Gi������@_^�v"��555�j�N&%K�%_�O�$j����qI�R۞��Vc��d.��R�;(��i&%	�o���q��IwB43�Y-��MgFa	�g����N�9�	���$�a��
�F6sU�=�SZ�Ty�=���<�p�I~i�o{�n~"��P"JKk�t�`�EI�C����Z?��� _���?F����@F|��-��"�\'��%m����9��ߺu+��0��oi
�6B��_M�I $������3�~
A|rg�7mU�1~�����0\��$	�n�on��s���7 �����f�
ןFk�0��RB�pB-�٘āOıwRO	��P��%�%Vp���ɆҨ��ɅR��Br�^K�Fs���-�w׎�wS�;��-���4�73��)n�LOq�KS|�mo��#��"��%$aL�1>/J��k�����z䓡[G'����y���3�/����h���_-n�ĴM�9�52"�+�/���e�i�0G}[Pw���5iiD5v�(����p�h;G�4�o��rVH^Ւ�$X𲡸4!9��S�����i?�J>�`%�x�L\�:u���qS-Ε���m����>l�����Z�Qw2�����Y�a�"}��2Hm)��n_��If�C>m|-N @�! ��Yi�1o�[3)'���6�Ό���H�풉C��bn��(�S�l�6��ajL?�dS���s)9�m|�Mu�|��w�K;pQ,'I�=�ԩ!c܀���x���+[b�힦E k�@��Χ*�"�N�����3�� ls�dq~�o�U"�v<���z����e��L[u)��
�4骵�:�;sq�VNS���ýGz�e`��uF+;R��?inn����÷�l��M���JNA�i��Q����?��>5�y	?0Ց9,5���լc��fz���WEE�qS]����:�+��Bф��&YB��q��PU{�{�^o&k/���.�l	�͊��y���\�5#�$#h���a�?B���'��&�����Cjb���s
��7�=䌨�A"
 B�E[�Rq���l�N(�Ĕ�B�dh���S/<�Gaů��v�&�&p�t��"��N����fH/��	�R��g��<c��1��0DކA�̉��c�|�8����Y;8�ػw�I�w��Wf���5P!b�f�۽�L�V���B>o�O �lV��.�{kJUn�SL��>�C(8�@K�M����K枕h��-C���XE褛?�9k--[������b'��L YO����|K�р�C;%��$���$`�v5嚸z8u�A�Mm��{���=�nu�'�D�&%>`���J�����ԏ�;*��|Α�,6�$H��S4��{4iۤV[���	pxlY����|�xj�K���+��3ձ�W|�x����d+��r�gX��ˆ��a���/l�F���|�B���#�P�Bv}�p�����-O���[Ba�*;��0`��=���7�ŷRU�z�z��I��s
�W~:6yv��[0kͣr[��6�-9"o�0�z���:��G#���T[B�*��#�SZ>Y����s���K�b&�춃�Ozc�C?��N�h�pܫ��0rēA��a���6~ˌ�r�Ġ�;��GIc�4��Rq$��#B	z�K�J�^����
�d^�d��ifl��d�L=��tBXۨ����ͭҁ��Q	q� �J�u�]�B�kN����,rP��[�����I�O�h���M��`��/ ^>���֒0=H�bQ*p�]�-x�f�,�+�®F����dj�D��3�v������π�+��Y�=�{�����D�3=�5��B&�\Q�	�>��$ޮd�O�J2�b��iK�o�,�N��e�}�W�)7W���g����)��׵���kB�4f�x���.���$'_��Ѳ�^�{um�y}�:�J���F�P=hM/*�CS�S�|}��1,��+��m�"Ɂl�×�@�mL1@[&xI�I:O��n{zE�Y}C]�9��j�������li�7/؈�?a��[��=X��G�)t�*����#$J>�"��/هz�C�����.y���7�=]�3�ض�\i�W߫B:Ŷ� 5��8�oyb�l�7T6YY�[#��_Lɲ�wa���1#��~�z4��#k�/�B�%�Λ������P@�`:��sێ���9�U�h-��
�f*��s���PX�Z?��P����ɌMh��$�K.�����'��bz�zrO0/ �]�vͮ�g8H���b-�#h�˩�P<�dسK7w/���J���U��!���+kb?���\�$"h�h
)�.{��9_�^8��K����9w�x}�����O���̓�-�P�7��}Y6��V�6��7�~��w�p��`�Q�<9��IĤ��$�PW~��ݯ
�g�G�>���H�ܑ�hg
~�+�k��2�&���[�6��_a�ap��S[':n|>�M�-oFۙ��"Uf	j�WB�8�cJ�L����kZ3��1��A2�2�s�W� �� 6�z�fiE�͉��e��,�#_a����Ȏh4�N����ѣ��e�T���%�=�0�ҕzK�4,V��N���)�b+��D�W>^�ũ	ƪ����xH��	
n,���xw&Q��l�B�F#��^���-P�O��oM��.�+�ܕi�.R�I؃�t�;�%�$Bu�����YR�^�2�О���@wz���!��<{�<v��t������.n
��G
��^r��cK�ÅE0-�	����Q��Q���i_vm�\��0z<�����9��&`�{Xe/SSSup�u��XA�%�ʕ.{4��e�)���eo�ī2���{�ؾ�e=D���)�	M�zܡl�[U�.ǀ	^=�T�|� �eS
�s�@��	�1�N��ìq�:��-Abc�z#�jv�������y~E;!�_Dl�S'a__��WS]=U���\������hkkc�Ǒ����d�Fë�]�H�+��>|X�Qei�0�����M�Q #S,�m�YV�n�,��Fq�[�O�5ڃ-�k��zȩ���y���^��:Z[@��wߔ/_�ͫ��O�շQ�c�ՓwI�yC�ȼB>#�w�<�传�w��)j�ͻ-����\���u��B���������P��W���R��F���?��7Ae�h�����%}p�ZM�Pi�Sւa���k8, ��z��*K���Hl�-1F����Ta������*���-`�y�M�x���vÅ����n�\y�'�ƿ�fa?^�~����]=��d*���rb�k&8�W2܁>gsK�L�y(&ѩ0��6����x�O^���d�t@�s<���1�5BuY��E�q)�k��=d�z�F(0�:
�I���@'?逦��9qѣW����y��m�+�H��)�,f�6	fv�S�Q��ᐢ�G���;�r���[4(^����I��9N�3|���f�1���+�1^l��[�W_U����vZ��-.NW�{%Wzi-k��+����J�&W�������w�)}{c���7_ٝ]�W��{��O|��-��EM����}�hZ[�Z�� ��s����t�\.׮�[2ͤ��s�{kϑ�iji��`�\B��#��o^Q�W�/W��)��y�!�(��H�F�Pb��MK7g/�	�/�a�pϓ'Oҁ�����ȣ!r��h����;{P}���ȘD��s����p���	}�;SzX�M6)n���É�NY$0�Rm�b�w�K��U.�.�����e���?c�|P͔�Xwi``������e�
bŃ��-�Z����@)�Ng�2���:����x"f���h�$�Ň(�k���ů�n�['�����Ǐ��kɄ�+T3�&A�>'�"}�`�̾�q�
3��2J9�s�]���cW4O�O�n��_��;��e"�gZw%i���Dۈ����I�j��"�Gݻܐ�esYD�K��| R�%�vQ�����Oâ���l��}7��?��G��O�v"� ���2�HF���ħnj��r�Dۇ�Qq�8�b����O3���;���԰%���,����LOK3��e���a����m�ήtw�qLF��2����C^O2)9H��y:>�p�L��dq;Հ��,�K��ˏ
�m�%!�+CE���)�\l���7�K�d���%IhMJ��2��$nn��+/�t�nS�D�	��}��>*�VBIfWc�m��B�y�l�}��~�ŒU��V�/V3�S�-���� F,'��+z�KK&F�B�m�<R�dxܺ'��(��"lD�o�*�qb|���
���hk��0�]��Y��`K��ml�#��Oe�L ��Ni� 2��/���ܼ��ſS�L���Ȇ��
���6�5�N�!kS������r[�*Q'�t���Z{?�5��R�{Xx�I~n>��gI�U���s�2t+�q�J�}n��Lt%F�P迣�1t����-+%����<�y��$x��0i���GK��a�l�_���WX�S�Mg[�`���i�]nJ�Y+ Ch%gѻ�D���C�&n��m��^.7������G�Oa`�[H�χ��vNR7��So�g�����*�l�ӣu��q/�̸� #�Y��{� �ߡ�7��ٴ��,�Ƒ�
gt�o@w�
&,Iu1�w���l��nZ�2_��A�"�!�|�:|>�FZ�IO��Z�~�?N��`�D�5֎�9�k1[��(*�>��/u��z�@+����Q���n}�h���Vd/ɢ�un�S�+����]E�q��k��a�k����bE-c�>L�:���t5;�:���^�w��<O�+�% ��Vd�c��7#}Q���R�Q5���o�BI�s�͔�!�v��ck"�1�-�v�q̬lɟ)���U��)�8�t���Üv�.��	~���s�4�[(����Ȳ;��t`DV֤�NMN1`�Og� gvF)=5UmW��)�՘��v����}w�Kj�
�x�tt<�r���Vt��	�Tb�&)su�<���D{���K�F0�"/)9�|^�	��2�f"��b��K�y�F��~|�~Qs��3tJw�z2�1E"Ga�V�/:J��PJd!�'��#E,��hG��!�~�Q�;������ %=8��\�%����*��VI�WVV��e�b*&	���շzJ�qK���Gijj.?�@�M��UM�mj�T\�d�[6�@���u3��"B�ڤ��)))I�J���%�Pe����=��:�g:�%x��w�����
�������ȓ(#���p���%
/5V����B�ק�R<y�^:
x�^�^���I�m�=[F]���֚{�3�	h��Sj
�.�*����)�0�XZB�;:��W��;���FԞj��6Z�6�|�}A�É��e��>�a�ǁ�����c�y�6�r{�n�ڥ-�)MR�E�C7��bF렶�𒪓�No�7^P��_�9#�!�~������Os}Z�k��v�� ����_�񸮮�!đ(/�o��Rw���WD�\G �����(�{�����[f�~/��^i�Mu-MMW���朲޲j��c�)�i� ���N>/����m��U��f�1�'�$j�K�4q�*c��`��-{�9I�I��ʀ R��O�}*�����KU�լ�lY���D�~OX�㟢�x�,--���s���~�U�kA��L�7C
��c{m�i~�w��Cn!)r	�8��gϞe��>����b9��r�,�Zc�Q�̶�/�Z�������﬑XV	3Y;��ބ\`�)�iRRC,x��S�w�1If�P Ly�3| ����@n/������xe���)�>���ݭ�]Ky��ƺ�ӧ�Y vz�W���
	9A�P#�A�Ѓ9@��{h���-tڱ��}�,����&n�ٚ�zrp1�����z_Z�U%R����I�ۏI<����]���LN�eItU�1;����ӧ7/@���%�I�}Nh&����hIͰ�*���?�5O\`h;�	�6����>��C���_p����H����*=���Oڢ�=\h5�x��	�?�*Lw�J���A����"�ҳ��һ��W�T�tu��s��/�<�����7�dK��d^����x��{�t�$�^J)Z��"2eK���Iyâv���T��G�����w�"��
ɥp�r DiG%[x���	��O�~*�％��qhѐ�~�wL#I&6�I��D��H�֯�Z��^����+>��wEid��̖���u��o�V_I�Ç�u-��'��.x�J\�?$3m$'�c#��W ����=�'3����99����t���PM�s�|�l$��͆-il�0�r/̖�ʲ*��yVs7"��^��4����YjH���8 ��!KEa�P�g>/��oP/�QeQ��+�}*���k#兑�,�����[�v3�m��r�����z��t���ׯ-�΢_�=�)�*9�>ګA�y��U����2���R�S�̄R�6�Bq��/q�94�ï�,�����2�ZEC�1,�ܧ�*�RgSJ�EaN!�W9�=i_�H@��tG�ֻ%Le����J�`o?��h9QJ�`N	�i^ҝ�J�s'�x��63���>v�סd����GF���'KD!EN1��:A�9e�e,-X�vr'��`�yqwh���N��tzN��v��1G�+Q'6H�Z��\ûh�ik}]�������*�Ϋ�o�B�v�B��sꀗ%L��I�\h�*���ak��Xc� J-̮�dM@�*�}��N�^e|�d�Z-,,d�_�Η,�0��:Ρ�	u����T�U�,�ws\���Ȩ���5>�D�Ә&D%ǒ(Y���dVٵs���wĹ���)
-"ϓ��Y	&�jw��@�>��Py��%$��]�~ɕ-A��݌�ɆHo�����.ج�!�zD�����Ѕ����{}p�y��ڝX��N7�����5����<�/٩G�M��dD�K�������/�|a=x�z>,A��l����g2י���ٳb��-��lTH���SKK�#�J�frV��\[H�D��MU�!i��nj��>[>�LM��Ԇ*�Ϲ*[��|�ߊ����{�����0_J��/����T[ufƆy�� \���3L`G�a�o��)Yr�oPt�`��=�r,0��ݳX��%g0.8>�}(�����n���z9/99M(L2)!��rU}yP��+�.i3f%'xI�T@�ܷ�0xP:K9L��9���ٵ�2�S��䔴rGw���*�cդiH.�>���~�.* ��H�FtI�����p�KLyN2p>'t�C�tl��j����z���NU��ʽk���G:�y�ƭd�B��K�C�� +}e�Q~FqbL\�]J��Y=�)���uq��9���4���eW=QDV2��jM۬-���cc���I�3�5	C���Y��S����ROi�Ye���ߌD�1���H��}"u�8���<�L�*)'3��(������ u��������ڎ�`�r��kkk��� �J�~�Q�qdA�x-�ɰ��:��n!MT܁c���������wB}�k�)Bs"�͂���^����ID�$Ok\�l^R�&;@���Ν5`�	�RR/����ͫ�F@Ѥ)��Iy�~e��*��%���3lQ�ѴvW�''�g57c{��)�7���83q-�l0�Q��F3�ڇ����Oi��p婴����swϴ���d�>/��Z��ݘ��ԡ#�1/�r`W��:2�:��ws�-�����Ɇ��X����[�D�Z��*�0����y�Gp�+�4��$=�)���~�����$B�3�eH�B������0Ԝ�M��B��k2�$�g�^fW!�Q�	>S��m���W�W� ��$>������>hb(O0�T%��%��=�3�����Ɛ�hC]Yh`�������4�)��|���m��Ii����E���yk��U���Y��H���=<ğ������yb��B�B�y�-�B�ZF��O~V��Q������*!'�w�} Q��	ޑ�1w��jFX3ԙ�İ�eG>��χ����C>ݝ	�E7�zDT�u��3[�H�b>R�
��1w�¶?Z�n���#��C��v���N^#���X�pA����:{�厴��6.IB��$:����<�L�Z6�'��i\B�K�JB]�,�jL�8|N56�@A���Ax����=��s݇��cS���k;��6YY��Z ��������0-Z�og��Cq7��k�Uq(�W�nT2f���۽���̮,����6�m؝�F�r�=�T���aNJlݟ�`H5��*�s�y��h(�F�Q���PP@����C?��MOi�۾����u���f�c[Yf.�5�A������G��<�~��߹��(��Ogs�sds555��Si4����M��i"��6)M��(����? a��0�lo����vt����|`6-�R����*TT��,h��C�v@��1�Iku&w�|�ip((�&��)t0��$�k�%���la�k�Î��K�2�W{�)&R=|e.xρc�e#�===��(k��u��o^(������tP����g||�?�kqT�}ܒ��m��Vp�����TQ�T_''�+g5�[�3Y�{����E�_�*cRr�&����%�r�ȧւ�I�p:���\��x?��Ǘ���u��yG��)~�牀y��<z,7��]W�����5"}|W���ں�-��*��[8�����5�3¿�;A1j<�ѱ��E����i>��k�tP�!�ʀ�.���Ӷ����������	M�
1ëX_��ЗDlkC�V�rZkQ����D���'���ebL_����7_oY5��܆���4��4<���� �Y��s:���]�K������k��o�U�Yv4B��ni��յ�1ޯs9�)%31<6b��&�.A�}�%i4����W�2M�NF��P��台�X�l�jV%<`�Ѡ?���<��s�Zn���������~�� ]�{1��hZjj�Ld:�٢��-!�����������|��BE2����3Sa:�!�z�z8�³5�E,��+l:���#H=:�IkzVe�福��x
���$Q�r|55�;��
�Hm�x�q���K��k̝�?GL�f��>w)?��95c٢E�9-�^6/BM}���e��w�Io��~~>��\M���KC\�٧n��8�=����e#������"��y�17 ?�_�~���5{y0p�'�4��q4$P�8�T�ꄃ�z�S�>���_C�p�t���t�UL�M<�3�Y�����.7�sFX_��liiI:1vj�P�`i�wb�1��<��kZ��C�w�eU��R|�Ӈnc�<A7�%>y�)��n�XOybH�����;+�j ��!��VA�jYN�����'>�\�s����Pt�c�6Ӣ�Xȷ��w{�\(�/�c\;(c������ҒٕZ,��;�[�0��G�%��D����OvgگǗw��*�~�)��p�_��[�C��*@&4��ݧ�A'�sbbb����k�ل�ߣ�`��i�.BhD|��h���#,�Ǝp�ִxO277_>�e��EY�#kO�������M��u�bSB&6�'#���R���TIg,[�Ty��ah|g?�2��HGG|�_�	���R|������ii�Ȳu8��昁ǂ��d5�8a/��!��8vj\�f�(l\mB/\��D�pb h��}�FwH�0��i���I������,�i�6!'�=_6dj^9��>D��YNn��<IO�P�@�d�ڬv쀎P3f��w�(p��jw��V���� �GֶۓN�8��Z��
�N�;��sxJ��'k%���C!k
�iI<�ÿ8��
8�n�R��ͫ��w���&%����%�˿7A�Pv�14�����/�{����IY�m[��U:�z�����7���w1Wk�¬�*,v�W�ε́g�.T8F}}�3%�~�u�p�x�������C���Z�̼��;�����㠾�Gy�95����/;��[��������~�e�n]@��4�j�������/�yٵ����y��w�ZeK�6��UP�?t�/޾;�MD"m�0'Z�~�e����T}����.�Y�Ź`kF)Xm��m��i]��+&q@��9�e'h+������u���RO�0��u��.W,`�^4z7fgg�U��U�h�=���7>�	�`%>�d�ȝ��3Fq3�M��Í��N��6�1�*������hS��-�;=.B��;�ᒖ���{��~�Ȱ���3��Uf�q�ƫ�� ���`�4%	���]����3)QB9U3�����E��U�����/��̄2�	K�k^�����J�^v��4v-`�h�U*��^i���������ސ��O�mS�7i���Zң2�!�ʀ�>�h6��XD����6��a=�m[�M��+��o�{��jq6�d�͓~���A�f�k���\Xi�3p�!����ͻ#lZ;w�nu_?y��4G��t��X���F��3�.=۟}���V�����������*��*S_%�N#�}�����b�椇�!b�:>X$�]n��BՋ]���O��j��Q�K��c�M�zt0�T�l$Ҧ5��u�[���6f���G���ܒg�yq~SOK����.J�����z�P�F�rS��G_Jtj���`�d�����=@�0��wcn�8����`�����������?�e������%��x�J�q}�����\�2���k�x5�����=zT	�vqfu:*e0���U�Ɛ�������$�V�msO���	'q��1�L�Y��q��98�σ�jD����.�\�>m]�N(�+JF� �ռ�|�&5�w�ɘ��$O $Xp�tA��]�9�y	�(}7��t���eqkC٬B�e��i;��;�f����O���'pDy���=�ڷz{{�U�8�1+�· |d�`Ct
;�OdV7��"D���\z��Q�"ufgq��8�;�sW����{%��;AxYz�n�D�hl'��lݠ|~vC�U�7*�N�]��a�>�	***�?;����^���8�C�|���q���� zm���D�pH�\ߣ���.u�Cv諎��`ȓ�ޏ!3�޸�C׼��@��^oe��W1��(�,�ruu���ه./{u�$rF�H�(��A�p�?2�ќa�xJ��$"D�X\��S�|E䩈�w��[���骯rA����}��T����	c���.g5'\���ާ��
MTO7���G��S{�1����<|�O�l����
Kޫ�k�%QWQ��?������z��6_���6Z��f����^Wm�.��ϸ$�0�W�W0�L��,����2��U��M7 ���0���ᶝ���(������#�~c���w#��N-��t�B)��>zl��ߦdV+|�	 �i,�f<8���16���in�4@�ر�o�x?�95���-�	�f��9F�o������r�����94�O����<Y��x���O���-2�s�DdeR�n~j3����3�gc������4�䬉z��I�Y�ٍ���+ �TU&�s�H�=�L�\k��C-�u	(ƻ�g׬vB֮�>����O^UrH����ga;����G!��5K�S���Ts\����ɘ�\:j|>{U	�����o��i���'�]7p�X����x1��}��DoFd6>�"�:��Ym��c��gli=�dA7zbSp�~b�@�?�[����#��A#l��;�c�)
����xP��7����������z�֟#��h��	�:8�zn�����D� зy1�{�ٯp#g,��G�ؙ5����>���,��������ɘq����5�\n���s?K�V����$�1�7�YѰ�	x��`Z���s`\~�J��
~��e��_<ϊ�P�pD��L��^���7:�}6�Ψ�ǐ2\koCX�G��3��q�)��<H�S�F�ӈ"�0�K���K�
g�F~�k��~AO��?�Ҍ��3	q�Ol�I�9&�E��zzf,�1ow������Tvz���|�Ljc_�ZQ�Uy��1B�y ��Ŗ����/�G�u�� -�<�ƿ���
�h�$hث�G�Z�p$��{F���f߂�۪���-��?�G �+[R4�ŀ�u�vw���
Cz��J����Z�|M�����6sA�����1��c8�~�ͬv�$��,�d�1�:�N��Ł�݉՟� ��Km�n�<���  �MA�jL(��:�kٯ3�`Q�}�$豵U�t0�rf!��g]��hn�]���e�^^�k0Fi��}�km|jf�23ҟ�R���FC=��3�V-C�+R"2@�� b�Y�����j��]}8n=����ZSX�k��[�� <�-^�������C�;�7��hGe������2t4vJ�{�l͂�-E�:%���ڬ�˙��� �܋�˔�}J��.����?u�do�������K�@9g�����c[
wuqY��Đ�y~}�������p��Q�;��g�%��w2+>�����ID����&m�?��\q������\2�?�e?����ask�����7}�q|���wà��N��C�l��683����C�cf��R;�p��~�
%ج��+*b*�Иd&[���{�p������|ļ��`�TYc�}����/[veuM���`?��K��s�7�﷏�.8��ӳ!"ݣ�C�ZV�Ǔ�R5P�߯�C��׎��rvn���}9�.��xJ�ec��
�֔�ŀ�]�n��P
��ql�Ū�� /w#^%6)h߅���fm�;+�,�� 1c죌ǻ�Cٯ�A&����g?����@��6_��v�7��vt.���k�y-���L$���%	Z�;�4�/=�(=���^�j:S�I\phX�}%���%��5��r�~��� PK   ��!Ya6֌1!  ,!  /   images/a0acbd77-339e-480e-a1f6-37906f79b183.png,!�މPNG

   IHDR   d   o   %e�   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<   �IDATx��]	�Tչ�{��Y�f�a�T�EE|FMH���R&1��K%�HʧyO�T��h��*EbYVi�b^�DcD&B�HPD�f���Yz���N��s�N�L��ՙ{���]��|�rι��������͕(�r�ɫ�x|��瓕+Wʩ}oס�%ǟ�G�7��{;e����$�0�< �L�= ��yR�7��Y��;@8u7���H$��P��q�R|V�O�Q
��9b(=(a�H�x<ݽ�ݡ@ �u ��:@�9ґa(�
�����x	�����'�q=T9����|V�R�D�NG�@�]�-c��=�m(﮼��]w>�P4����q�^�
O<�):ztb����x>��/�דP
쪜C�&@�,ǩ��S�������*+wu�{����rl�鮨\W���'�)���_�ŋ�{zz�}� � �f���M*?�@F���,|��(��F��\��� )`�,@
P	f>,ӟzJbEE�Q]-��+-ӦI���> ��f��y
Ǿ���r�% �aP�'r�իW��<S�LQ&�¿��`�=*�x��={$��)	��0���?����wr��(������sᘄ�/��^)߽[*P)�JJ�m�d�h�l�`:J��"��6�|����x@�&6%� ��
J���
@�{ <<��:�
d̃�B�D��dg�$�Y���c�"�o1ţ���0�z���۶���ۥ&l5�� ������r�ziA���h�	������q�����㥨�(�+���D�yn:"�8��J2�R@�@��~�0�pK�O�}�t�'�zbN  �*.�� ��8V���A�������8}z�����e)���}���ݻW�;��bI�3J���4�6���믗�S�JAA��"T6�l�N�y�u�������G}�Hh�/��+.�@y�++%��1B��̋���k��@�#z�A	Q($��"1lc0�Be�8/������JT�ڼE4X����g���r��˥�F����ƃ����˦M�d͚5�}eӱ�A���E���o��x��DP��bj���	<D��D���0|q��������T~5J�&M�bT���Z	"��������	�9m��8'�mj�n�����K7|F���Y&�i�p,�PL��bM��i��"9t�5҃J�FS�������Z����U�V�\w �Y�fɊ+�£��{��~<k�S6��۪-[dܳ�J	Y�02��'�c
`��P�fΔB�Gj�b	�O��[[%����J���A!�hT�"��% w�g>#q������7���7�g�~�߫��X�pנ��׿�l�.9�t��Ι#oG?�+��?#�ZT�o}�[�_�B����H 7��/|A�n_�B�4C�mw��!G1��c���aFj�n�8�"�s�̠I"��2� �H�ĉ��&� 	P=�k��Q@���v��1�0[�¹�EPP	��X<c
nݰA��<1<�Ɨ�Gl�(��g��N~�1)Ӟsw~���i�'�9p��hY&��K�,�?��OC��Γ	�U�IyCh���ꤶM�r�u-&JF���&3R�
ʌCɁ�*u�%
� 3��8~%�y�
^����T)�B@X���E�sK'p��������u���%�}Ø�u�I��Ș�e��Y��C��f̘�*s]]]����%x�k�J'}�P !�nv�&HtP#�T?�|�� ��?�Q�':�����qC��Rs��2r�B	�M���� (4M
a !+�H.se"��ɲ�P,!�ǖAA�!0>���/}IF~����5����1>+.3F߂s����o��96���;�#���z�r��@��*G`�H���� eeeif�f�W^Q`��7�t���������Ȇ���Y��*b��ϟ/c�C�)FA=0I	�.��ёc�a3� h@�
{Sb�aLb���k����jP0d)K`j�|�W^)��WK�K/)T@a�������P���xZ�L�o<�����@�*S��8V�l��U�>÷'�|RE_��F)�Rk�t�,y���f�Y�o�Y�L�`��8OϾ}��ͫB0X����f�E�ñ١�����2@���k !K,0T),�����&~��R6z���;�cL%[��OE�ݔb�wxJ/�ɱ��U�'[� 6;MmCۊ(gpj�dD��N��6S�(�_,5pd5���D����D��###;4,1� (���S�/+��8���g?�C�>*��/��:�T�%�z�a{�0���e���g�GEs�sn\d4Eنj1������ �b�ɇ���
�!�^
m6s���Ҿ�1Y��a�*������5@	���53�� ��^���J`�0������?��Y�0�_tޢM�w
���5(��L!r�� aSGKK��_��Y�D�`�;�DEP��jo�A������A��1��3 �!
̈́4 �
D&�LJ*8 k��0@f �����ϧ�������_�J��+�o���@!S��\kp�C�)�"9Bԅ�����h��M0b�ႚ���% �z���lA0,@h�S���>&1��<z�P��v8�X����sΑ�?��|�$����yMҔa�C��i�9s4���Z5o�(�
 v��Z`�-0�l�!��2;��V`�T�!p��_��$%#��-�i�x_�4se�a�B>V$�6�s�]wɞ��\�`�(ԅ�)l��	��  �͔%@�=zԤ�@)�I������Id�joc��ب_�� +L>�I��I����n�AVv���i%�)&���S���w!�0�ˀ����{8�n�J~?�@�$���e[�!n44f�L��:��{��`;� +R�i8��7�f�>3LK�1Ae���n�0�h�i8e�E��*�����À��ն����Su"%�`�F�.]�jx��I� �>ÎtN�=+F�~#v�a �|��[YF_���1�?:�:U:���T`��=�ʴٳ�� mq��ȼ8���:��R7�&�-7;�I�"1��o-��=�ܓ�X���}5�׬�= E��{ǳ'��Z5�� �A�b�aø��.�bd�t�QG@�i�t���������a�n�)C�Q�b�|�!�5)?":C�S/@PD�&|ٻ�R�g�Tm�.�C$�:t���iӤjʔ$3p!��� �-)��AӰ@7�Ь�B2�	��U�Ρ���i��i@<�wF�2�C!�
m���oTϝ�@�����`Qy@I�{��A0��-�o�E��_7�Wq,��(t���K��t���gĭR0��{�ĕ�:��0�����c3�C�,��4��T��}��ej �bt��ˠ_�x}��� �zjJܪG���7PSJ�����^�r2�>�È�g�b3��Y��,��eiU,\(m0[�d���8߀��]_F��c�� ���Y���W�c����b��O�X��`{���
[�mf�u�K��F"C{�M���;ɨ�?�>��4��$ฬ�lӥ �'R{��Yx���N�bE�r�p����C��g���5`hf0o��~�aE�'K�WH���+o;J${��(�9��JE�,lkKb"�B>߅ �괦t��	�&L�HC�rV�u�q�-��3�����l��!)T���8��c�j�q!N�%�#/HN���f��
@���d����]�i�g�P7l-��@���V����^*-kצ�D3��WP��Q���p�a�ax<#���<n����f���I�q9��DE^���f*a��c���=�P�6lHv�I�(I�r���`O;+�/?q%��ʘ�"��9(�h(��ټ��m�Li �z� ���N���󭷔y3CV����|}�i�O��D����*	����UYe�j4L5�OXy�|vG��@a%s4T��E����7�?�>��� �i2ǯ�y)���v{��/E�u���%���ڣgҶ���Κ���}�8��r� �J��[��;�ɂ��$��2���Rpf4�w�J
 �Ec>TWK	��Q$��xG�.�f���/����E�#���Kt����E�� aFa��fzTMٜ9*{�_����"! LC^�63��b�@���g��B����E%��)��\���/��m)��~yo<^�������d�r��kL�Jd���|�(�����T�o�-L=|K�����M���b��a�`�&z�D
kX�
����I��k�N�۩��`����(� �!0�{e�T:�2O���|+�C3�I��S�w���I�����KR�{,{�f	M��,�e ���8�ɢ$/C�1�	�q��e�;�\�42�������3��8z,1a�Ra��"�b�q�h��4M`��h�f���3�Pg �u�q�>8si�� �G��&CF8z�W�d1̣"�2��V]�e�T�k��`H&�L,H���%ݩ{��8~1f˼�e ��|�&_p�"��o7�P�װ�24Ic�5��d߉=a���d����l<	�g��7��C<ه��Ȑ������l���ű@H�z�:u�'�	FY1����rbX�C���}12�o&C0Q����K���<�,{�n?g����t,�!1�!����2{RS*�w0���A�p���9t;�f�J����=�ٻ���L�a,��Ӏr?0,�D9͐$/�!�,��84W��%�:H@v��wՖ`�7�������Ğ^�[�_�|=��+[⽛����0����#�6��k�.{��^���Q������;�@�]�$��5�MB�ɶ���H�ى�+����9|ˏ����w@iƇ���c��7�����D�(3Bޫ-M׾}�	8]��������񶊊]pޣ�oyp��Q)�Hk(B䞯+�(�yOCC�C7�pr��pOO��{��U������A����dy�>! f;3yZA��P��� �%ؾV=��������x��X����
��S9/�2I�Y�H���9����ɠ�ߠ��2��Iz�����
2��s>A�MhI�6�kn.FV;v$���C뻍�~�L���ǄB���%n�Ս��@�7[9�����\��0�y��k1��A�� 36��F52����]ϟ�^�o���۫ �KBse����:�ys��J⊲�l�T&����{��ap�X���G�#L������'��֤h|7G���;�)�ә�m;��F��--���J���*�� ���m5����<�O2�(n¹�^yE�O���U�&�_��:���������*v<��@�؊'��q�@0�ܳ��$�\��S�p���M�RS���U_t���*@h��?䲪���il܊��4QV�,݈�uw��<K2���e5L�WTH��K�5�찚ܵn���޿ŭW� �a��#A\{�p����M���@�kM�� XRG���3��Vx9:��wC_-/��\�DҙA����I$�d���iRSk�!��g�\��!pi���$�uuɹ�h>���@H�
����I�9;��L5���?tw��XK�6���V��!�} �Yf�BT�K��H9��΃���f
@������Fi}��dd%I ������+�hw�2CwqB-נz��E8Q����/���pX.d��䇚�|�`b38�GO=��LS�2j@aP���Dr�C�ލ~���r�w���ع��'B�⳽0]S�^��f�@�P�GK���������?,� ��zd;��T��ܹ�9P%�����d���g+(�\@�p�pC�4Ñ����9�;P��͜�f����Y��S+�,_.�m��Znn�d;;;���g�?�s�~����1j�Æg�U�!ߡ� (���p�"k�d=e�ib9Q�ĉ��:�<�D?4Mn���]Χ�<Ffᜳ�`0����3EpĨ�@(3�©f��J���'�B�v���!�����}Wz�o��^�'Q���Y�>	M?���9R�['�{ů��:j�>]_~���j 	��+VH�����n�ӟ4r}���PK�xP��7鼃����hܸQ���*0, �d2� ��0�jU�AL��#����V <f
�	��z��g2(�5�f*8n����0r�ַ�R�0;t+z�x��V� 8.��0�5%�v �?`��؍�W��B�~��E��F
�C�!�=Sn�0���S���[6!I�!G��p�� �̈́S����ٶ"S�<jg4�(�3%��`��&���R�v�gfX@PE`���j��Ar�ݎf���$���Œ�f���c�d:@)�K\��b���(�2EM'�����\��P��3����7ˡ;�0q2t��&r���\h����N3(��ovj��/9�v��FC:�R�<ϑ��V�0|�X���ڧ����ʳ%+ �	��\p����O�$��Y�+Is&�L���l-~�W�f&��[t�0A��G;wJ���
 ?G�d� 㿬y��9uw������]���Yf��ld|T�+].DQֻ�a�q8H�(@�TT$5���x��oѳ*��n;�ƽ���������3���zW��NG�Qw���u]d�+@�,ᢈK�.�}����^ՉQV�t�k�����'[�7_`�t�������ߑ={�ѥO/U�39�E��H|���\�rs1I��^P�,z�M��>�[�R|���p���o�c�=&��y��5��g�p>������m� `*ر���Ġq���z�CE H@��2� ��*;���������]+,X�@���/+�se��mhh�z+Y�jƻw�V�F�yb�į��2o�<ٰa��E���_����r�w��s�����ܘI����I�Řf�
������Q����R�qߝ\����@$�l_�m ��׏���\�������ɢE���P/xZ��kԿ����R�����n�-e�[�̙#��:9���),+.tx��~�Eկ⚤+%2�(~_ Pi�F��1��C��NT������]��
T�"!��
��+D������8������5��r�c�^��7s�m2���-�hD��f��^ʀa/��C�-�ܢ.Ƌ�d.X�\�7A1�Gn�Y�a?K�|R:����t�k`��3}vp='��R��W�<@���5� T��Y�S�E�^(���f9c��ń4V�X?����C�m3f(&��Zz�S���`�x�9�0���lٲE�9"���g���^

�S�/�H�ӧ˘u�DP�a��6l��f ��@M-E��݈n��3���0l斀Q�~]s��ث:�Z|�ۼ�j*E���[Lp�k0�rP�.��W\!Q������K Z��7����o�BV�)1<x�Z�J�o����-��jHck�127v1�7o��E��9�ձ���oEt���4Ź�i��ەLh���%���g�®ֿ�ao�%�ii̸'�Ȑ`0ReT�F2r@)�t0m ���Z�:����9���bk��� ��_���V�{�Vp�F�LLH�
.j��	����=X��7�P_��'I
%�A�6I�i���}(E~��ٳ�H����\@�|Զ�m�D����ັ1�'mN��FR���A2 #I?�
B{ߋ��0L��*�	F�yh^"ѵnݺ�ljjj�>�w"�[�l�m�/2B���^q����}� �z��;��&�<�Wj^�g�m}�f�d�l=�C2�����V+u���7��ɓ�&�J�s'/����O��믿�mǎr*%����e˖1���R	�E��4{�4#"+lm�6�׿�,Y0�OS|��Xc^��d�bLL|��-�f�k�:5p`��5��r�FF��d���r!*X�ʕ+�T�)$�s��𹻢"�
����WO��ۣ�i �B 3ʙ	�L�vJ���f�ӓ|�{/ʻ(o��^��կ���9g3�U��՛c�ߩ�O[�Ͽn�]J���Z����
�o(�4ùN+..��	����,�*�Q��:G�R�A��[ �l� rjn�D��D��?_g��sk�e� B�-���/��N�`����x<��Y���?��&aL�&D���+�N��N�S�q2��I�a�-si��DE&/�ss���2|e����B�u:�iș&y@���?�L��aR�    IEND�B`�PK   ��!Y$�8�l  �  /   images/aa130aff-16e6-4627-9689-819d55b5861f.png�YUL
��Xq-EY܊����K���a�RtY�_����;��kq}����M2s�9�L2�3�/Z��X�XHHH��Jr�h��[0��Ÿxl���d������?�m����p���d��e�j�����e������ي���&�D�	�F_YN����3�z����k����Ԏ����(�Gǳ��R��7���c�JMNf������a�\w��{�I���kD�b�K@�)u+h��,?I9=̚;�����[�(6-�r�d��CGG�%��+��1A������G �����B���	�A�eF,M��Lo���k�=�8%_<�3��5���K4�AlaA��~��V����6�~nU���٤�:Ƌ]��d*
����W��CMy(%.KL�)�U~3"`��&���Y�t t�I� �Be���qkP��r�<f|0$L(��-+_�a�� m���$�J&�a���%���}$?�}}����4��ۏ��˜
|<gX��m�/���&�f27��+F�lȏf�{L�4d
�"��)"eN��_���`��N� �W��ܥ��d
ڵ��Ϳ:��-�^���X*�^�☈"G��oւ��^���i2���n	�ii��}I� ��M�L_�n
k|��g�^�D���Fg�Y�U��'�Ԥ��������$k_{���A��G�1�F\���uGLvaf��<V��W��f^���2=Wt���\C<�m&�	@�Z�O���g4��͆R����թ�#�7�Ȇ�A&��f�vf5
�"����0��hż_�z�@o*���I�3Mu�l#�c
���H�Z�I�C3n���6���ﴪ�	�,�@_�7���E_��~��ܫ�[&�N4�X��������'I��^��D��;�d C�uI'��;�����L��ږ��!�@7�<�^�����	�ʉ��!Zv�pt6�L(�QbG���Y��XHZ�e�<Z�L�$��K�V�jN]��{��i[E3<ӿ����R¼�`�ӡs@^��pv�Z�#�A��4d!~�D��޳%�{����i)�*7�CՐ��\,��{�_{A���>�Mu]hm�w�bD!�$_`�12Ő�Y�D	�,��&���W;��uo��oX���N��������c����`j������{���c�sH8�0'ޠ<C�ȲL�Q�ۗy�ߡ`��#��Q� ��y��IX��L�J�{�X3�̓0�1�|'��f�9�CC�U{�'T�K�c0�W�&O�BMJ�7&�꠰l�j��������X.7��k���leY#zu9`�4;��w�}U�@�l�`V�[�Zl|D`�eJm�c嶚��lnQ|l��;�l-��|�8�Z�-b�P˪W3��OIƭq�:��KS��d�iؤ�)��)hDסQ����UU��e�K��iKR��@�^9���� ���7G��*�p6�����Ir����1�q3��	
�Fl�I�=m�h	� }9!��m�W�:�1�jC�����w�(��b�������l7��2�~xJ�֛}���F\��w.5��ߔ�h)UV|il��;��cL�{K��ty��{ �``���C��p�w�kz�����I��g�'y�h=;�@�D�{:j^.�m⅊��|Ǚ9����;R�ȍ�� 3����xw\���CTl�y�,u�v�e����Y�(Tc4@X�l?��%:��v�M�(��� 8�TZ6�[��_��Rz�#�E)��i�{�5��.�X�uj}\m�w��~&�e/���H�8���Q�/���H�R��5���_�5�q��i�V��;���~�++�9Q����9=�CK�;G�T�N��㥲b�=;�p��>�3���W��.1���E�����|��Kv4/�t��XTJ��6�u{��%Ǻҟ.���G@���:� ��y%��
��E�N7(�� 2�-���]�H���Z�  O3�*韭�<m\�����t�pz�#�����Ց��Um���C�nĮ�$�e����uesM�����?����pc"a�4u�hi� L���(|�ϯI�L� f'�E"��*٩��ծ� 9�-]�]�������S�;iSKn`Uȏ�=����R��8�b�96K�A�E8�կD�h�⢛ns�/4��b�#5���6�R^&h`�j�y�9w�T��ێ�Gy�x˞�iz
z箹�c�*�_�9��Rg��U]���,.V�m
g�H ��rK[}����цQ�I��X�H�����rZ�y~ 
�6M��
򗢧���A7��!ܡ1�@��I�ĩ`!�j}���%h�	Hm=M��ğ2�2���I	��F��[�!�Myv�LE)v��� 3���>�xj�+�Ҹ��_��a^�h�$�ՖL����q�Rf�.��� ~D��O(h7G#�<qF�[)�������k�mFG7fL�o��k�1ջK����r�W��o���2Q	-��k�z�Phiѕ��"0����u��{���blRxk\�SK�.wFM=gx�)���;��(DCR���=���}���ST�P؜f���M��9M��X��Jlָ�.�1Bf�b�^�����g���H��(�_��_���	�F�(�P��}�y�&(�$՜D�Կ!u�y����e��a��,2�R;���ٯ��=����"3[	���6�rm�E?\L#vO0Q�3g��ˁ��m93X��GS�=]��F7/�=6��z�|�y��0�7�#�����7�}m���4t��`���H�袟���P�N�ɖ��{[���4xʨaO�K3\�qd`��R��sL$����;QE�I��G)o�LQ�uz+v׺,��L��X����%�\��p34p��Ѩ5 �j��Z��g�<6�^ܘ��岓d$^I�@//�!R}�V2qPN��H��b5~�q�@ ��>Jɒ��3��?9��yb�Yř��s���1]%���Pf���&O��O�X�����S���cܹlb��Ya��@E>��7X>�J,#�В��s�*.i�JeyL�P��N���	�@׾q��/"�M�))��u�:�����T؃ZV&���b��(��h5�]�+��9��0�Y`/��|�~�<�����d+�_?{����@�U��bꎘ�״$�P�`oP��R`]���;1�9<P���Ιd��`��rCF"���\ջ�(d>�M%DiJ+(63�Cb|"&��x�xL2%ѼZ����CV(�(�aW`��m��R�E�o�j�SX�r$�h�cz@�S��.������/���kW��z��[���z�K[�tK�f(��z�ôڛ�I�����r��,�*$��;$�|�q���zw���ǜMh =J�"2�Ƥ7���"Q6�˪]p̻�Aզ�s��:�C����w�5�hxa8B�L��n{�?���(�͸nu�$��Lt�z-=
>�EO��M� =�=�pΆ�0٠��Q��e�Q����_����h9>�Q�?O$W�d��/?-��uh�4���)(v�Uh��CJ���/Y+���<�!�Uw�~]PP�����Qǟ:�Ǟu��o0��|j�sv�%�U�d16͉-���Ze��Z�PR�_Y���7�������}���؆X����Q�������)6�	��N*.)>�.�G{��3�L^�u��p)��ÔA�Q��yM����Vp,}(Ll�xh�����---l�PT�ruru�ޥ2c:��n.1�N�\�4�M��3�ť�N,��f�e�����5i�@�Aɭ�-YQ�S���fƎz�
�*w�ÌO�ƪ�����'�J�/���#�%��.���U/��G�+;�ET|VP8�FBM����k�WY"���>ފ�]Rl2�T'�w���QK~���O���҃��b�15fBv���tA��g�q�<QӳRolև̅����A�D�.`7����B���*��R��$�ka]|o[d��J�=Q7�FbnO��I7#b�F���3�|�T�#1��D:��/MV�u��Be������u8T��'�&*�c��/C��̊�|b���,5|%���l�W�d�_���V�{������)���y��4C�dZ s���NX9�[T�W�⍪��ѵ� �"*SPÅ+W!��q#���[Z?��Vl���{�w���	�h�i6�XJ�/��I�\#�)짎��~��x����@�'^�u�! "F}���P�����@f�kM���������`mO��3���((��MƠ5g������본��N��_�b�mjВ��W�O�٩�7W�}I�.N���وa�lF���ʔG���N�$so��]�S�ee���=~뤶��@��N�z�5��:�s���ĕ����R���5֣o���laӗ0���>��^q�������3��2��R�7�$�;;M,ˈ����B�������`��W�p\4�\�qH��� `����1�T)!ؒ�Ak�J��b]��%{���DW$����~ս��F`(��ÑuCg��F�(�+g}}��'��- A��x���6����n���#<�]��a�������{�c��J�,�5�p��qp#��R�ZX�S�/.t�Zr�]A��a�N�(6���_km�mR�c$�<Qq��)~�+���f�Z*pk��Z�f�͞Ff�/eꝻ!Z�@�`ḋ,����?)�*��(�<E"�3/���"���"��o�{�RX�N��/�a��ZU���xm��iX21�:1}�,aS缈M�rwg�xM�u��k�Ѯ��e�k��V���S�Y2�֯�Tw������o���];��nf�/��ŧ�A��\��W�o�@��sފ�H�#��3��m��{"�E�Ӛ�G_�U�]��K�i�,�E���6��tl��$N�J�%9��{�P#6��䓏�#��.�^YSx��WBI���7m��O99.UϹ~!�t������	�[z~� SX]�"{��#���7��4w�M��z���$�o�,lM��u�D�Q���=429~� �����AŚ��Zo�Fc|��a>Bz��
?�.j}�"�F�4�'OdZ-�QB����j�IF���{$��dֵ~�l�EV&y�˩ XXy��DJ��c��_(}��s�T��Ҕ��[��D����Mfod��%������Y��cZ\���$�1�\�Tgp�ڊ��-��I��*p8�C��k��Sm6\�������<� qN�&,&L��0���=��M*�+Nol�X�V�ډ���b΂��z�o�����ӭ�������YĶ��U$��H��)�5�:eW���Z���<��c&j�0�b�m�վ�s���X�O�0!R+"����U%���a��b)�[����z5g��x�$����Ke�����d�@HN����c�܂ח��):__8�$���8�+�Y����JG�짽�4�E�^y��5p\���h��VU٥���h�븏����|��^����ЉO�I5'�V�t=`�},R*G���8Z�]��Bg�X8�F!�E�����t���2;ę����+ݘ�V��L�Cc}����)[�-�� .KfwG���<8^h@`!;��6ͮΒ��z�Z�%݆W�Z>;�[��#���0�%�o~���<;z5D�)a-��X߼}��U����[��̸��W>[��
���D&yY��~�}���cx�3��Ey�1�VC����wv�Ӝ�)1���Ⱦ��L=���V}8�LRo��N� <���5���w��x�4����O�߆��Hc���]H�Z	Qi�{�������ɳG�լٲJ�����̸�V4�$E�2�z�5�|�R�$5R�a�qL�qe��"V������X��	�y_6�IG�41��n����@l"�oz�i�v�ɤ��KlP�*$La��B��g4��i��/��<�:�\]/����d�!`7��k��J�AVf�����Pmܠm�g\|����"݇�P�B�?� �jdԇ�-�#u=
n��m9/.��\����\�]��g5<�����y4�#F��C!;I�@&0S#��T}���wd�@C��{�K�H1��7��,���M/�K>���-N<�6��"�wqN�5���s)��G�q*%���9L�Q��0�wk��w���x>0.A$���-�?�˙6/�PDH���>��2�P����Eiap�13.�U�Yz�C�)|�s�VkV����#(V�ʹK7�������ߗ3S��n��?�p���gҏ8��Bقo�'j���BbZ�%��M;#w�"�⮣c5~���/��IseIu�/�}�m14ƷS��b�#�<��k"Vj�͇�[���V�o묆I��?DoA	�Sv��&��������d�~����6��v��h��=�X�?mΜ��k{�����6�c���W�L}c�w�.�S�~�Y�s�_ٴF�u��;��8���g�����QT�0�ap2�;Z�1''����>���˵X�D�%!�$�ʽc��V�/&^+lB��IJ�(��y;����+<���V�ܮ����z���Evu:��2����=���!�K�[�xWK
�il�����qn��>I���-��UI�rub�j�=Qut9�{̝�#� Y���r��q}�V����� q�n��6f������O������e�� �b����`���g��8t��A�ש�x)n%�W�7'��C]$�3�������M�s���-|��f��9��A4K�l��@F���D�����,��ߜA��[/"*����%�="5=�He;�^	1#F�,"�e���Zo�^?TV����_��z�^ЦE>@�
>�$�RtF��1~vu>'��s��K��Wk�pϚq���A?\7�~ϟ�_�G!
����&h4�[���

d�.����g+�񿩧z�N �C+�ޛoxt��mS�j�����;�'���kpڜ�L�]��)V3�� ���R"�@(����l��t�O�;���;�
Yͣ>*'�a^9&۫]�g�7p�v��W�&�C����C�ޮ�����lloP�H�l���(�����X����}�`���cZ��S���h݋�e�9Am3�P�<(�L��ho�|�h.Ϲ�о'C���F�"�ʉ苃��7�Jpk�xsJ�3I�U�X��V�D���6 �OfQ)R�R������r�l�i��Q�u�)��-�a�5���D{j�b���5{f����컈@����㠸.;����}l���p~�;(�:�6���,�y��{?%�9민
�8=*��I�)is��c{�{�#diۥ��,��lhq���W�!��a s��[q������%�U�?J(e(�T�sZ�%�����>��RnӺ��j�ܿPs�>��l��n�wEl1�u��O�!D�	B��Z���bC�~�3Px0{�#�PR�_�L^��,����A�ǁG�	�?S�א+}�PK   ��!Y+L$��� �� /   images/aad47697-5cf4-402f-a095-abba84463b41.png�wT�i�6��;�#��*��2c��T	ő�z/�k:"U 0��@�ޤ
��z���K�S���~�)���Y�k\�<�������~��B���_X~��������TTJ��~?wx�����/���T����[����j:QQq|���{�����,�tV�3sF:�R��h�W�VNƆ��|v���dq*�_�����*&a�ۙ3�%>�Or���������~�����~�����~���������~�ȾP��~�����~�����~�����~�����ʾ�?��?|�p~̘�����\���*�Ηsp��"��'�&�m��׳���C�d��;'�G�=�Z�(���/l���d
ʜ������K�Ͻo<�J0����̚��#�s>q@�}�OJY�n������dR5�/�|�(��'�����ȏ�c�X?֏�c�X?��k�'����?����=��$K���8b�+Y���L�ug��J$L�R�(���2R�]�������²��7�btU�謫4�
.=>��~ӹjWS7�����y��|K�]U����Aw<)�~���w���WK����b��yf_1<��i��\b��}`�/.o�U���(��ͬME�������Ͼ ��+8M���R���XP���m��FC�����Ж�D%�w��2K��e��7qoޫǉe�QfH>_'V�%�oכ�)�p{��ڡ`FS��GՕ�ᾰi�)A��+O�`�+�ع����U�&��:��#�S\-9l60�f}u�����P_I�?A��4�O�����#�W;:Hj����Deg٧���S9�C;�IjE"w��)���0	*0�du�K9>�~�\&�A��L�#��|���+�R},����qM���딴��e=W���a���W]zx��K��G���ޑ��:��=,��j*0���{t<H#f"��rT���
t�՚^'��k<�	7��xn��_����8´vsa�r� �߬:ۛd7Wmv��V�#�u/B橉��x�p��&�r��ix���v��Ǹ�#GY\��US����d�8�Gf�`S�����y×3���O
��:
�F��[��{�̱�Q��.Tb.�d��gh���Q��aQ�]��_��|�Ȕ�[�H{�ȱdo�7cγ�5=g:Ԕ�X�e�+�e��ӗ��ĕ������h
y�E�6�G�g���K.s@�'�K��Wk#�\�ʑ�5~�7�/�ݮ���*��Xֶ�1��\����xޤݮ\}3-���\�����x��~޵$��"y���^���=�}M�4�P���=H>�`o��9�/�k��i���#�B#(���z�~⍄��Edt���'as�
A�X�G��ZM;������{�?]�����	��,�N|9жo�ޑӲ�[��n���x.AO�B:�F��C��7�D���;��2+w�}����g��+��fHVotìkP���Â��%��a2�p��M�[��w����#�������!v���,�$�.��� _�����Y��� 0��uW���R�(RN\�M9� �ò�eūع�����7ޫ|w��v"l���ðw����Z���o�yb֏L��ߍ1Tҽ%�O����Z�:�*��\�)2�w����eb�x%��T�O����&γ���hL�l��Ói?�8�S�S�E�C������{p��s���RS������@3��9�j�㉪��5��5�#Q��gGM�\ݘ�v����;��3k�H�>��ZU*z�[�|��>ʾ�Ԏ�N��e{U��`,d�愈���(���P�lA��K�y�
N�#��x6��+��hQ�J���8׆-/���c�=�?4ݯ�2O�1����lP���[^�K��C�h�Wp,�*A��K�d�mx�N��v/�k�cg*��j�_��t�撃�	P��1��Ć��m�d4u��e�1E���?����~%b��m�����P����,�N�N+$�� N0�1�U�8�lX��vq#����`o���nkJ3k���A��T�L�<ذP��#�[��'�g� ��ڢ��$�ԕ�f�iZ�|?L)w�u����2�*�$t]e������"ߑF�!�g!)	l�kʶ)!C�C�jQgm�g�J�'��&�����q(f
v��d�H�^O���f��yL�����HeQ9� fC�Ͽ�]��n�l��̶l�Z�_�Ex�۽���u�)+�
�7��ǵ&jF���"*İ�Q=��"^����°1����g�8M�j��|����g3��>�J(�՜c�T��kt?O�uU�����Z�C��:\v�S=���	."@r���ӂrT�O���3� 2���!��y����3Uحɀ*]Hyd��/�x�����0kBɽ�9�)�\�5�KFM�1).f�V�y�+�[��WnV�9٥_�V��+ڙ�-�o&�gM��{�����!������z��X�Y��ײg2#�T�e&�:;���f�k���uQ�S�
_�j���パ9F�cL�Q��X| a�ev���_T{�+m=>d�_t�?���b�./$݄���S������8���O�F���t#�F������vQb�򕸓���=[�i4��û&���ڽ��,ӽ�!q�}��(F*ka���?dӯTu�5q`vZ���mp#�N��9��-X�*�����0}�������ai��Lr ���mWg���IYm���Z�=mRyϘ�R�4��A�J@ ��^E�Sl���x97��Vƅ��F�������zեh�I	�vt�P�'�%�lk;�~��ɨ���`WԾs����i�^N�ڍq�S^��x�O�)�%���rH��\���l�۾s���^c��OT��z"���}��+*#�K���-�E�p�5�j���5�+�m G�~q�G������k"��s�뙺��&.��-�ʷ���b4�����Gl`9�x,X�#,%������T��Y���<�e�ۓ�WR��Y��V��G]���eȗ��L��̈:��¹�fqoCMa��p�����-l���W� ��	Ѩx}Kn�JL����,����9�k[��z3U	-�w�l,�$	Ի熸 0�Z�	�06�G�i�s��+�S&���6��n��(��@��j�Ż��w��V����6�>q2���O��+��T&�%�n_ߗG���$�$B$%9��H|ЮEP�>�ZF����k��e��}jx`mU~�j�y��/eAf�)T��ؘ��ƻ�,t�������*aBn6��X��n��;�b���ų��u7�K
��Hv��S����T��	�t����⧖��
��,T�܈�ւ_�b�'��k�|���(�i�iO��a�쫊)v�|���ηzV�
�A��h��K�C�wQ�s)���(�+�s�� �2��1��{�f�-�}�I�"��`��]\N�co�W�������`��4A�z�T<�<5�u+�[�m�Wo��.70)Wǐ9w���5wѡ����\�>�6��L?�:'�|�h�PP��d���m٥.�GY�g	K��_��v]	�C�b��`�V����%/��O�灐0��6��O��9��&@��a��� 5��8�+��\�����;u!�p�P����H�i1���x����FZ��ϣr��H�J!:O�����z���`3ğC;<`��ye+�^b�!e�bq��O�t@�*L?�%E�}����|���ia�P��O{>m$�E�D?��ǚK�ӛ����$��Y,D^�K.A���K�[����:b
�B
pAׁR��� ����i�(@��7��z|���:/WG��s����&��CH�~�'M�;Aƍ8�uo���0����"����Y�H��^G�n�fN����#� �ˑf�>���2�c��$�54�����у��b<[$2�{�A�t��:��4a.�k:��p���b�ݖ{[�ࠚ�p�q$AN�fh�j���F.oA�rF�g������ �9�P��>O"��9^�Ɓ��
�%ȩ�#-�M����W'	i�\A�Y��$���΅*�t�"�E�A7�FRC�Lp�Ǚ9�+1�ϧ�����<�o?�Q5�����e/�pm,�oz+�ٳ7܉ÿ9k�E���s���Uɡ�!o�����]w!�(f�cH�����Â��a�x"�i%���PZ�I~��sj�N��7t��Q�X���������'}��ފ=�+@��=k��M1܌��u���Z� �_�=ߍ�*�{vR�v�rMF�)fҿ�,`�m�,�i �(| ����}|q�s���BML�GR7��:/7�^�d��I�:f���g<�,�-���.yC(��qV~�T�&�΢�7A\��Y�
��uQ��t��L/q�|�ZuR��WZ����Q��L�7����#Ō�e뼕�m*����w�2�)
!PU�/W�p�ȸ�B.*��ʆ�6��k������*3�O��B���tx����!�U��z�eє�L�c��)��<���#O|�h(��n���9hâ�ⱒ2s�����O��6]�A|����c-N\/��h��:M&�d�vg��=�f���}5�W��rf�Hg�IW�]�0Iyu�J�[���*����A2�=��,)�v[:{�i*�K���{X'�����n4�n�v����!YS�`�~,��aS���;�"_�M�o�I���8<~n�G��%K�7H_I���KT�v>iwL����r�@����6��J oĥ�|�Jz.14}�1�&�X_������WΘ�|-� `��az�\vޠ�u#MϏ�7?y��h󛼚oREٓ���W���v�>�boxSq�2�?oN앁��o�۰k��Cɬ�I؎�����^ �5WT�M�|��;��G���?�6"�B���J�wt�������#��r����MO;������v�n[�Ȫ�+*�9|�j�e%)mƶ�/|O�q ��>��W��')�z1�_���f����y��B��ч��4ss�\� �30�y�qW7�_��/���{)�.P1��0{����m���M|���y�uMI���zۚ�H�R��$�4Th���O�i�������/{ގ4�] �xw6�ރHʼe�QF�F/Y�ߟ��Hk�ڱ=�|��==���8�S���W����T��p�#ө~���]��aq�|�{|��W��-����!3�Iv���N���o\YlC�Z򹛗��CB�佅�YXގ�X"��ӥ��C~�9
�ט�L6����{g�����JY~*1zԜu�D�t�'Ɛ3ތmF!��$�莶k��N)~�� jM��J�,�l��h>(И7ׁɯ��+!˷̵�%b*ˉ�Y�A-�\z��@OO�F�Nm-�XH��VЈ��3F�O�*����"L��g��c�c^0�5)�u��_�$emo���,G�1�C�q��1�������ݜ�߈�(��M�� x�qlb�_m�&�w�5z�,��C�&�{�6*r�RU�d�ɗ��A�K�C���>"����_���ʯ��C[EY�1�ַ7�vy����(�;e�C;]�Z'
��{�ϛ�W�-6$C2�3�x����93vF�x�OхS��wk�k@8��l(��ǵ"q�c(;��S?L�6m,���0�N]Q���-={ �?l͠�6/gw�4g�+�F�<��μ�K��%%w���TC�n[�|�������ea?��t}=E�-��_z]���kf�\M~h<B0��L�HL*�o�O��0p��.���f��EY�&��������oQJ���,���3d��'7^IA�XoCO�#_Y.�S�q��{tn��2?���p~�0�����w?gػ����Օ]��`��zKd�d��Y��r��#��D�h$��B���=���Kx	kB�)"1�Vy7=g��z
Q��V�=?=�LHh�_r���"����4�B�z��U��"+B�a��o�Y���>��c������ʅ��=��`�P2s0�q��av�z6��m����N	��R��E��a:#n�|9���\����d�'��Y�\u;C-�A��}��4�X�r^3�S�`ʐ���Z�Q<��5>Sb��X�EH�	���~a�DW/�d��-�ŋ�$�ҧ�i9�k)�=Վj;�>麨�1�Д6W �x#r��s5�3u�B��:��w?}���(Kj:�
���U�;~*Q�t����B�����b� �mx�	t���g�m�r��r~8�`��cJJ)7O������V��͇"�3���^f,�>µ��H���O��H�B�Y�1���x�O�0�)�:����(yM�s�.)$�ZC�Ȭ����!��Yܧ�3v���s�7>IA�p+��nJ�`���p��96N*��Q/0�j
�ǐ�fZ1��&��n���W�{�ǲ3���1Z����"�k�!�>C�<�K�Wz�7Nv���«�tbɤ/�")�aw���D�鍊g�,��*�IR��_���Pl����^�w�o*h�x�����A7N|~G/����o�f+݁>�R�d�d�-��d��R�OI�ba"��]&M�o�����OJ�ӡ��[&ꊈ�Sn�ʦ�d�����qrJ�I��K������w�f6�TE�AG��bPH�<<:V.ܺE�hk��cM9���|���~�XS1�C�R�2��^3�}����f�GU��cц|��Y(��+@ 	��4n���r!>���g7��|%8�ش���1����4��TkIg;�c�Xw�3ۄ!k�-��lo���C��0EE���{�!��Q�������cI���񳧗�tVlI�w`?�ƈh/���H�m-qQa�ѵ��wBt��. �v~����������1F��]_��'���E���ψ?�'9���J��,Z[��Y;+N��S�%�����[tE(:8m������g�"�hE%s���z9AO��۵R�֗�/� vW�O�N��P9ϝ���Ϝ�.�Ij��,oT5����bo\v�`�)vk�|�9��-�||_���8������ڊZzyh�G�̀��=�aŨ' CJ����E�N5ȗ�r5��NN��H�.��5rP�r�Bȱ�
�c�R��O��|g9�����BMTH�P>\��p�ˤ�@S���NTO�$�R\ʑ�.��8麆E�e��1�����d�� VyƓz�i2��Iڐ��a�ZJ)��P� �%g�Zݶ��A�gG�w�h.hc��L�~�˒�_������^y�r����)z��U��=~����V#���Az>%���ҷ�(�&��(�������w�Ps�J�c{�G	�5�F�v,���kP�St*�m��rJ'[��Rm��������h��G?�Ÿ��ny��n�H��fr9xG����
���}I��o�*=�F�[ ��L���|z�"��E��d_S��!�|S����'���ә ����k�����A��-�:�Hs5w�IW6sY��H����堯'T�"�"�6�7<��I�zI[Hs�-n5!��+���Ch{{˨��;y��$�.�5w��M�#/��3g�2�[����'�R�y(mSe1���}��x 3^�X'
T��[|�k�Y��IiI��ꊒWO=������6�{c�xE�p(��Y��J-#r[�ɴ�������)�3�.�sװ����؄�ն�N8O����nο��B�� �d@�+at�qeȩm��B�^$�Ԇ�(��Wi;­":ʯ�	��i�(O6l���L���6�w�P��l��V�w���Pf)���D����QΫ*;��#݋~��.-ʹQtvl�,":����{T�� �0��d�k:���o�`L!0��0���D$����ֺ-4�44�jܫ�M0?�{;�yq���}���{,�ջK�c�[��[���]g���OlSG�Dj��Mh����+�����f��
J�?�'d�<o��w���}��3�*�&��j
��g�bsb
봚�q��kO�O|*У&G�J�+����`Gw�j����Ɔ��>�Ҋn�<�����c�ׅ���;-ꗺ�%�!z��`|.9��Վ�bҸ���̟� �3�t�EڕECA柡�1����9!�r�DOM�.���"(�n�JTey8Z
���˩�c6[�ō+e=����FĦ9�����e뱱���ǯ��Y`�Hx��9~��(K҆��`⪥��0�R�N{k�L��wM5���W�Ym������G�Wd�|�o^���M���RXH�%��՝B�����!���w_�mnV'���f�� w��W�ǵ���7���cY��r-�wJf�h�0�c����I*���΅Z*�m�H����'�ls4�Tv��P0,�'ꉢ���`���w�`�0�;i�+_M5��2�2�{�x?���/��|�L�e[n�@8u�.d��'��4���h;����F{��8�%�Ks+1��Q겨�6���O�[��Qo	�l��� �B�+�W�xK�I�u��a�R��7x7�V4ὣ�����/���Sni�cG:|�\K�����W_WK�?R���([�],l�3rMĊ�ڹ�юV�]~�7�@C����?)�`7��}�T���}�,�#$�$Г����N�߳���e��=7��|hx���w����-�"���T���۽�Ǭ�F�a���8�Kz^f���irճ�(��_f���,U[�R�`C�E@C�qY�����ShƸ!�ɸ����_8m�aF�+��a�]�y;�a���?k�H�nh��aޓ:4�	��oIc������� @6�oT�Ӥ
�;��a��p���9F��cu�y1HQ�٧o%C��@q��Zc���3N���,ݥ�Nq�ec� �ym�Lڥ�j	r�A_9Xr���b㸫�0�Y 3I�������rJ�m^J77��m#p�FRB�������3箿�녲���Į���B[x��~ ��P+���-2v�,��@��]�ud;�ٰ���X�i�����k|%_��|�L0�E�jmNv��)x��G-��m_J��t�*�ɻw@~�q7k�4k�iԕ}�l��43#�����aJ�z�צ��~�;RmI.�<9�9 ���pȉ���8���h;K�t�I�z����fRT���U�c/�sM7)�����?���ƹ��N���L�����+��H!�dm�����`��[2 $��U�M�D*2ŝ3)���n�=��xu��pΏo+����2$���eh�z��`�J�ӚL�>#������;�����J����N�S��|��-��'�F��p%�&K���#�3��)ғա]�)�׸�O�z\��F��D�.ϻ.@�QDqe���؇�������؃&��ͣA��k7W����Zqc�����5|��Z�gQ�C�"���������,=Y(���4'��JD2ڹ�{Gpeʕ���.T�x��e��q9���=Ѹ�� ��`It^j�U|����6 ���8����*�`���}���3�R�I�X��/�'�zH�phC[R���0�KPV&Y7�"���ֱˏ�% ���r�'��\��T�^�r�=Ĭ�3�U�P���f�NT�؂����*��6j2L/�P̡!���)��Q4ԒzAT�T�wa������	����MF�k]�D "?��4�E{�a5�e�Ԡ-�ܩ@�R�u���ĄV���A(�^������&}�@���dN��PkY8fVa9������	���'	%��\YUS�Ͼ�eOW.��2��^��B`Dw��t�wA]�{!\�K�}N���J�tN�ƶ9�4�)B8xB�dfo��C��(3�/�}}����'_ٓ&i���|������^&HzL���pB��Cd�D�Y���3����=q�;o�U�������S_ QP�{��:雏YuF�����5u�������NO|Lg?5֪h�V�67�6�p�7vPt\ך��=3�@�. W�%���؂*m�E��Λ�*���P
ʪP���`�
�
�qN�e�פ�<c�#�y4or���Gib�IZ\��[�X�-�Ĳ��,���������o�h8!��l}��)kzZ-��9��khk���O�	PA�\hC��1���3V�>1�����������w�kN��#�Fi��t�S9������/O(�jm��3o�x����=�v��QT|��϶?!m�2��IO~E�	�5ƛ��`�7�w�Y�g��i%2p8�Z��nsp��_<�fhB�VR�=�e�S�[��?�4����5�B�ݎ�'j�{��Z��x� ��'���2ɯ�N�2�g���]Π��`�q>#�Dg�,w�j�r�Hh�o�FG�ǟА�
��s�^��p`�J�:7��,�MT�r�M�e��Mg�~b�Z��}�Ŋ���4�����*e	����ӳ�5%������I�]g~�O���&�nڦ��c$Ռh���/�MX�}���s����U�=K�ܓ׌灋˂Y���c5�m�&RP3�t>�.�6$��Rh�m�c��w��4�d_#��A�	���[c���'z�ճY�f�pׅ��,�GP���Du�DGO�g���:��2�\���0n��_#ra�J-V����.��{��Ql����LAV牓G	I	>|96L�@V	q�;ܪK�m�42���L(xV(��Yr��m��� lQ&"Gʶ;
��?��@)��5�Y��me��lG��~z�{�G�F2U�n��A����Pd�k xkd��(Б��tx���]��~�>�����q���+.<y��fyl`,/��{�a��f~\�]��+j�����KO��͎3{�if�W_��~��/�3X�[{{b;(���<�G�uj��L|&:<Y9$��Iln^a���@,�ns5�����?�'���LG����^��Z-���\ʖ6Gl���N[���sT>���m�C�f��j�3k����x�+!ʷ��Y ���J:��r�0Fذ2�U%���/2i��::�R�=d��C�.s����hX�.����������oΜbH�]�P"�3�OOS�"�8��o#=.;],r��@�!Ƣ�H�UH�����Z��B�4���^��:���3X!�Yx��`��Hi+k=�r��)�dA%�oL,Y���w��@]�zڼ$�2e�1j0�����x�jG"��ڠ�\j�m�av���D�fGG<��_[���Q���Z̐65��¬Hu���2_�[p�T�S�7�3-��I�w�y5�o��y������@�5���y��*ooJ��U�Ie���"A<E�o�F=@]�'��o) �,�㙜p����Q;��t�X!H��ǉ�����\ȫ8��4��=U��<9ꈫ�+a�C��b�Ni�%��#��Ѱ�2�H�k� '~�k-Vu<*��*5`}M	*�8>~/�R�LG�R)�"���u5�͏���F>�����A����!�ȗ��G�0�H�.xH|��Tg�[�6��b�.Z/�uZ:@z~�S�����tE�/����AM"�au<,�wH�~��
#���CǈybQM��!Es�ᶖ0�3����U4��$U�������{��� ��C����M7 ��X,�K�nS�܄+� a��!���ƚ���,60M���w_���_��Y��cz=��~%)nx�Dա�l��n=Dt#o��q#� i�G��-�y	�T���G;����2�U4A��ШW�'�>yr�k��f�NҨ�O���s[M�������m�g��Dq�҄Տ�q��7�_G�ԃD��5d�A5�t���r��`.S�]Ͽ�S>PR�j�u����\���ۦ����5'����d�[KY&m�]GK#hZ!�[�s�g�jX�.�������������b�.{��=�!�> W��1�8�@��R�j�h%YY��2,f�C��C��՝-� D��m8k����t���>�0�;�TL�b���s��Փ-�7�&����r4+�y!3B{��M��%�駠}�ųGw��".��f[6/q�3!v�DW�+�����m�.�UA�?􎅽�dn����V|��)#�J0`&|���A��]ɚ��ظ�廳X��&E�%:�������	��ꏧniIp�D4���}]/�~}�5�3���,�ƾ�د�V���h5�,�Y�۫�f�^�,g���g�	z4'kT&�/]8~���u��O�k_
,���S1+���O�{����yC��8�xt��T��xV�	��5d�f+� �1�F�W���pD��q�N� ����́)��+�i/`�B����E�:����D���[j5����g��3@r�'��o��I�t57�.�ÎDeFY���uG/�zrC@{�da+x��=Լ��E:��/�X��w�Yɑe~x��K�b�ʥ�����*���ɣ~m���88��7�Y#��P�0��BF��^��8�~������M\lP%��W�@-<G|���̾���jw�E�w���+��Y��_�{�{q���ˎ��l{?��=Vj��2������-���z�]���%��n�����z�JJ���ᜎ�����D���gB�Om�f��s-��]=-����K�Y��h���Or��Ǝ�Z,2fJ�O�]�����Xbи�d�׎6���J�,{���}ח�Ŀ<M�8̘,V\��,�݀�ߞMY�\-�ag�'�{%ӳV��5���rbQU��j���i��MX�o��F�M�!��\m4I%����#c��H���z+����k�C�Pvi��~@�N,[	.9�U�1A��Bw��f���|M4*��3nc3��>��3����Ab���Ӡ�[F�t�������E��B�@tq�Sj��8x��DRDBD9����x�\�!��� �W��m�g�¨�~ٙ��:UH�~�n�|���$�>�U]� 8Ưd�l��)�Oו�JE��⪌��������C� ,�hD18ΐ��j�"����c���`v��J����ma˚�]R�������P>~�q{?/�7���r��vi���-�����&;[ړ�L���{��cu���ǌC�`p'a?�����g�������;�Ͽ��Re髷l�4Nو�X��,-����jl��=��0l����D�(7^��w6�I����{�%z��J�*�V��OɈ�/�wrX�^VƮ=��o�^ך/�L�r�S��B)���)*y��W�q$�l/�}&{�[@����z�%V��U#�6�hm�簅W [u�c�G��\N��_r���kz��2<dw�*�e'�q�%k�/9�b���������`���Ÿj�ib����m�����rS���'Pg �˨���xr9�u�v3_W���� ��bA�K��2>v9�H��5c���?�QG�ԫ����v�#�F)�kV󭔸>���M*��*�z��.���>G�t_�*ky�u���H�T��<�1GB^��H�y���}��Q����[v5׉;�`%x�ؙ<m���v3'�7Y�����_�e�m{��6(]�fJP�捊�iR:*�t��g�s�g{N@����5���&)K|a�'�M��HE���d�}�Ez��\��1����c��j�]S��!������>�1f@�%%����z��;��`zz�z�lQcM̛^�w\��D���~�l�8�o%�@0�n�Y_�6n>��mhD�t�z�.l�$ �`(.{%��)U�t)mF2��o���Ãs_���Y�Ð��Yw��3J䪂���ցd���Wm����׏��\�#Ս�h������s9��ݮ����ݴ�,�4�P_�C����m����!{�	��z@��:�+%�K1�RL�3T<�䷞��y'��u�p�8Ǉ&�^��O�O��xiu�1~h8f[�����3H��c �M�W��K?.���Zj��D���L�z��gd��q���y�h�j�qJÀTe!�|�����i�
Rf�N�t
1nPS���nfꀷ�r�8�G����h'���e�)}6�W$j}	��[ �Ç5wP��8���㜕<�w�詠k��,���7�=��y�����*
����l��c�� /�
�M96U�k.b��`�dQ=���)V�5�gUl<��^�F���=Za)�n�+)͔�h?F��<T�2 �!Fo@rw���4
�3��C�`��ƨ�?ap�zΜ�k�jljѳL�yx���v�Pf�����N�H� ��/֥i�������ԏAId5~�$���2j����C,b���;��>�?�����q2�������<�pqo
�X���Ɋ�#��*P��6�S�, W5u�(Ιl3�=��5�wc
w��L��V'���QQ)��hK>��֮ >�w��Mwn�
�3@�����q��q�*]9������4�k�{�O-�y/�G�+:�Y�ZD(=�a��i�'pmk�P���bB�6k�J\Bt��k�oGx�^=6!�G`dEĜ�E���-������\H��������8�N���h%���N��t��"�>�9�Ɖ9Ip��zp#f������3��n��&¯�P�!��$P�����x?�����ޠ�5���Π����������?�u�לc6f e*����儇_v��ٸP�YK˕���GgRW�w5l�>��·�M|��l��(М��e%yO����]\BY.�]�z���7Sc��ٓ'�f�:}�jw׮_�J���-om#5i�*Ė�N�>L��t��>D�9jY�R���bjzM��㷵'���=����L���g��V��H%����O�:Х��>�F/����Pk�f�
�^=!�)�w���Q/7w]_Ջ��}_�tD~o�6��e�bSb�OSNo��O����zj����Ē�e��M|��j'ܓ��5�E="�T5ʞ������=�Jr�Y�;����[���I��9���C �mi�T>�Si�y}�/�R& g�Z-}%[~F����m~�b��|B˷m+��4�*�\�q��+O2DA���ة&h0u6NR�{��+,��s�=�/J�[�t�F����=�ua�9`�l!Ro��y����݈X��f�5x���{p����&��RlA��F�c�#�\��
�|<Zʥ�}��ҹXn����7���_7Ou�a�6#al�d^��(���8/���ҵ	�5�Έ��8���5�L��;̦�Q����o���V����1JzL�zx�&0�ť�6�aa���C�#��<\��jG���^)h��}>*�����
��m���R����'(��g���2R�Zm��t��[��ֿ��Al����o�m��5�Ey���]��MC���� 5��G��u��N�����-Zݭ�v,�sA@ y��	��0I^O��g�vx�O{��p�s�pjM���A�
��1�G���ذ�_ٴl�C]�{qGF�(ag�
����8yt�|�'��[<$h��>����&}�sF�6��]����F9 ���7"�[j�w���U�E�_<�W��
K62�lɣ�@�w,�z[97 �������?i^�hBHKL��BD��N�s]�]�;�wR{��8+F�@h)M�-�\��4�-��v%�Z�Ҩ'zid�o_�83?D5���&����n����N�%Q�e��۔��@H+�C9ȫ
|���͒�U��Z)�3΃1�'>�f9�Wtf�Tz	$m�q��LZ�C<NF	g���h�&�sR�z<�$�s�4-�)���:Z�u����}�`����曒ݯH�k������Djl/���yos`Llw��#��R�Kѵ�Ո>�'�q��s` &�o����r�i�0@��*���s.
2_�%��n��O֭VVR�F�!Iy@�"�m�kjV,6S�G���P��j'R�� ht��U���ΞϏ��sn�H*%����A?zt��l �ރ�kv$%)���@H���LW.~�YV��iп� �5e	���8�>#�G�6sdX/����\[n�O_iS��#B���0��̀F~+��̭�|�u���A��/5ã��w�A%|�*�9���O���?�(f�Y��X��v�:Y��_�E��WO�]�������*2���z�`������ snN�M#;��(J<K��pDS�s5��ZW��<	WtJfW&sL�p,���sOree�D�h�}�:2����FE�W�ֹ2z���n�^B�3Z喖=�je��#�	�nΘڠ���UFS��J��ѻw��<-��͝�J$ �MzK��P�x@q��j��|�1�ܬ�'Vy)(^��=z������10�M#�c�i9m���J��-T�>��/t��t�=]����gD��,�򧙮����|��c]�u���@��S�瞵5�]�����Hv`5��j��h�N�2�P�����)+(�o�}5�|�!fP�N�<�q�RR<�G+�8�n)��O�TYQv�4���A�$z}|��xlmE�[�Gf��/4;�l�ύ���N���ʻ*����Iz��:�7U�PUZ��s�œWfT����'�kO��X�t 6�̫��
=��ڝqx���� �2�Q��Ҹ���5ۙ�B��!�m<Wj*4��K�D@����}y\��
U�g�$i��G^Mva�1��t /�u�M�zM\ q��	�_��8L��ʏ�8�����<�{��7[���"����#˩$ �l�q
�����'ʋ,����LP�ʳ]k/�:E4�k�u�|���U��2�Uݨ�Lo8��˥��x �0&�<�P�Rt���mfU4�׳�g|LM~�I�*9h�� �fA"%@�����>����,>�ZP}�܍ O�톽���
�ɞ��w*�1.���8��W�׊���-� �����t��C}ׇ_Q!�O��+6ˎ���̀78�}�%�:{d�r��jRb�G 2�,�mR*tlxY��2�Dk�+����潂y3o~4����Ti5PLC��X%��x���HpL���K͖ ֊c�u��U8�[t�"p�z�֒��<�
��[��#%7��͎�����P���}=os<c���p;f�f�wN%~���c;���N9�̬I^�(�X�d�[��Zm����$5a=�����G��偁k��h�F��s���j+R���!���1�ׇ���3�T�ż�F�Y�Z��^�+@_S! p���H\u8��bN�Vb:f�T��jc���#��_�(�3� m<K�|?߸�pf�%��G���ʖm_U	�^=b�̭�]2�R�f^�����nD�]g�{ZTBl�ԏ�=���M�d�`o��(/��v��d����!�-�݂،0�����������2]Bu1.&Ք�ǖj+���=�^�OO�6�}�^�{X3��"3��s1\O@9�H����k�� =��L��d�[V��U-4e��.��{"a�U�!�RJ�PS�iT�G�K}L�$�dn�l��YE�/�A�-�Ԡ�ط�L��\����1�e�}$��'SK���'S�yjc������|�zm���S%w�D
��5k�̀#���ɠ�7�n�O��
UǳL=to9�*v�&��g|:�027��[��g;��/�_S/لz��m��b���4���_�)�@�M�V�����RL���I��!�=��	t�x�/�_��P���nM� q��y<�P�wW(60��mKm�k�0�sã�kFT>���.W��cSY���=EQ� x�I�r����e���R���5?��q`l��ȵ�n����q�JuX��T�S�w<"��τ�Z�~ex琊jO/��,"ȒLg`���6��@c�` �/'���t�ݹڶ?բQ�ë��P�ށT������T�]YY�ܥ�$١��E(���:�cӝQY���C�������{�c��^�����~V������z]
�7��K�k���@��.���H��۴�C��":ǎ����Q!�����jҬw�~��s ��ot�.�:�.��[j��7\��܎�p7L�����:�? 'R�x/R����Rݕ���[�>�1����C�
)�;L�R^���+�����=�I��lzw����s���-��2��K9�8Vվs�hT����z�����>�
�2u02�;��w�|�k/�����2o����#�/c�G�L�6�h�:�D���'1 ����%���)/��<_ � ��0�>._�Ɲz�O�F�\�^�1.(�fV�Ր��V�pؼ��lg7�b�O�'vY���ޫ���}H^_�aMу�K;s_{A~=�}������?�3�wK�(�h\R��	&�1&��=��g�]}P���]PVy�f�����E9���4�S�O%����٩e�_�&��̫ϵ(�0���*��?=�u��e���E>�$~+E��oA���yB �u�?

����go7�v�N���	Q��,�r}1 rt�y������ �;
9�%:��8�15�=�>�$��"��~Wp��}�ܝ���W�	g�	@���x�����S�.�w�z?Z���{�E�5��`���u�d��F�r�I��av|�^�y !� L��cL��]y��RV�b��h�o��Y�=&����2����MB+MC6ǟ�z�MxI:̴߿�v��`��{�<ψ���?���0��
��6[���?���)س#���9ɼ\W���pPoղ���o����&>P���qQ�D���n��z�3��-I��c�2/�ʞ���%���?k�ﵫ�[�W��×��nC�wfe�I����N_��,Q��QbY#6�"����s�Y���t`#���*�N�-�����(�`\":� ���-����g��@�I����Xd��mA>ݛ�C�� &`a�N��"�La0�k�JR�"e@3�z���8��������{ۥ����U����Y$���ֿV�e%y����M��`��s��c��M����bΝ�1c�8OӨ!�o��=�t9�+���o{� �rg���Qw�����c�
<��lvǝ�3��ƀ��_<z����F���9]�B�7��_݌7��Y�lɀ��}#F6uB^�p�ޡ��k,��M���c��CW�v��=���Eʖ���u\���з1���Ą�e�pb�Z�	Xjc�;,
n��Pޥ���VǅәvQ�yݢ0<Z�M�U�@/��v,��7B�a�d�F@r��{��Z�2��f���?H���I-����YxW��5�*r�⸉����Z��Ԥ����=@�����>L���i�U�8�s���j�FW�&}�]����� �I?�
&��'#o0���u��!�K&8����)�y
��~a+D1��c�ɕ&L�o�I�4�Y��?�uI2���pպ�������)���gg �����6�8=`A��%���j���8����Q��r��m*X��WS�6ʊ־��2�E�4��!�{���怟�#s�k�K�JRNJ�>��`o��|�w(�&�+�?ʓ�gTN~r�KP[
-W��6�rfT�g��"q�z�*/�k�'BW� �����5bfT������#�ɪ�Bo<�6Ad��%�fv��vl׮��P�$t�����냤���Ñ�N xs��D��^ό4�=܍$��m���m���mN7"\}9B������6�F���^�2Ň)��=�3�J�qs��L�ՈW�,�I	��rK����k�����Sr�6~��ki�K�aj�)� )�O���\�L��|�ps"�����n�����ZX���f
;��7HW^sx�;zb�i�+&=��3�=4%�����e3ҦO�۷�<w>2a�"z\��{P(��f�S�H��YԄ@�d��Oxt�C��%�I�f�~�JP��VLM���#<���4"/�R�z!}�!'A��)6Q'���s����YJ� ���:�ݫ�A�s��`�-l�#,jc��%��b�G���L�� z|���f-Wb��8�iO0�
S���4�?�R"���/��ʮـi��^-��>��MB�j���gApL$^{��?��ln�;�}���X���4����^��p�h�4f\�L���$Hp�~����騛��(�q�Bmǭ�z��Z���C���P�B�.��{���B����R��%���fO���']n��g�U��4�Z�p�5��N��/w��Up ��z&�U����nCyc(�$��g9W����G�{�������;࢝q6�'�3�n�ìAd�>=H)�:.ۏ}Ks
�N���qK�u�+�-�"��۩�_��'���6���6��Ƶ7��4X I�/_9���+��0+���ejql�hsd����l��ݍUwS*�ސOc�i�_��hg��1�~|�E���H�|,k��Ĺ��VBwK����FB<�f���jd���|!�a��-PZA���sa�D��"�SBHN�ﻙǍ��~��8��OcNri�J�A��)��*T �$46�j��U>cu�P_�l7��YQ#���BN@��en���+.�uE�BS�E�E��D��M��k�����ӯ�U\a u�+n��/,d
+8�i|3����\l�w;�{��*��GV%���+�.g�B���b�I�olnpE{�� eʝ�]���W�w����[����!����!�Ғ�'Ѷa�	�4��<+2di�&�7�X��+��{�տw�J����֭!{���E�R�L�����9������z�о��>D�[Z|�X-K�;r�Rϴ����0g�g����6���i`1h['��,�G-�2�e#^�ְ����[���aL^��[h��Z�?i
}�a��Xv��kz��
ĀV�%��#��G���%����.�g�Ɇ|����P���g���}��݀iL}u��m[�`��H�B�z���n��v���� ;S:���C/D�/JX,���2f��)��9~�k�:���.��0^��~�2⡤�T	yI����?�FE��M�r��D����uc���r1#rN5q�B|�C;���|��C��i7Z����c*6v�T��w��wyG�Z6SY��}�#p��s3��`�5i)���Tx�������%_�e������3���r��������c=��!���x��_��2��m���P6����U�K�H���^�r�hk-�d�}D�����bq��þ$F��Jk��75"<����n�)!2����o_���6W.�z�vyV���%(҅��[����-���:��L�V�b()a�$-���up��oE�F[�n�k\\|�{Z����,hi�vd�d 4�N�tݮ�����u�v�x~� �hI;�~�ԣ/=�m^��1V�&qPc[Ϋp�-{zSj5���K��{�}�)��f��Du�L�,��]���n�,���`��;3�GO����`��;5V�����ln'%V��h�_?��&rh�R��:�]�����'Y��v4oR!�vǨA��sBh*�ƞC���\�ʿL���hp�^����)H����U�� ��=�<&M�v�_����8|o�pX,+���҄����,�r�WP��Ev��R���-��0�5|*�{��:�=���`Ux -s�����P�a4�fxز�G�G��4�Qa����9��'���HP��{G4���}�H���^;4��������h�2�i �|�H^�Y��r'{RZ����ɜ���yx>u�VD�
 *YǳomA>A�	R��g����P��x��W-v�[l͋�͕�q|�:�9�?��?�-X�?U��C*�a��T��N�:9��M��f-�q�@��韈�81�m%��
�K�1�7��z�+w�G<�3"J8C3Y��@�U�؇?��Ѓ۔�P��Y�[�&7���Go�yZT��]%�g�?Xw�w�2234)'�ΝU� ��b����gC��o�ϼ��z�k4j�G���ĥ�:�����i�z~ކǺ=8$�,�@�N�����Fj�w��$~l�VG�Vp���*����ej,��^�e5�k����g��8ۯ�."í�	�k"���_`��W�a�l4����d���~�8��ʣ�&f.��>�����
�ވU'�Ӻ�R�r5n4-vhf��G�,�������ЄC��h/r����ݲx)V�X+ɭO��®�T��x�p�@l�����=F*E_w7CEK$�H;`�5���!)�K�U�}j�Ǻ9[���*[��6#��a۫�AJ��h um
��e���]�'I$��O�P���o��3��q���e �
+Wǘs�Q��߼1�L]ݑ9Ԙ�$���+���WC��2c���ͥ�]�.Jk�{���EBR��Q1vL���T5�ӆ�8����g��?�X�����������X���8�6D$��ɒjQi:+
���Y�KO�];��F�����}N�Զ�p�s��x�9Ah�w���w]NU�l\���)�*��?����Z�=������Ig�﫟	[���@su�CF�. 2�2�c�C�&���@���ծ�Tp]t��al�<�?mҘ0���A��]��<@Õ@�,�M�T�:wh���P���
(37{!��M����l�1����u*���T�o�xF�\��\��b�b78���R�Q���c����;K��Z=ɖ��$��e�Ԫ� 姺쭝y������g������!�jO�Zmb���sd�o��-c�q����K����'^��0�sI���G0xÏ?�2.w^��+���:�\�v�g�W-@�<X���,ÃÈ/ˈ;�Fai8��s��1�m�0�E%D_�b��C(@� 4�HK�+�3&4������B�* %٬�:�lJ�?��Q�����p���Ѫs8�ׯ��{����S)�=�]�̮�'�B�+-��?'-@���s����v]�Y��3B<�_�j6�g6�L=8�
d�t
B�Gޔ�S�-a�J�� ͒&vv����I��0.��Vo��]�D�82������!mg�����+�=��ly��T����B:��eKl�,�-+�K�Gc�^}�t(̈́k���M�q[gש�u([�Kv{����8&���s�y��< �(�1� V
���W�N�����g����H�%3� U�"`�g7,5Z�xlV��Ց��ͪB�
ڢ~ێ.{��50�Z�l�ŕ$>��Z8@5�,���&ٓ���sX���$�D��ō�H�C�nva1q�/z��O��y
�[Nu?�W�Es�ΰT�]V��o�_B?�6_�A�1v���J�h���ƿ��Q9R��:8ד�э�h t;��8�l��\����3��vl�Ƿ�	]����;A��D���q��s����dcݽm%ԐZ�gYN��k����#�=����|�ŵ�
���O_����ڟ�\���JI�����Θo�c��w�˕�*�#�}�����Th���r�O��-�@'%6�
&�K��o�pn_�f��:��?9�oc�����<v+8�E` ��^Zz�ȸRh�~�� Ԉ�������v�<� ,�GyG?K7	)�ѻ�O���uȶ��Ӕ�����U�0b���M��L�+�ƁA���kV;�J�g���ߧv�����E���~�&�	�PT��y�����h�з�fhg�C
	�[嵢�B&�g".j�QHo���A�{�ʹH�����
��ۥ� ��������+�UZ������0��,�&�ρ�aL��<�N��f�~�*����Y�M��W�b݅FE@zN��ތC7iNsK$�-֙�0�����jo'Pm��NBj.>������_SC�vP>��R���ǆN���Vj���7%��H�O:yW?��`�|�.����T{V�1�~�b~
��wa�0����9r���g���D��=�"�l�����\�����o��al��_q��fȯ9�F����I����o�PZ9���?wl�e��e(kw��v}��ؼ:gn%��iɨ���a����il��̧�o}�<�<�t_�(��A@������9�K����*/�����b9�<i;��;��'����i}�(l���̩v�և�J8`�Dfc�h�����ꏓn�UlJ��/'?��	�Q9�QU����~��S랠��z�|�-�p_n3�6&��a9S7���l���~����?�`cZ�`��o����>o����\���ѽ�����yCl�
(��ˢrq��}�������;���Zfɼ�]�:�`����²ژ�_��,�@�4�e�����a�uVH"&âfl���RN�{}��q��6���H��E���3>��C�'ݼ�6��cs�W�i��lZ����t�F����0��:8���;i[�;:�oµ�wٮ��3~|���]�ZW�K���!�r�,�	�Bګ�Ġ�^���Gu���V�E,��s����`c�����"���ؾR����r�r���`{H,{�z�����a��q��AۀN���Y��:��$8�&|�~����Nw�͓�gX�g�׮~ϴ_����|�g��R1�Q�	{���w�����e�@T���<���t�]t�����hu�d�8�A�I>'\ @�4s��W4�>��{�iK�ci�G��\���T�W�U9Fߥv��3_6@��~=h`���h��PuX+�����"�4^O�ߕFK�w�"�*)����Ӹ8�����\v��l��k�&�[B�����۹8:L��o@J0R���aƩ�l����83'��6 � ����	��,{&�Z�W��TY3j�.,<p'e�'� k���|���r��'��/M9��pɛ���,���A�&Q.�2����3�hg��j�m�I�V=���t�\��E:�M�%�n]�S�е�.=h�l�<&����\2���j}�p��?4��>���$��>�DVIs��o;{&��]�,kbZ�Ǹ�V�b�{���i�N�]�=�a?Cc�J�k{������֘̐Wj2]?�m��][��t(ЪĻ��E	�uNq�p���D�CY/@H��c����v`L��z���>��y,���+�^�dP�h����	ԓ׭@`�Rd���$��؈K���`�v1?�*�c�����[�{��� ��P)�zx�=]&�*�Ze�	��v8kJ�H��V���Y!��Clܛ���.g�;¨�eTo����,�=G:���XK�!®����s�U2�r�d�-�
f�a����<�3L�C� �Cc��>�бس,-���V�Z�������3	����{�jl:�D���VΫ�(�_
�85őc��r! :��k�I�5h��+;�H J}c���<�������8UhS�
Ģ*�U@D��y'�8s�c_�}�L~էn����Q���ߨ���z���^",�n>�To�B��ͲvJD��ݫ�% �o/�=T?�Ϡy�*:w'��l|3�_�[�g�:rX���`V"��l*���3�X���ۯ@Vk^ĳ��~b��4ھ@Gn��8�]/�6w}"��ԟ�ʩ���'<]Ӎ�l�8l9=��;Fc=�2w j�~u
��,H�B6�����K_ʩ���Xc'=_�@Dxp"Pi���܉��ˎ{��K��b�.�"���������n,�h��o�Eъ�� ��vMi+�1ʟ	���9��~��ȉ�5�I=;�;L���L&�~'���UcMѓ�H͜{w+��E�$���G�t��l����06�a��:�3`�����Ʈ�40������a4_���Z I�(�A6ZƑ��1�/��0�ИƔ��|��_w�n�d1�0I�E��hcS��ׅ|-�ʟYeE/�P�Y�M9��C��3�=���>������e�����x��-�dc��'T��Z��Րx\=��d9"���z�Y�;�R��Q�,GD��^Q9׀i;D�Qt�0�5�F�#����W��Y���W��R8���){\����S�z��K�z�
i�.F0���V�����n��x�I��As)��߫��7[26�?%�6g!���Y�A�D�OL�Fb�Yuy�2 F�
m-s1�����/�;�w��$sX�VOU�q�8�g���>L����ż4�II:L��c}kܻ��I��+S��藿��S�.D����md�lGf��>]0?�Rsl����L�T`a9!?���AװY��x�%j�A
s��:��g'&�'��2�s<�������讎��<@Xeھj��\:A�P^n\ނ�ݘ����D,Ml���{�������z���n�����B���ZB���9"lsh;#]�~��������^Ċ"/R^m_pQ<�C�wȏ�[c��5�[����������DDJ՟�3y���=r�h'PG^nx_��������/BǥA��M��b�t#�� �%}���6�E�����V��n`�'���:��K<����;�E���d�h��<��eX�*Y3��G/���mB��h��`5�U�h�D(p邕(���O}�C��T�jfɊ��ү+�I}���D�C�ޣ�`�j1l��U�	"�� 
�=O�QH��eѫ�`֥$9s�z5��VuE~��%�-n�խ������wȁ%����c�+_qAt��o� �m����"9�v`�<@
����!�hR4��H��qIz����0�g���6��%��?�wf�߄��Ӻ�=� ��� A��ů�I佚�&���˂,��.n�V��`�j,��h��m�����k+΋��%�.�ZJ�
v�x��q]�E&KBB��]S��4���
7�:n��ߣ����;��VSAY!�B/wTx���$[��:1k��Ł�DU���SX,��o�_|�j�/�T�6վ�p<���B��y��c�Y��~����uL|��;YХYy�Xn�T!2Lf����.���K����f�V|�s�A�[�B��L�x�4��t�dX������Z���4�%W����w� �f���<�O�o9Ԏ̟�5e�x@붼�>���=A�e\�h�pV��)`*�0�o�F��b�B���t��8C}v6n����=�?�{6���^��I`��ͪ��tM���",V��c����wY 0u��|+|��ց,�A�y�u����zkͫ=oU��5]//VWQ8�`)V��a[?���8�k&%F}�����!�l���㥎ڽ��7����I����P���Й�Θ�2=��"'g��Jkw,۫]��&CH)Q[�A���m���{��^�����C^���}ݵ��P`Vl��Wn�y�d,��L����������T�0�����_#��Ǟ�,�%`1�pU�T�YRآjO���� h���?(Y�������yc�\��YX4}����/>�^p��j��r����7^~nw���:��; ���V�,�0�@.#��|�ݐ�013X)]PY-ړ��xs�<���ݸ3z>^,hdz\-�o32��Ǖl�*���!<2�������F7�1m�F���]st���F�^�%-)��$�Lԥ��jQ9�I�ݙ{b���6gD�R��设$wӠ�b��X"��}5�g�W�fk-�V�#3�O1����L�ح�xz$Č\�]��b��BK �K��m�0�w�q� � ��O��*&�4\?Z7���y�����<�\8�g�n�w
U��V����r)�r��P[�=�14����
=�h9����G9�4Ϻ�`���r�Q�BQj�_��L�eٔhV9?��{ �0YU�n*��t:Q=�o��g���lDu��L���k�����<�ߒ�7�/���6p?�U��f4���`Ajʼ�X�]����?`d5��g9<�����7���y5�UI�{-��|R,Ψ�8����GJ]6����9�2�I���``�v�ی^ο�6a1{/���&��oB����LG�\͜�k��m'+Jp���v������Y/��c�k�k�'
[�F$��+:��p:4�@l�ޖ	�Լ�tt1`�ް�p?�q�/����f������,�t����Hv�-y��yJ��e7��թ�� �ɓ^�)����E$���]�����Q.�p�Rڷ�y��r�j����� Q8*'⻲s��7T���ZMM�dms��ԥ���$ș���q7(l��w�.�@���׻�`����D�[4xL�h��]L�У��{�F���u�w���H���u�����u��S�붿r
c"��o���$���a��鬱�u���`�˃1��M��f ���G�ۋ��B�"�C�|�+�qs��+k��ͼ܌x߂�w��
�ˤ�N:�(�zx�������iwW?.Z���]T�r�dx4\�����u���mz�]���ٙ����Q�BC�����?K��~��y^;��Z~:b��s��O.��d�ܾ�x��߯��{N�<m�6@2�AH� �=�y=���Oo���Dk,
N̐�:��}d�y�t�`�v�8��M�<�$�,[>����Ҥͭ�FV���$}�'~\�����ӊ�i������X�F����m�tؼ��IÇ����0�҇s_��9�4���q��]U�}J6qte�;�E�`sa��i7�mYp}S ޠH挺R�����I$��G�?>���1��D&��Ct����{W�^��ZF�Xۏ�hh:I�2��T.���tp �;ʸ$;n7��C�.��fֳJ)lBy�P8�\5s�"*'�Z.��_��A$��]��bm[L"Wv�t;�vu���L�������Qb�Ʌ�{�:���^��21��0� ��y#MD�}�e��ٚ� N����l�к?�����T�E���P�]L/8�:4z����l�l�Ʉ����((���͉��I���:5�>%�X�`3�>�.�%i����_O�K-�11���������{�3��Y#*�Ի��\j9�z�fWg�Q�7���U&�[�Y
*Hy-~��so�s��χ!]�2�z�>����I�s2�,��g�qÂl�o��F�>����8�=�aa���q5!��Q�����8���f�?�VA)X�闓}/{V���&�j��{mj��'a�U.N�����2���i�h��WSm؛A��i���J����7FN�@���
&}��w��w䊔#��:W1���=rNc�5�}`�G�f͞eR3�0_��ED�3_���������@D�T��퇫e�Tq���`�{�����A>�v=��k��ށ��Zf�VH8��B>6���ں���/���Q���ݡVy���=�[yS<�D�ZP� <{�-Y�/����d?j1�X��j�k���TL�s@|�m}qq�� ���j�Xg/��PHr�WƷַ�2;�鹖�=`���%r+�-ez�m"P54x*P� �QÏ������U�g�� ��+H�w�]u�B�:4�ٯ�ǟ6n<���5rRR��R7��J�c�XS�%%�'ٸ9�7���,/�)c�f���$$( �l��n]"�=o:úH��`L[>TY���C|���&���OԘ��RZu����"J�n�F�ÿ7�`��CA�<���]a�]\�9tԄ+>�|�`�pfc��	]��A:zǉ$2v8v/��k/l�p�'�D�?�lR|_8�_������P7�o��| ���	�����z���zdaK�DS ��W�u0�H�=wr28g̡�8Xj��+	�nT-4D���8v���E�,"8*X�	�9��}��t~\4d����2��Phrw�V�}#�g��ſ�.�us��f��o>򀿡���\\�&�R��b�����8��%n��kA�F�ZO_���7�FJ�v�h��[O]X��\��3(��O�o���eP��8J�����'�~�*.�{����� �$Q$��[�\?�e�zS�VK�w
��YV��؎��rYc8����Ԃ���?gʢg�|e��4���ER�m1�Ѭ���W{����8 a�.d1L�1�
��I ��3�MF�I8a��6%!<~ӄ*�&��l���ģ�n��U��M��j>��q��d�!��~���O�6�����1f"�oɁ=��ɴ�`Nda{���V��8ũUE~���s�X6ݹ=�4�m�����I�c��&:�
KwuՒKj�=`����j]��n�N�' 3YubyǼߘUm��$��`
Z��ɏ���K�G��,��U�`$�C�6Rk�eH��Q��<7��E�oz�qN���5l���3�6�����ډ�,-)��A��������'e�D���|M � ��a����VSs�A����>�N֖�/���'R6�FO�~��Ǽgy`��U���>��@�g�oz1� �q��a<9�a�v'|����GOXPܝ�Q����@��1�IΜ��c����
���cNڟ��;+	褄�MJn�3Y�2����r~�������+�R��>��`��{�	!��˸~�Z;ڭ]�	����<RZJ~�� .Y�!�=B-+h��x��֎W�J�b�168������n@�4ܨ�����N�3��7g��Dө���O�&��/X������.�
�E���ї�o���?�ү�0| ��l��ݜg@�{� �4/_���Z�0�J*ϳ�/���>�1��r:��[Pk~E���Nɸ��Ԑ�G4J6MU5��WC�\�ω���U~	��2�֟��J^%����ШT�?ljaѠ�w ��N\�E���6۴��OJvl�Cm���iҢ��W��
ɛZ��IRh۶��֟nTn��5�� �1�	b�|�kq����{��w����L�������|�.���_��4������Q�;�
�k>�[n��k�� d�-��>~�^�z�2��gƇ���UH�RR+_�b�ڇ0j�6@Qv�q�-�c�����#���8��[UĆ�
`귂!s�#S`#���[�Rn��_S��+�H��v�#b!w����o׾#�gt�������]����-7s������@��T}�,��bzI�G����ו[z�� s�U�ˇ��P2�5�Vs�hW����e�>8��c*�bci7�sgG�]m2C.��bi�U����ԔP��ɺ��Ŝ�]��+���K��5����9�����I���.�r�/f�1iǣ�i0O�i�+�ce���.z~�c��U��>��wZ!�ܑL�|�w����x8yb`u�r��a��}`D��p�%L�2Њ�ˋ�sj�����(��iñy�б�9��~�u�/� #��%WE2i��j�w�/}��"�*_�p��J�n��
�1�>k!@�v�(���>�a��&�;�wQa;����O�'u��
D��M�i|L�ꤗk��CL���t�& �;�$��� ㈖6W�i/�i��({G�]Z0�����_��v5v7Se{��bu#���r�[�%o��t�~��M�<��9���w�cb��g�W}�ϤYw\��i3�&���=0:����6���}'���bC���l�g��V�\�?�qC�r����S������ݘ=L�]�y�-y}n���_Y:���RQ���
F2����8�8~:g�i��r��A����ǧ,-'�f�Bh��I��=���k��[`�~�|H6��G7cFj� ����c�%dq��#Xc��.�=������_ ���� �zm<�9�n����,�N6����S�Nu���KKzv�J2���Ĝ�{��Ts4:3�),L������O���/�����aj�o2�9"���^������>����H��#�R+��]�i5a�k�b�����Q�Q�݆@mw-h���w��r��ӟ~���U3�0�e��<~_tO�{ C�~�_)�� 3o �R�G5�јN$�?/p /E�Y3-kC~��8���1d�l�xܠ:��_�}̧s ��c5�hIH���;�P8�j���y��Q������9��J3�����P��b����pS��%��Bv�'yo����  u�G��=uP%X�����#��Ƽ<N3JZ]��V#�@Ka7�����'��z\C���0��� M�޷�m��)$��DaϺ# V�';	  |������DJ�JI@��/&��o�j��j�T,��K���xƄ��?���|h���s��ˮ��K����7�T�Q1��P�VqP��+A	���n������V�@�U������If>��J���a���a��x�u~�w}�@�u���ԣ{xg�����t�_\�U�������%r���sTGc]M�7A6�u���c��.ԞcQ$uu���:Cmc�ʼxh���vM�su���p��`E*}3�Ak[hV�_�d�����&u�V����]�ov�?@�3d��W�n� �
(�5�̖�u�F�L�>�u�)�}���@۾�v?(P{?@Lv�)�i���Nw�0�;���$Z��U�ǜG��cO�`�����YK˨�{`�J��������:d���?���xG;�dP�����]�\�������oz-�h�#�{�)�B:ߥ�V�KO^�@g,�t���?�����/A�A�Vjb�'3�����t	��R�1�����c(�9?�.?���Zކ�'�{U�S������^�
�5��l4��U� T�ĺ5l��Q���[�]���2D�nyW<A3��J^��_17rf�O_���@����,�Ժ���D���XۖŦ8v*�hA��(���S��ʾrrէ���j�Ő�=�wqi��G�5����f(n}��ܕ
�t�[�P<xk�e����TY�b��eT��'�X
?_#�}ua�vWG���;0InYhǡ���Q�O#��{%���� �K-�@3���x%�m+�����Ղ�YbY6c�h���Rlً�JΥ�Q#a-W�1Xb����6�@�S:/7@�z��d��Q.;��I/�<������iW�W���e�! 1�j�H ���ᗡ{�'�nU >�ҐHLf-F��2��C
����]��3�Qs�C�c�n ���s�h�nw��*� i��IIYa9Ǜ�����8�}����Qwմ�Y[����N�T�ǔl��^4�os*8j{I�i6y�f�J�2�>c����%�Y!��������~z� ���5W�Z��{�jg�B�M�c\�N��!��qd�@��*�ul�����% �\��9�d�u;LS���4�J�o��L�6X��I��֒�t	K�ޚ����v��pnlO�:���$�}<��X��ٳ����^��#�Vb��W[�v���`fά��ث�8��4�B	��e-�u_�&�a��Nc�V�"��8��w��0�&�����I�;}I��a�J��1}=����]*��p�n����o��i���7)CŠ�U�bM`�� ����#���������q5ѡ:_F��,��z��O� 8{v�WO�qs���W�̆�����k3�>�GG��_��i���j !X<���9��A������d�δHY:J%,nU��cYk#(8殳kI�v. Ps�G,�N40�� �$���|�,B��������P�<-��lC����������?�J��;����}��u�l��%-������w%3�Y~cӆVXMA��e�Nw�zL�n]���{��O�6[�M:�Id*�v����)��Hvq���cz��e�֏�� D�ų�ߡ�+fS��(�
��%]&@]�����,�m�0�;r����+Y��{��ƃ��ONȿn�jo,�d���?��󂩕Udz�"�"r��9LW�$U�A�+�����ٌ�:���ߡ�8q1��:���%�R���=qӐ�0e�k�a4�l���[��솮�Fk(oU(���~�w��;���x��?�Au�Y����%�ٴ��Xzz���#�a:��û|h�"=���e���d���W�°�Լx�0�}LG�$��P.(Z����D�'T{�o�ܣ���܀g*��RP�5�2֗L���;��)�Y���ӊ�8b�RF�}���J0��	��h��[啨�Ͻ�{��Eq��3����h`wd��_���@꬟a�����d_]�$����n�n��ƙ�?M���=�L��|�H�٠WZ����Le��B\�*�m9>�*]q�J:�nl�D1�%C.ۘO���D@�k��\����jA^(U��� z���h����W�eY͜���/�f&߽��޼.^U&Ņ� OQ���T]���Q��2-Yj�Ļ�RW�WVe�&��������V�)t"�U�V��W�|-�FzZ���lV����}�3P��]���<����ס
���ր���&^/�R؋;J4�q��>���1�-tU9��y-͟f��B�
�Tv��V�z�/�K 0b'�������F�ҟl��6f�SA�F�� ����(7���s9��̀'Y坯BY�;^f�'#j����	۩�������*_cƋ��5�[�9jM����6t���-���F��1��`ʞ]I��/@�ٚ*��xKdSu�2=}��s,���_j��2,�:���Z����L�N�Џ�P�^m�mڍ�x�1�/]�4l��̍�zh�=�,�Ad���&�w�ܒu�������Eh��t]���Ը�__��3)g툷�1bU܋��G���0��<$i�ao�� ;��$�ۧeX�~Śf_����?(n/�(t�1BȲ�fu�6}��Tc�=��- N��?վ簯koi��y��HQ�4��a�j�y�c�t�X~�ϕ3��B��Fc�%��%�R�y`(��s6��g�"�Ƣ��VN�%��!D�GMpgک��uv�UQ���߄4JYՉ�'���Q 1�����F�ۀID��??��y�ެ|'��� 7F���V0�Sl,}G�mrb��$�u��>i˂�^Y��6�{����0�8��O(��Yd(9�����N>S��m��!,)��Y���k]�E!������{iC�l��l�2U��+�,L���vv�����S��%�*}ߍ6�s��PL�w�x��IC@��8�tx����sڹ��<��ޖ�����,Z���Le��ܲ�V��S7
�<./9�_K@MSb;Y3�F�F�[d�@��9�Y�ᗁL��&ƨ��͗7C����S�����7<ng�\p͉����ۢ͒��s�`�\^��%&�=ޗT��&�ip(�ߜ��a��%�kw��cҎ�e\�8��l���s��e�Ia7��tJ^������wIEъ��I��Z��~���6neH�B0��嫹6�tޏrrf�[�A�-_M>�M� $b��O��Mr\{8)��3�@��{��ʐA���Ŋ�?t���xz}��6� �|-����m"��NqT�:w})����\��-�c�7���=^�ZS5K9�]�X{����e����$��g�i�u]�Q󳞁�I�>zҧ��vh������qQ$��𸸀Jr Q�]�$Q�� �"� 9���s�AQPI*9�䌒3��"Ir�4�0�a~U=��|�������Uu�9�[��7� ׼���嘪�Pg%�����\��m����n�-�{���/�������"N����S�����,�ŉ��J�D��Q��`�E��@9�Ԑi��A-�$r�O���te��j��dEհ;�&Eu�5ܕ�ӏ4=�G(��(�+�cx���b
��y޿/�5Y������-�ݻ{Ms͑,X���O�p��?Ű���&����T+����s'	��wq�t�Ě�6C��0��N�2i����)�O��p��1��$��JE7g�mѲ����GqVI���Be=(��������-�k3`ť��Ӌ�7'�����*��J��\�K�9*������W:�R��O#]TvJ9��n�+ˀ�D�B���g��K'�nE�<2&U���h�J����DM}jsŃ��m�R(� R���Toh�����^F�s�;A�b3�n_Z@��
�&R��NͩX�tpM%��S��DP�V�zp�k��B����C@�M]~�X\������p����ƙU��ߚ��\T�g+W�x�����#��Ovg?��_�r���?bǕhjy��SE�?�#Ҿ��ʞ����q�������fU<���y?ٹ��#����YO�럊ˬ��!�wh:cgy�V�;�c��:?�R��n�!�e��l�Ad<�0ǃ�<��Q��*�7�jno��
�T�Avd��������>���X��rr�ZN�0��xF��u2���L��{�3�U�5��kBEsobBf�3gC6�s$@�8��&�Y!/���'G���O��WGG `���[x$^����*�����E���E����)�M��Ծ�ۼ3��@g��l����Q��!�:zb�B! ��%��!���tw'Qe�!]j�Z�"��*|��'��:U91mC�zu�e=h���1�<Ms����˟QF��]oDX�R�Cޥ�e�����$2V~���x5j���<#7s�UÚMT��T+���)6���5X�:(H�ฎ��*7���!ۏTn�*�{��p���������D
!oр^�:s�/��a�P.L�j�uX����ޗ��w���_��C�w_�n^��Y��	����%�r��х��@�6l���(�T�,�R�h�y@�}���g�.B���'�ծF���%k������xo<��O-�ziP��:������z��ӝOa�"�^To�*RNqd}烮��nX<`}�O��3k���QJyp���ȇ�S�&z�X���d(����wǚ^�@CD���6t���$nӛ{89�w��acz�:zN�X��s�|� �v�1�,$9�dY��k���0�O���Q-<9��qw�X�R<E�$�h�W6ܮ��|e��ˑ��ٔ�瀼t��J�2GL�-��T�	���ʭ�$�+e�*u5;��R�7��vܕOfwd�������:$l���Kc%h�+�@G��]���1�����cp� K�	��K>>'3?U��YleS���Q7��a��ٵPk�Y��^4�/�B�{Ng����;�����q�MSٱ6b��1u��f��m��Dt���f��;!�x-i���ܽx�}���g�'�6'z�)�_/�4z�	~��2�i���`wP�r��BY;G�v=���3FO��7�D����&�g�R?��j�|_B��@AN�0��xP��Ձ����β�d�$�5�{#Z�n*Q�cԯO��8i���ʍ@n�p��[\��'>l5�ӥM��,
8��b�Sӛ"@cd�^�8���|�H��#�RLfn����5%�^�v�]ﾏ�2���N��[si��^��J�@|�wծ{5�BƨREm-�^A�R,v��_
�GNS�������8��_�v�&��-OM/z��w������o��A��Jޯ��P���G��/�X.dZ����ֶYD1��τ3;	nP.E�d͵���@������v#�=K��e�(���nފ�A�ɹ�z�y[^�H��gs���|�+���z�[ӣ;��d���7��]�I���a[�S�7�R��a��H��'�)�����N��[��tu���.�vegg"����!���O�Z*I�zގs��`p
ܡUv�J6",��κW=�6�c&��p�����Ҫ,첥���m��9�NVҸJ��� r��.Zx��!�����{8x�Wu��PQ��%/`�VV�%��"T��N�'�7ÌR[n�|������~
�{uS)�vU�y��Kp�8�b	[L�vp��A��X/����	9�m��i�Z����\�L��t�����ˡ�"z{O�ijp����.E���(T �,y'���rv@|���a'/�Gߏ8Qc�	{g��n������̎�*/v���Ce����$l(O�~��<�O����x�Su�
V��)�+���������� �JN�ɖ~�6�B��5�G���8�!yC�f��SQ�h(Z�T����-;�j9��7�l{3����*�Ϯ�>�q�ZB^�AQ��l���	L���ލ�ao��H�!oB�Y�t�JhoV����넕��q��ZbHk`H����09���~hz�d����$�>}��k�"�W2�> ��M�2�6L���qǤe��G�6=�y��}{Z1ٵ1��b����Ĳy>���쐓���wqq����f����c,!C��5�.��e-������<�+Y��dl�^z��892��KiE���6@g���Wfm*/X�H;�����
 �3�'�;�C6�������If����Ip�R����fa�ލ�����s�#�
�I��(�Xi�����_�eQ��"���ٍ�Y4�"�{�$�����3t5e���l�ӄ�dB�r��'|>�2܇��tZO����vUR*��I���͛� ���M�uq[$�yQ����k?x̋���bzGdA|�16Eԉ�M��3iQ����� ��_�硛]L����ʙu��B�ԟ[���]�����_�%ZI�U&|p]�b����<ؿ�3t��!�}��-�&��_�lǻ�:�.���RN�+���H��U��$Nu<���n	]M"xo������F��g-�������.�/l`�k9�ްz
��|3�9@�ft��r,"g�����w-�(�\d��|�hz����o������HU��T����[�u�i0��-;��p)�ߦ,������{K:��)^fh;7�>pTLE�a��>cR����>jԙ+�O��5XK�q`&�����9����?�^Y�8t���e���v��Cр������x�\�Ârl��G�H��C7��{�})A�y�Nթ�`S�ޭc���ǧ�V�;�3Ww��g��IH�P��/U���?��pNNn�m��+`:��芋��(�|�qʄ*�TS&$c��l�-6����2�>��vܪ��E|�`ٜ���i�2t�g��=|_CFT��7����F����l��c�/���|�O�����r*d���@�~��
dԍ�����h���̬���t�����3@�z�g�1�7�d�&�"o	Q�����v�=T����]U&�CMG)n��͆g���,����k@л,���M҇§ʍ ��+��o�L"�3������5 ���mn���!k�Ec�v�fV�4���/3�J7S7�~X�]h���?�Zj���Ju�n�:�R�6)��/'�mʲe��8��R�5�����O��U�%Z����~�RMW[�k�����n
ɝ���P�i��k��'Y��B������h�2���vhZ!�9�`lcq��9v�Z�V���~{����F͛k���8|�0��]��H*f��W���4t�+��	�;7I�{ER��ꛗ�R5���&-�����e�~ys�ڭ��P�U��M�e�I��V���}I�N�ѱ�KT�7j�Tc�%�w&:�ʨ!��8�#%:�����E<���_i�\8|-�@q7/v �$K�sI*3�?��2k�iP�T�m�BXO�njj|�-�?�z��.�7��Wa�i�so�u�n��@���`o��!9� Kl�=��ul/5吾���}��`v�^OK�ow$�ߕ�%�1qϛ���8��/_�7��7�^�L��x��΅{��zɖ�O�7�P\]s��u�V���;O4�z�%��fs��5[U#`��IĹ�Rzn�]R���a:����؝���9,M�j��i�Լ�P���t�e�˕���Eh���_κ_r���iZ?�4W�S���-3=�$dq�<3@���ΎӅ
�d�OG>��Z�&�:�z�+p�o��5�X���/Z%-z=q?��nq����DZ��B7�����G֙�6e+�@���j�z196��"P�B�����wm�a/�g3̮����g9�y��#.?3lrr^>��f���o �fWlDp��+����h�����L�%�n��:��%aNE	������j�(�D#������y$�1`"���7 ���>~�����)6�bnBo��/������bo!~��F�@7��z�wb�]�ٷ�ub����E��m�^lR'�,)�lr�� P�N7*b}�]�������[�	�E8 |�RL�,L���Q�,�bl��d�I����2å9�˲u4��� �-��C薕�p� ���r�1�}ʆ����ɢ���s�B��V�	���A$�$�q1����z1/ďQ��g ��h&H�ϐ�{����
��L�^D3����<��wǘw��e&��@v7aB�x��m��s���D���ٻ�O^�|[d�!�Z2|7BD;����V��|3\��#�F%'�u�8-k`]�e��ߕ�.>8��aN��1���xW�}7����*6�
U�P)�s*�1��58�+����ŨSŖ���QF"G٭<r	V��2#s��)ݰ�����[L��s�3��?����������m��!Q�h�$�r����<�������sT7���5��Ow�I|Ş�s�L%�w⣖���T��cf�x�3��+�<~_UZ)�_�/�zt�b���|�X���tѯ�i�h9���n����0������>��v���,�\�g���h�qT�mwo����=3��^�3��c��/Z�mS�mk��Ź��z����9=\c��+�q��
$4���Z� �ɭ�0�>�4� ,��)�Z-��@yv��|�n荎���4`�"�,�ħ��tɸ���Ġ�����M."��m����m��}��f2��o��>����P�g�鬪�.-z��t��~ΞO�Y�)��sH�x������d��T�<�x@�^Ui|�V��	ź�ȗFQ���3�t�@��ނYk���}[z(���k���M�zw�3�B��r�j�ܧ;�lw���sY�!N}ƭxʮV�R��:����e�Ta̻V��e��.i|�p#����s �f�dd��*&w�!Mg���l����}��T<��:d�%x?d�K�.��8/7��|��g}��g�\�6��Xq]K�5i��7T0�Ҟ+t�`Q�m�9����g3�� Y���n���A���{J>).���i�7ދ���C�;V�>X� v������Z�D[) q���w<�wy��52�]wf~����;��qVg�t��Z_�$����k�V[��1u�@�H�y���c+�����Ob��%B�wg�jΈ|UtY��t��D({=�	V���P�?k������u������1�X�[	���W3��
�O�<����4QRƵ�e�R@}�>�&��c7����X/
�H�*��C)F��Ύ�Lc��l�y>��"�n����t�a%\����x���ݮ�ݻ��5�Q�7�ݽ��<�}apf���>^��>����'/��s�|%��2O�߄[Xrd�a�7���K �I�;�`��y���x	���r�<M�p��2պЄGiP<�PP��T�Xj������Z�9�Vw��=J�y]��y-V�*����ur_�8)2���b7�D����\O��̹�w���PV�3�?#�bq�
X:��-����Q�ﻗŭ�ϚBݤ׃/.w�ݓ���e�1j�)X����vu�I�5%~�l�@���I��?��5t�j|@بa�8�@A�0��Jش�Vl ~�5���.���C�F��>�`-��Y�eߟn�cpf��>X&a��i��Ic�^�Y�]��T@=���	'�<����P;_x�L��lh8͋o����k�����Yj��e.�x���q��բ���& V��9�<hI�����M6�������i0�o���E�[8����=O��cz��C����v��j�"]O�<5
�\��(��B���dOJ�
4�0r�~�0i�����xi�C%^�U9>��/�^�Y��kٺ��H�%�A�)zuw[�C=�7`�=��;�eP=ja/�G�Ul��T"�iR��c
��TV���r�g%��s!��p�%�t0��d$��°�����-�d�*�������=��uu�H�&��P?w�t��6�kT�?@��R�vDH�{������8���9��冷�:m\(�@�?4�--�љ:Gg��ۍY�Q ���|��e�%ȮY�$%7K5�Q��Ke����ʙ���v< ;�ɸ�'�{s�!�P`����Ϋ��C�^�Ul�ԔO����2���*R�:���"����o@J�����Gg�n�U�Z4�%�v�жLͽ�O�SN�~ҡ��b��\r��ʈt��n�����d�UX���&�NX���w��T��b2T�X�Q?R�"�J9{AL^}�@�nfo���'/�σ�MM���/D�]G�qV�{��������\9�3��g ���U��gs(��Q��	X؈�k^tM����K�a:[`}\�c"p�^.�b��(%&ġЪu
��nO�7a��u�Z:�[mR�$�F���軄蝚��f�� ���:g;��	���P�]�J��z��橽-��_nSX��0��%P�,
'��پ�K��#�ًE��Bx"�"`X�(���?
����wy͞��%�[��fQ��I����n�nX�G�#�&/�?�n�=����#t[˔���U�M�AY�c@�+��U(B��P�d�t�g7��LC�����TvY�!��B�SҘ�F@��}���5�o��\�͘y�P�D�� Ƿ�`��+�[7|~$�NXظ;�߲� �*�G�>z ����("��.�k؉p��-����*���t����ށC�v<ē6TC��s'�IND xѠ����h�q �WI9�y�ݦ�E_P��l�U�i�Z���&;�(�"X@F3F�I�s�2����ݕC}{�.yu��"�ɍz}}�<q���s�֫L7��n�P�����s�W�5�R������^�ON6���B��1'�U2ӻ���-,�����^�7d�$�R9�w��{|�9!Sro��/z�H�Vi��E�*�ȣTf�d�<���� <@`�I��?ΰs�>�f'�
������v"E��D,�)|mU�����T��S��]rG,����7�e�N�d�,���EK�;�����-ܑ)��q�/�_ƛ�a(fŷ���4��g��҇?&-�b��$!}�Y�����!�	E�@j! ��٣LۊB���FJ��$�:(5D��lm�ƍ�X���bĘ�N���b@8��>�d{��!�^-W��!9��i1���ы�C�)�^B��}�:}P�
��X�+�J��.ƹ_d�D�/��{`����֙����	�.ŴIh�ZD>j*�����7-��$:đ_l6،X� �S�R�N)��	��{m���}�Hbaьߣ�-��ߪYF/��Lah�(�>iH�R椂��x�����5I"��.;P����r�e~�%`�i�~��4	����R�k*+�&��~g�_w�@��%���p��c ���lZ��K���{�Dgl��q႕C� �T`��^�����@E��,7�\��o]g>�K�?fF�8��2g�]h�`��{,��P��:8h��ijzZ�	���=.�v�5�	�E(T�C���j�MqZ��j��̞7�4�X��P����ooX٬�;�IA���M7��g���O��'��4(]�14�h� 9,�ssT��;I6j͢M���IN��kL!��2HTJ�1g�l��ʋ��kb2�K��ސ�[w�])R�d-�J���-��uޮ�"w�;�c�:��[��:��%��ݭ���D������I�<�F�)NՆ��EJ���(�����X���|�]J����i��Dr	։;��ðc�YS�P%|��әX�Oi��������������F�1U�|fծA�H&}{�eF��9��� �i��(��s���4�ޯH����[_��/B��9S�Oʲ[��8�E+�$�IH�N�u��lnW����*#���pΖ��6�K�����#�ࣦĀ��v*ƽJ�e�<Hz�����"qmw^�� .9���ΦU�m ���a�n?�| ���o4ܾ߲��d2�Ñ��qc�eb�~ā�I���XQFl�qB� 
5������8�^n�~�Z��"�*2�%��a�*��ׯ�����zG9��rj�dA�I����j�ì���ү��?㴺�H�d��rl��!�@^�}�ZL��a9�B�n�������, Q[�S?�>�P�Pc �f�>���N#z�$݄H��L�|�	��?���,m�[;.u�b[���ٸTߠ��I�,(��]3AҾq��NW-PTh��e��ϱ&��ND͔Џo��ޖ"�B�b�WF\�1X����u>���/ƹ�k��R��M�,�c���[�p܌e�]���¬���y�U����sX����|��T���G��*U)&N�*���,fFG����X�|_h��� O���l���qGD�x�U��X�
�6�u���t-O.�c<L��)�@k�������S�k�j�Lv�CC��j�uN�BU<�$�/�����`]��DܷVLC��9[0�h�;2���g��l��5�@�NO/.^N�D=~��t6�dO��0Cߗ��R0�����/��! w��i@��d�
z��b�j�z.?�A;��%�l���ޯ��aV�}Чښ }�Grُߍ}}�,8�=m��=��K����no]�\[�>"�lw?]d�о�ߨ�:E�\8�$s�p����<ii:K��^ �������3'����o�p���D�}�)?�|9��'^�d�1X�[x��Oo��R{��@#����7)��8�D�t����i�d�	����2v[�ݩ��=����R7��Q޿�Wxn����򽟢�QӍ�P���V�S2�P��H�G��J=	]��i5{��!l
�x�$pu�7�䊘iE��n��M_-!3xGL�{��6{x�~�����s����MmeP�ɤ�n�6����k!�X��JfEd&����k�2� ��
����٥��C).۔�����?��خ�#T����I�E�&w7�H�
�i��:�����o,X��`�\H�9�'S��$��
p-04���j$
��ݚ�f{P�E���W�{:�w���F ��#Ce�M��0�^�8�~�p�F��)_E�S�H��t���ws���R쎭�������X:���vPyoM~���XR�Mҡ�޺���uFF�V��D�ѯk��Ѳy�~J����.]��.�S�s8�hɃ��ǲu]g�"*kw&�s���!�E��| Lt�Z��<� ��Ώ�FEm����c���_�M���|������z�#(Æ��'��jݐ޲�]K�e��i��<�C��h�h���X �+D�V`i?���:~ �O��*���7��V�v8-�煮2$���ݟ��L�� h�x�$J,.��4�"7�mȻ��D�?5�Q���HSr��T B�ݣ6�X��	:΂�5}���`!s��v gʤm�m�����L!�\������7J��o�X\�b��2�L�bi�%R�Z��f�^�/�D��jTL��>��S5d;���|��G��ES޸�D���J�۷�)�P���%�bI�p>�`մک�
#��I�8	�	�ЄQ��OJ�Y�,�/�4�
��f%�k��y�Z/��A�O�'~}��8��ڸ��
B�G��}T���~Ҹ(��FJ���5xx;g,@� ?����T�=�q��n�1z&"�#Ч1P��W>M�/�P�Ӱ�)�3-H�G�uf��)<�c{
Ghf:��ȿi��ٶ���K�:O��Y��'�)Dq�0N�=�E�?	�%��D�؟�����h5�xBj��	�*[T������XS���{�(���j ���}���sp�WM��� ��<�����t+��)`�I����1��|̧##�ܬ�����|�$2oI�L���L=Bg*@̮�q�O�Ty��*_(9=g/d_?�E;�/��LZ�����z��LH�]p�^v#>�2o�`�x�Fo��hD�ڴ�?F�m�v�%���"���7�s�
DJ��W�f��~�FR���$o�J$�7B�D�Q����*@�%�g	f8��w�`�1h���TNf�.��[� ~��ӡ�� �J��<��0R0�bS�z
7���n��e&$t�T�Oӄ��P���3-*pb��En�ju�t$$0f�M�I�mS��3�3���-D����2�t�p ��t���9�v�@U��9̯ˮ�%Bd� �M�!a�4��P'�ר���s���9> }	*���E3"LO��(g8]܅���������2l����!�5^�Ϝ��R{y��s����Nɖ^�M�t@q���Ĺ�d#�T��ƻ�c���0�obBჯ�~{�����.;Ӡ�;2O,l�ʐ����������"�xc]')�U�cu�,��bت�v���gia��>&ٳ@�����a�AB��}.�'��p}.fg>�3L���O�u���/ �&��;ޞ��V���q��U�f��-my���$t���b�3��t7�j��#����M����&!����1Н�TV��1����K�`7�=��T>L���9t��'e
���B��A���2���Pv>����I�,`�� #2�D����#�z���&�^�-]��|����O����gu��ch%�.��1�\]�$�\�e�ZN���υ�q���ۻ�d�*�n<m�1Q"Q�#��u5_K����:3!��Uy}eO	�ӯ5 xՁ�M����=]1�9j�@n%$�M]��ɽG����7�&1a�Qg&�x�%�.F�NRu4�yqI�\3�c�-� ��t��6�`ǫ�
0�ÿ���n6a�b�@}$W�W�f�AY�$��N 	��CJ"��/5���
���!MSѻ�W!�� @�F��:��|�[���|2զ�6f���]r���i�D�'w��fe�K�����^��-�!�βȁ B�\��*r�ut�fZ� �b���ں4*���(j<��N��P�&g r�JT[���g�����B>����tk�L����>Zo����0Cݓ�. ��-��`a(4�����T�C�Sg#_�6�e2i%��t�Q
��haS�Z�G1�5_Gr9�k��+==�O��]'l6�@�o�ıN��i�ݍ��1�m���8b�P ǩ�����
ÿ�O���`�����`H�Q��&���~�*�;���O�8H:ȁ�7_�~�+���8̆:�!'���Y�q��t�dT^���+<yk��Q`���=�v~��Ab�U��}���A�6���RlbH�{��=���ٱB�J&����ן'�v�9A÷��,�� ��~�z'p7gw���h��\)�7k��+��'���%��J�	�|�L���6�9�� O���~ޝ(JG�El	Xr���QYP�a�R.��#ϸq��D�h�mk���7��R�]�Ӓ[*�7ϑD��R[@���1�F`����9Ӎb1q�"�F$8<��
]
���EU!o����8�w���UN��i���8����Ɩ駞�M����+����:yP�4�����UX��1gŋ��_ix\haU���X9� ��z@3�޼H?���c �M��GAz,FM�KDBP�9T�w��8!J�jf(e��
:��u�XRrS�I'@��۔�6$鐇5�a�k`7����o�tmJ*Qd�u�b�EdKB`K=���` ��wY�����Tp[��;(b*����{'k��	��L�B����"|^G��.��
�C���Z����&��;PVVI�%��?ݶ���yaf�"DU�Q/�84aX�Ab��E�����yE�@��Fd��A�	����"�bl;K���b|�'�6�	h\��E�@��Xd~�\b�Yk�����z�,6��~Ŏ�柃 ��m"
�
�;���y���`� ��ʆi����K�D�"f�k��}��Od���a�9Q9��P�X������{$�O.�,����k�j
M#���(@�_�R���>����a܃V�������O2��	�͡����] �� ��Z�rXʿm�.a��DiN�e�v��anԑ��M\&��|`Q{_�*p�`���'Y�+��-�H�f�Ɠ�uC�II�� (G=�<�0%�/�j��f��e�������P^cc��_�V�{�.:�G�n~��Zq�8��?����re��%`�5D��`A�s�f��O�cAfE� e���f�9P�᣽3�5߀Vq�ƾ��4�EϺ��������D�]��;M`F�n@>0ǂf�4|�o]��*�2�L$��ɽ�rr4�>&{Q��_�qp6�y�`��D�F�~�NGJ:�E%$m�.��F���2_>�+	͟L�o��qU�J���D�h�2;z"��� �7�L��z|�G+�6�������x��D)%��b�I���Y
��o�'�������ƒ{��或/3� r	1U�h 2���=�7��=�Gu"��(so��J&���\|8a��������=�J�
2�w�)�j�`��\�Q[R@�`S|B4�����
�k��]��%��2��K4E� ��}�6K�F�J:M����>���k�6b<H�̩d��3Rg�����I���$]4�?'m���Ue	�Z}-����Q2?��cD��R������a����:I�-�֕����^��P�~`�V6"-N��ȸ�e�&�T6�t�
��%��vւ�i�`���xݾK��/K/���X���1������w"
���G��0�|�p��p��7g)�T{�\i�G�Ư�bc����8��Ѷ>bS�qc��!����_�=���s.٣©�*:�zK�"�ܽ�׋�o��elOq�������ҡ�򪝎\F�X"[�Tg�?B���pa6�2�b���Ŭrmn�O�
��Z��qHオ���',`�{?�0��]H[�:}dҿ�[��������9wu����wJy�8��=H�5�z��-h���=�3h�A���;ҽ�]DN��?	P���6l�[��a�;�xKɒGG�
��>9>th�yot!�T�`P`^��#{2����.P��n}8G���̌+�����MzW��9�4?�;K{�-�g$��+�y[!�Has���E||�_D�B�<o�I��C3.{���4b'��,�8��8Y]�|ʑ���~~���j��Ü�x�����0��Wh�xө��`IdXslL��v��t��Xn�j���Aȷ��=Db	o�ֽy�G��՘+��	a��DD^��1��W����~�3E��4���--[��X��bQ��u�����&��U�H{a23�
�P9��4S��i^�v�R�/dO�|#\�$�V{U����i�i4H��Q��hGS��@���<T}7%2=�eq� F�N�W�6�p�0u���+���og���pu�B,g���O������ XK��L�d�]�i�8�b�F��+Mu�W�6`��h�֯�Y�!_��\>�͝���I��o��Al�_PI��xK���3퇂;
�� ���z�Ņ����G:2�H��d.z�D�4 ��W�
2�̭�S���z�e��Ce�����1h��q��ۍ��u9�N����N�������+��o��`#�m��3P֍eNI�`*��䊾09C�U��ŷ ��u�2[�f�l�3���[x�ԃp=���{�.�e׵-�|���Y�!��e����]�'���=:�`:���5����k��V:�5{���*F���t-`��eaY�*n"��"jkw*�Cֿ��^�d�<A�Hw�&)*}�_.^�j��PD���c� �hj��?�F�܄ݱ��S4wʤ�k�m���<��r,���>J�ƀ�����:5��؂��:��}%��Q��r�ޱ-�cNB����6��_����b�O����&,%�fl?�v|e=c'(j�^k5%���DϬ�ܣC�r�M���!#L���z�3��a��a��!`�m�L�R��v�l[hZ�ÌB	y���vwC��(�����=�.i{���v\!W����u9��jPX�cw�OY�w'��}��V���#� ��;۵3��J���ɤ�T�M6�mA�F�ֵߗ�v@�I-�f��b�2����z���M!Z������y��Z�1X�`K(�Z�0�@�w��-V��d)�<H�ӧ�(ں�v����'{Oמ�Z�n��1��V�a3�#�l�;{��kO>oѳ-���;}enh`���Ə�1��k���K�t@Q ��sx�~���C(�`k��
ZS�k� �$d8��S\4�J
{���=q���Au�L�X�]�$��þ_���44Jy�a^��b�IQ�-\��&����RnP�eNh0�~��RH6I�x+U��b�\*�@��K�9��!I5�o����R(v�J:)��\�v_g��Kh,$��R��+O"[����#�`j[E,
}3;IE� 7�*�6S�i��]���
��W;�N��R[U�lQU�_���8T��pngq�:]KD���"�?z�6.kW��T��&q�אۻ��.=�4n�C~�)
��DB?VU�n�m$G"��u�2=�LQV�gh�N �g�B<�����ˇ��9�z̭;!*���SvIp�V��Is}��g�.�nJ����U�F�`�<㞢sU�����)�S�(u'�c�H��A�K�h�B8*	j�z�	z�
'���u��
�ỵ�V�:�DI������p�'���s8�b@��	v�u�ťKҚ����V������=C�-e��N�-���}<F���-�>4tp��-`�[n8�c��_M�	v2;y�D�,-b���)2Uz�rn_K@8
t_R\�_��8���+�`��`&1]����g,D���o�<��%Q�9�%7�%Go��$3zk�c��奊Y�R�� ���I]N�H�M@��זn�_K��{Ҭ�/����[0��;�G�-m�~%�P���J;Sݟo�wP)u8ϥ�z��l��0ɜT�`}?�FUG�8�=�\Г��C�~3���>纁�a#�Dyu�e7���d���j��\=Tf�&��K�SZ�Ɏ`���a�"��P��'45A%Yۘp��Bo��N�f
��ն�^%[����wk@���Y����q��ѥ'e;��^��6]jq�g{ 8���‐S�&��%�5	��fʌ�X�d�������UK��CI4�îvẀ�	%lKݯP��D-P��Wf����GZ�˖%�=g��%�-��Xr{�^hK�VI͇����G-I+�_��8�Pj�0t�~ �m^�D䱯.�?�XN�U	��'��i4g��Q���c��j���ޔH=��]��^5D\�A�K@s
��-�n@^��
�2�[�:9snu!8�T���(�����H?H�v37P�a�{�3���z�*StT� "훽8'H���:�mqE�^j*{l��&�'���a4�A���7^^I�����`멜S>����f{��{�٘v�ZZ�Ǎq��L^ۮ��g?��I9�i9 ������o�om��`G��\�������b3�)q��u«NBP�:�d�6 Zo�*%���wڤ�&��&���ý�8�j�+wl����N$<�%����-/J��"��}��'�g��Y��~����!�$3�k����u�5&�t`�&��V �z���\����~
X�B��Pv@p���N��lS����.�k�\X2��U̫h��5�~�|?��o��7�b�^)c?oX�W��}�G<�U, ��l� �;�����$���Í�0��*7���;�L�9��N���t8��w��^M�����Y���]�f���z�AS��֑���W�b}��� (��@�:��La<c ���vo�a���i��L|�Ui�1c�`r9�1�5el[�I�s�a�U"���#w
�qP��
��6�2��du?h�S�A�
w���� ,����MtH`�; t�K���D<���3���׊��N0�-O��$��\fwH��P�B�'�Ã�f
���P+Y����s������-Q�K���@y���(�!H��L��uA�|�NuŦ���p_�rX	��U��n	�� ��WP&����m�@�a�������@�;W_,�zt�7��7������a���O����;�% r�O���Ђ��\���,�G��4^c/
�R�-S�� \J��vY�i�$P�Z�w�N��S|�BTD>mP���pT���\</���M
��qD%ᮬg�C�s�Ⲫ5=�n��u��E��M�M��g�M���v��b��x�2s�M�}�
��vGi�KRa}����;���M�G�Ѿ�<��Wjȸu�� t?h$�;πK��)�g�_!���=^Y���ֳ;B.�Ly����7�����f� ⍭)�����D�w݁���k�� �ۺ/Ht|^oC�t���򕌻{��{�VZ�~�e�)06w��z������fD�)�ϑ&�B*���x�#����������uW�4�mP����h�ڈʔՍ�������O��1?�@��m�����Oqۣg7:T)��������K
��ʮp�ܚ1O���M,���˹��Dn.���!]W�Ө�G%���:,��Jl]d"��Q����<���j��B�<��`x�PZV��f�� �IW�����ӂƵ������zt뿤�%}�uS{���Z?�݈NRQ�H�����b��&�W��Tb���|�dܭ�;�;�qU,�VPK�^������S'@�֎J�%�l����/�m bbQw�넧�ϭ�~ᇽ�-���X�_T�Ӵ�i$��RǛXLд����,Qx2z��-^��?����_���Uۍ�h$��.�I:js-?:>Ls�J�y�h��+x��6q��b�?�K��$�
ťTk��\R��:P��č�pX~��V����f�D��F=<H2�ۅH�L5=���n9f�eS��B76s��i�-��X��[B�����bs���u�x�c��nm�,����V�]����영Nb��1�ZŃ}9��ڟG 󵚥���0ԩぴy&����?k&1��?U�}����Z_��v�������L��'�嬔dHf3>nv�^%�Md�2�2}��4��p9�x/��q�eg1Ym�YX�=2����qb܏%��*�KCCu�&�9쏉�� �ۤrG�H�+���-�(}w㒪��Ĳ���Q	v`ij[^�g]�� d�y�o&�����ub�W)�%J���2s����)z��s�*�S0��W�<3�����\`Kw��q�J\F����]�o�ג���Yų��뻇��w]l�~7ch���$\cB��W@A	��K��f�3��r���yKMR��=�Zu�E��v�C��{��幞���>;�X-*��Hz*��r'�o���287��g顿�����p[��IM�+�!�;#i�%��,E��I�����j���s�6�w�;�{,��}�������?�e-�y�n�dp���#�Թ��jb�OW����w`-Q�j[	�S�e)��Ph��s�A�s�W���z������u����\a�ҙ��K+�J$y��M�~E���'�`����3��Y5�լ+�w��;1�� $�ق�p�]���ݽ��fC\#���Ϲ
(���+Tևڥ�w���'/a���iR����]���V<P���{?�7+��aVs�׼�$}����Yw�m=a<�L|���>���*(�g��<d���^k܄��{-llE�U>�GLR�� z%9;P'z�G�YF�S�n[#�d����]��׍V��`Q&�[}[����s����9i�Ѷ=f핽����4�q��������33�xC��Ps���o�ՎZi�حng�q�d+�&ƀ����LU��]����d�T��!�)��fef~R3X���-TGo��8�=ʇT�G��tn��O-x�B�r|�m'���DHٔifpG�rf�Í�π5�qv{I�!J�9T��KE�\��+�k+Ʃ��O%+b�
���q[�r�xB�\z�_π��1�T>+U�D�� ���J���i���Nm�jo��m?Iqg�, O\���ki��!�~j#�>0A}��u.�|��ĝsS��T���	�;Ol���I�/0燛��E������x��7�so��[��VTJJ��P2��m�PIȘB�1dO?E7�.�2V�̉�1���J(2�$�1�޵�^�{?���������g}���}�����*_�� 3���v'�˘�Ï@��}}1�����[o	w�ybG>
�+��z���2FTCދ0c�����6>{� s;|�{d���*+]�ٝH�]��<i0E���~��F��Č����fOl;�����%�ڿ13,�㬿�(.MƖ ���>KH���0ad�J%����B�녧�~ �o}k�7�_;-r��O�nJ��b�v��`����|�P`:a,� �x��Ir4��,Y����%Z�N}}��B��r�O7 X�Z����IL,#X4���6|��U��f��	�7��iH2$�lqX��K�"��%�STJ���T�+�뛋ϸ���V;b-���%�j�~t(,�B�������v	Pw)�BUװ��i�S�!�Yl�;����e���R4�G�s����R&���A��)�"S\�	�;��T����mT@Hqi�y�ga��:��&��,�z�
�zJ^���{tF�
<�?��"��/gO����w��xU�Y��#�bi����^�84�+����~Ք}(�O���@���ҹ�͏bJ�re�UJ/�q��8��w�H5 c%�8��	�u44��Xu��!#\QRH�8٣�̕Zc��S%��|�ٗg	��p�p=��1��롊J2�}�Gkp�N���O3�l�T�ʴ<'<Ɩ��6$��'x�pUZ�<���Aȹ�|�f�����E��s2k�H�R#@R��A��S���ւ��[��\��Kq$���)�����xH�uvV֠U)b����k�7r��[ ��S�>1렔}�ίn�8���= ��U0$�w����"���*7� t��v���O* .��7��N�8g,��7R��̯?�A���c	t �"u^\U�ʲ׽��w&�rIي��^O�[��m��.�j0�V�m���圣���,�7�4~8��~RS��'A�tv)�J�; �Ȉ}�>Tx���{�z���p�n�b2������V)��V)8L�m[eoo�G��KJD�?�v��5?��˫�I?��R|�#�����Τ�?i����+#�{)�t��/L%<8C��Ɲ�/��6k#5�4v�2q
=���l�uo�/L9�b[e�����̯z�ƀG��Є����d�NԸ[��6�Wӧ���{[�L���5�n�1�U6 V�|p�X�⾆���Θ�#������D�#�p�O<����5�E|1~��ͱ+�7�^?�EX/��ǿ�U�-�4-��0�aS3�@��ӧ�+�$�
e�I����U'�U!jqj]2nݭ�m#+�����c�4�Fs���ރ���e�$��^�x9��*UF�韍����Mw35�,U��r$����)-�Y�p#���{�u�K�,t5>�M[����^ԑ�{��a�z��N5���s���x5�q�><��68/��E��F?�oߦ�	�Ur]�}�\�UO_E5X�-Y�f����}Ʌ~���J bo��(��DD�7�뢈m
#3'y�B�J�I�9C��Dr�l�s^�0棹�{U��0�wDzM��� �< ������u����v;旳oߴ��vϖGj��=v_�����NKň���$oϗÐ �ג.���!R7D� C��ex�ǿa�p��z��yfr�*���`k�}V��N������Gtoh���-`���%�N/���4��_��K��/�^.s�耕���%��hu�I�X��nL�u���g�6�R,�>�{԰�.�1�;�4�d�Q�]:�0?��� #u�_�v��m�I/~��DaER]%�A.��υj�O�ֲK�>s�ݛUU������77�Ϥ�uț�?'��<
�j� ���%�G��]���t.��ːܮ�^�fߛu����ԩ]�!��~QI/Ĵ"�ވ;Ʒ�rD��\|G�V����?_V~�w5(���k	���_����c�����������~�ߏ���?�����~�z���F��ܲ��}5����{�	x�?��d<F���"Աd������QgϜ�����=Q7r_'����^k��b@��]Zk3$�m���`PǨ��$��B�4_Y;$��,MS��rjω+{&�"�M$��c/i�y��D�vy���oX��b)>�48b��k꽋Pӂϻz'+8��/���z̎��>\���Q���?�Y,H��@VBM�A�⧭wE��L���O��61�;��sF*<2�\���.��,��#�5N9S{F0#L��O�ч����|�9!���_[(C�;f~o���X��͏.���`���7�@�{~#��M��kpKt�u����Tǵ��Ϩ�*�^��DiE�%y��fGJ�-�6~�&r����=ﱥț��r�����,�y���;�	2��������71	�\hLa�/��&.�>Pݑh_*r��m�M)��k^���"rY�J������-bm\�������hB����\TQ.fJ���ٴ�/]�2�/�_�W��v�\���C{|+��R�H��ZΔ�������zXLaޱj�?<�s���/)��X�}ؓ����	^̮rQf��k	�����}�/<�4�i����_���B7�j�0)�Oo���/A�af4^|����욯ƕ��W�8���Q��U�r�]�{�U���Tj�8W�>�^�]�Z��p�3��?�͸�9vL��#h�-u2�W�
m��l��G�fv�;�\lx�O�o�L�������W��G����n$�F5��qa���W6�J�:��m�ae��t���u�r�� 0�8�t��s�^L��@l��u�u�:��.�&7�z��A��a��/�z����h��܌n�>�!���eei"5��C��[3dQ�`��o/���2�X���g�]�2\���N�;`�5��Sȓ+PL�cT�G{G���2+i��d�`�������?.�W}�f��(�b��r���Ć����.�	�����5r�~�ƭ��T��]#��:u1��Z������+wjB�L��].v)%=�&�C;8�U�e>tG/|e�Qs�rًS�T=\>��Z<�"����/�4j�"���Z��t���S<�%#�D��q�j��>]���Z�A��'�C��%�h���(�����$kQ��� �D���&�~�`��&-]#��\HG���l�[��4��Ы7a�o��m+!�x�Ջ��N�&����4h��Q�"��j�W9_�ӶR;a.�Y��ġnZok��W]nl 
#_��%�fT@SUw{���e���*x�gZ(�f����
f�e��5-��?�I��L䉔5z�����fx�R�KZ����x�)l��5���� 
�WjS{a�_�O���ܛ�;���S{�#�qD͞į�I5oe��r3�֪���8�l�]�cba+���B?XM�'f�vLˉD�0̅[�9�]58/K�ay�E���,�j�U���f@��Q�-?Ř+ze�6��q[�?|��/R5���EC�/��-��� �2� C|JBw=����vls6��$��԰<x�.E`��I	�}`4ou9#�ί��o\�K̼��D��'�m�X���&#��8��C^N~f{�\��Q�,	m�}-ݮ��=��z�T޲��$["�=�r���Z+���y��%��Cͽ�-Z�J��Iz��ݦ�H��%�ư��.�8����e�l9��"sS nQ�i�Bw�h�ё����㱘�_?���P���q�� �o��iZU��rގ��n±`� �o��Py_R�9�'|<��@D�	����O�����r�'�6Pِ��ˌ��n6�ij*7�7lpBȾC�ø?L�:O~�8�r&	Rzb�q};hԝ��bq6E��K����7�f���n���E�4Ʃ�FQVsaL�t�v|�j8=� t�q-3����m�h���N�\�z�\���t���7Y�����6�Ӵ
��@1�NO^�|ޝX����a�Y	�/���] �M���	��w���7��5��6�¿�9��o��7���ݒ�1��uMQ7^��^������/�in�>��>�Z�?�^���0�}P�n������/�����)R����m��k�6����H��<\�� ���x}{E�iL �XP�9ܥ�S�:��w�V>c��BU��7-_��Y�ϧ�ǅ���? y����~�� E�;�6@/Tyf=�?:Tje\��������謊�$��<�Ǭ��������G�Sc??Q�6���?B`�C�D��pg���q2l��.�~��2���%��{h�(4JB��(�{YF����J/S����r��w�@]��z��1]]�\��1g��h�e��Bb��փ�!��?/�v^�6��i�A�[�V����/5�0+o���v������gJ��W�B���N�8+���(S"�s|_0��+W��g����n�z9g⫓�Q�~ʄs��d{MB�-\��B��K�MW<�U�b�Ɓ/a��{�D�h�iQr����b��\�B�\�B$���D1��Q�� N��et_.1���_Hjۮ�3�zq:�]��l�v���xܷ͋(B�r�����,d|�A�T����emw�B#��8��!SGm�U%��R�#�8��)����q[�S�n�-�.��\��[s��ͭb�& �ҍa�5쩢B��1�}�\dzx����������&�·���ޑ���Z���1|͋1��2U�!f��)�����G{"�����DP��;��!�~V�eum|'��4�3�%\���co?;�Z���Y!�;�t p;p������O�!�

3}�P�n����/WU�E�i.(��n� �J�c$��Z��Z,�mw?�A�j�<���r�\�ǂ�NݵP���bx�j��v2�N�*�����0��:����d���@���j��.������󮓍7���Є�>�I{�r�g��q�&��K�}�m㋑0��6�Y]�^^sã�% ���<ئf����!�#P̓]!�%5�d	��B0�bDA�g�E5�=[�۶m����G0A��HO�P��'�O���e@��<��&j\/��#L6Z�h�vt:�#+�o*Y��ǣ�>��ͷ�5]�A����]�75�r5]�#<7>Xδ���	���mkZz�o��&��w�XZV��K�D������8���P��D��ti��RU�d�gM������z��W�d&�)]�N�_�O�"�ޞn�T�*������A���8���]Z3SF+�~�-�p��6S��S��^@�1�w�?�]Z�YPu��3?oR{���'�i�ԏ��m-�:�:���Q�����,����e�J'R]�^���s�"���PI�x`�o�S��	�\�I��eX��)�(y�}��#�Ȧ�Ar���.��$O4�w��"b7\#�����u��G�bXWi3���IQo:�r�c�b��1�84=�H�r�[�#p��e�� ��3�{ŃF�1�]f��� ��KD����Q^+;��9�~��&�U.�W�b�\��0�M�%�z��X�;u���p�惤��MZn�Q�2�ۤ�t���4��!>�pi���vm�MѰ��@�m�okT������y�>&��%�1A[ZA����v��qW�����6ǽ�d�H8s�NT���J6W�+w��1�R�d{:�$9���x�K��/8��ZV��{��Ymz&]'�sk�Lȁ��������t�t`Ya9��1c�<�a�*� ��M�-���sig��Ʒ�Ąw9;��H7�]�=YI���t�E?���J+��׼�r�ϟ,�t1�J�	ty�_ENI��z�x0�Ct>մE�,�P��i�["��xX?I���d�`��6_�������K�������?��1�b;Y_��6�okoh����oQ^�V`����1��e���Ԫ[��]%vXhCy��z�{@�l�ʹNUb���K�p�����oZ�E�Z�f�V�n���+�J)������
6�sl�8�㻣�l&�쉣�!gC���q:��W?��0V5�W������E"7+����
�Cb� ���,�9mR�[���ݲ{�o�7e�^�ͤ�(��d��!_/N�&׬c�&٦��3�*�M&Q�'l������C�w�n�TG��1q��5���DM�y��5f0i�� ׳��1�,���Q�
�_��4�F���~c����\����6>;m�i���6Fo�SC��	I������yե0�`���;��4=���HЀ��9�#1���/!�w=��`{.��n &*�/��U2���Ӱ3ig7b��گXb�bc�����V���%{�cD,8#>	|�(Ӏ��՘r��aʟk���4�n��s���C�Z��1�ˣt��S:zl|t�m���ʵ>�@ڐЦ���M�P�7������{�m�ct���>B�%�ٴ�.g��h� ޔ�ؼl[}����2�0e�O��fw�ϥ����9� cV�E&�>�x�-nߍׅ�h%�
 ��a�ܬ�E/���Maʒcv`yG�-'�`�Lq�̮1yU�<$���&o�(�΅�� ���-��$�%�N%G9'C�`-������Y��.��ECp������8����U�?��nw��d��
�����Jx�C�{B��e6>xTM�/��߾�0�M��p�K�Ʀ���n� o>�ax�~��ݔb����=����<�� ؼQO��=+qs�Yk%hg�R�����l,S�b��o�U�<\����o��S��ȟ��M�-hq�l��ܴLL�R��X�][A���B+<�����Vc��5�,��h۝`#i_T���AGK��Vt��}��{�rtDBR�$;%��衏��� �a�5ϛӼ��j�;��;�abp�A�V���~�������-��	L��Z]%^/Z�\�*��Z�x�~M���y�@��1np���$���0%�5�������]���?'���f�%�7��z�ѳX�o�q�F���I�o@f϶�;�q VU�@��]��nPu_�@\�'WE/&���}�5ƃ�+pL��'�B��2�����r������;���N�a�&6Uq�{�m?�o{uDɳ�|���tzL��苨82+o�v�Baoz�`�@�� u�0���b��W�z��D���U���'"9�w�[ԫ�.Nq���di������d�2[�Nnƽ#,�̲*C1ꃄ�o��;�����0�'�݄��ԝ\`Ru�E7�m�"e#].�{[$�O�eMg�MQ?�Sv;\�j�dP������2�*y]�	Rɍ�Ó�	I�X��"�s?�7����o��F�v]�����y��}���fc?5�<K`�{�
�d�HӁ��e]�&A 1��#=�o	��(���`�3����Y��1�Y
4ܰw�T9_�H��ݍ10\����%vPo.an���D�NƃӍ���I�E��5Ly�!a�
rVL�^�Hvx��J%S�����)RHy�܌�����)q�}�"*�M������j*Y�?^�%�]�v~^� �~��i�P�V9�\�ĜxM�{;[�2Q2�Q�\ @R�^�e�g�U��jƱf�&�M���6nH�-��\�7㹊�$����ʲ��ɦ�b�=.��E�<1j��u}Co�E�X�����@��Et�7
C�4$�����u_�Z�&Z���	ZS�M�^��tQ;�Ά^ÿ��v�X���ޞ񂖋�$�Z3�ܰvv8r����'Ԏ���poJ��H��'.̺Be�����W�~5���>�H��\�d<H������� 8v#�AkH,o���D���#^����o`�O��Z�d�as��ôF5�ީ��.U� �vk`eBF]e�/?���7L9ɯEOQ2��]w�l�zE�%�MQW v�3��4�i�R���d
�e����[�p�|P��0���G��7�}���F;p�ob�ڍ�>%�V���ז��i;�ڇ�ə�%#ҬvH�����(>�v�l�O�f�{Q3��S�X++�� ���([2�����ؔ�Y��)���Z	U��٦�o���\^�p��p`��&���֍�2��:3%�V����Ԥ����!!���ۈ7C�e���F�����X��e8��f1d~핥s�J�i Jd6���(��L�C~�
�N�ץE�4���H���ca�$��8~�qri?�����<̚��1��K9ylh�)�&���h����O�*d�4��Yax�MC�
�mf �q��ݩ�;r��1�Hu���#�"��Q����KY�\�}%�}��.!xt+t�~6���!��-����J���.�Ƴ3�NTA\#�f�7:�����u�J6���8��纜��!����s�&��x?afDd�TFCN�#\ْ|�{���H���|����'jMO�5�Z+1�ؿe�j�Y}e�0nW�U��Ƌ�,�$�|�>�%�>�i#�>y)jn	�&��niN��iDhRX���� G.�����@tġ�G=./EqF��g,��*��ɍ@F/1�?W)/E4y��_C�0��w[��8���9��6�|-~��Z�EOh�*䔏�.�$:3$����C�$l�0[I�E�0�iI��n��Ʈxd'	�"3�k�h��ů�v����CMV���q-3g���	wbz�A|�8aj��KbX��2�=M\!�F�.p��pjA2b�(��FH�� M�~��k��^����%JJ� eС��[�)��5(S�mS�WZJJ�8���(���N4#ޜܾ���K�<��%`����Z+��#������`��3�af�zF�N��֋��q�,�[��H�Į�����bI7䮟FH�	C;���B%�4g����61D�Ǫ�w���clG$1ʼ}����&��\��d<r�A���!,�$$�F��ɷ7�v8X��:�E��ߚ1��U�*�!����]׀&�)�y<ćP2-�i�x('�GQu�F��w&&�0ٲ �t�e�����X,mKI��M�:��������'a���J]��(�8�O�-�+�o�����Z�R�/�`>d^#6;��+�]�|O|n�`��-��Er$��J��.:+������|b񚘿J��H�f�\H���b�r�J��]g���s�7+\ΦJZ�2e�oVR����7����`���c����c��ذP���Bt�n������~��n�C��G�v�N̦2mBp-} �����Ǳ/j � ��nݍ>�J�Ϙ��Q�j�!u_v}������ ���'�סX�)ȵ�M��O�N(>��j��e&�� ��e#+�ݴa�z���g�ŗ�Ѱ7Zg��2]@Ӥ��~���vπ!Dh$�'��3#�J]g���KV�H��ã��;�V^@MW`��3�5��~�	���x+����Ճ���X���(,��!�_����b�r}��Y�mr����d��-�F:�mA�Z�p���$yo���-QӢ~�`a�+?xǟ0 ���9�5P��j���y�a?�H=n x?|3_���rb%���e���`��\�#������G�f�24�$�a�ċᾀ,��pl�Q�j���"�v3�X�	����347��W�}�ي��s[��Ԛ��;�Q�XP�T�����cs{̴y	��:jqѳ5=^�rǁ��u��/w���p�����Ȍ� Pn!Z�7���W�يE�C�bEE�Ǽ�L#G�x��.=5�0�������%�~6먇����F�a9+ݼ>\ݓ���a��@eS�����<�2�Z�����¦cĳ �����q:'0h`���$�^�/ʼ���)��P��+��\��f>��-�*����̜s�H<�����'��`��"��^�S�1N�,"W7�E���`�	��X�2�*L�a�}���F�{�}��ZVe�_u=�
�g,���0�&��=e;��◗�P�H��3|�w��\�%
�bv�`J��^���`�2�A��֚�|�P�Ա:�a�8,
�]R:���&bUab�`]�ƶO�j-�=K1F���GB�qU#<�++E�*`pV��Q�5x�#dĵkq��p[	+�/ʮC%[T�˽QB���R���@�J	�ׇA��;�E	&��j�����6��H*8��Uݳ��<S��e��7��VĶJ-Ω��Aj�@�����5Q�tB�$c^t�@�hA��n�6���+���M��fk��(�H^�5��}C�l��7�� #�8���0rd.'ZF�K"��c$�����Lb��eՄ�E�� [a�k�}�}���z�x�|¤����1{�~���g?`�8���;�u"�> �q�N�0��t^��K���	B(��V�M�pR���I;:�j$9DO� ������xT�%Io��_䰼Z�xz��������)�E� ����\B�|	��" �@ ����7o�(I��g'y��6��m�1�vPe�\)�V��M�*H�Ы��z��^{oY 4�k���>��3��eYab�c9�����N拘���b��q��J:p	���wk�ܨ1D5�kw@��(��91%�z-/��F�Xo��1�>��5���F9�Zk`o�S��+<R�"ho�	?�
7,��Y�ȁ~'u��*r��
h�T����A��������h�+�^|S�D�e�W(�t�Q�0#�`q2�c��dNx�ؾ�x:�U�H��!Xh[ޛ��)r��~�I�`��2ў��
�jE7;�~��2��$o�ްP���f�|�S��w��
� �S���*̓>~���K,��2�&F�k@L�"������6Xc����ɲ`jڙ�G�'��D����ب41"X�6=��G%	ψ��`&��̤���/�"��&��v9�`����}B/� ��yQf"��6�7�����k�yyNs�]��G�n �\Zz�xO�'�yjl���
�'jί��Ѝ�cqF�Bl�;W:�ܛ@����b���F'��A�N�CkBq��8�Qö��0�ʒ�ѭ`ʅv���5|�>=�S$g8�a�&��=��>��S��퇸�1]|��M�X���ؠI��!XV7}���;D-i.qQF����wE��k�M1�oBya��}�
�c�BN�����̏�7��S��ߏ�W���}��V�|�W� CRl�j�V��'7�x�`uI�z��4*�Q����M�Y3�*,��B��Q��`��Լ��4Zz�ۤ�ˉOD��~Gt��eK��4�t�B(����]�o�rl�D�ƫ\M d��4��hg���!�_�@� ��i����G�e�ns��Ԉ�!�r��M*��t%1����;��J�O��J�:����M�w�/u̡�
f�Řo��_Ҟ4a��ꨍ���-��g��%h敿�̬�=��E&9 �� �JX����L��m�s�Kx��=�(��F� ��B2&���9W�ί�Κ�#ƃ7�m�>'3m6P�U�15?��`$_�mP����
��g�-[�"Ttb�t���+�����"C�k�1"��Y~_�'q�丶�7����F�<uv"5F�{HMx\�/u?_�l{�8��dXUk$��KG4w�q���j_@�/n������G���炣��w>�7�1����ݐ��V�jK�ܒ��Dy��sa��^em=eI��R����!�=+����+XV��췚[��q��l[h�4�䫊,�M*�o�[e�����{�ݟ'��Ow�GPuE�-%�)�,̝��EN�̰A;?���xJ�F�\qt����ϚL �J����o��a�NG�-a��c;�6�ǻ1������-�,�뺁1�F��g����^sK,}��t����n�H)��K�����e�a-?��0P�|�d�N{ؗ��"fv�X;x'���Ό�9α_��Zv#[8�{�K��l��}�Q5�(����t*�N�#�a>3e��e�ߙ�64;6��K��Ʊﮊy�D?�Y1=��3�4�V df6�0}f�7g�Ydۛ7=<���h���a���w�:�S�B�@��p�l��q���&����*����h�����q����)��������6��(%²V2(r�8.SxЂ��4z?o�Y��p}�`E�Κ�����S����h�^��ͳ��3f:�\��BG{:�U*��{����_9ƍ�b�f�P��
ռ�`�D��ݿC��U����B���K�b�Z~Rq25��7���zF�C/d�sU|y�Iք+PHD@���f&��ۯ_�ꚒEǰ��4�?X�{z&L���1�ì0/�y��T+��;����j�KD@�څ����X
�fz��J�n)�~���=�YhG6!�(�d��]z8kz�x��.s�����.-� y�X��t�L���,���D*ϴ}�x)#4,u��(�TyQ���x��q���7����ǕE���uVNuN�X������Co��- #��#���#? �A��q�eH���Z����Z�P8aέ����2�NAs�_�j�_g;xK_���{��/����/c�ª�ݠ/5;�2X�����tߡ;�|)�N���w�S
oJwD4:�rTfN|�E��5B�WT�<ؙ������X'���ΓE��n�
i��k��#��Æ"zsw]����/�<�s� ����([����f�p�ه&g/�ȇ�A[E1�>w�[8p�}�l���3N-"y�t'߅��_��x�ܨ���M�e�i�����8�E����j��%u<�ͻ_��?���L�k�С���;�J�6/���0^����7�'~s�a��v�~x�O֤�[�GV�e�7g�^�ΛG����MᎰ��Ǆ߬�����U�%����W��o7���Pp��'w'�d�j����o%3���dl��+�3����vr�D'��Q�{��)׎q&��H|�t�7�I�.�dw���RvQmyd�p~���s_Ů���w�s�t�����]s����v�
�=�B�!St��Š��?뙴���z����i�u��d�lNM �-���T:�x��-�yBc󏞚�ޯeT=�VWUUj��?ک�5��3'f����9o�@�!�_v<4���n뜥I��g�5��B<��^l�J���j�gP*�J��^�5�!N	"���u�Ӝ����������z�w�1��e��n�E1|)�U})o�s���qZ�l4شR���d��~�/�0X��,�D�i�u��F�]�Q��F�#�YĜ�%�&�����P��O홟�����t�wt޻�f
�Ea�ofEv������T��%�c���:{���Έ8ģ[����ךª��J��rL�+�N���Z
\ԉ@�F��}��)k;b�t����wz�.�4$?)��<��ɻ����w
o>�jѹ)=&m�1�S4m��~�%@:AD,˫dc�����Zz��-��^f
�I�d�����FX�YS/!H���;eg��Ɨ���Kۃ�~B�P|݌o�2�_�lKCy���s����]��X�Z�W�����C:�t���҃�d0�
�b�.N�=�I��fzk���5��\�B4��r�8s�e,�$^����l;wYTHPtX8�CE���e����,�6n*8}뉟G�tJS�0��]�[1|T��YOu��f`�˗e
="w�e]�w_�B��5�|�v�Ts!����F����">x7��dP���PG��4�6��4+�69�'{M�s9g����݂�a���ԂN����t9-�|S��L&����ҁ��j����3�O��q�����r�)kl������-�]��J,����ٱO�I���{��p�	�$u7X�:���
�W>��m����m�"��Q���ck�a9�V��Y 6Yl�s��=~�b�a�oS}�yƪ�ƌw�Y����NU�0��5�
Pex�S�C�i��G$�����;eş2ݓW�c&���.�6k��I����s�%��z���zs��X�"�Dq�:\��(���a���3�\��0�,�:V��p7�XK�_�<��U���F"��mb�T�tT���>1>�^%*����Z0R-��a�$ �'Zn��ʏ�0c��~����uq����tܤӄ$�n�Ġ#4�oYN��H��.Ȋm!|8`��l����փB���s��'�k�5p�D1=�f����cNn����|^��G�/W�̌��r��Bu�����]'_��DjE�wH��?bg�J�%GǬ-����D#/�]�oq�hֆ��,Hƚ���՞.i���4r *R;�����.�0\�������C��˨ҋ�8�Ӱ���ؓ��3&(�ƣH*q?٦��;K�	-+v���0�~��Ȅ2���=�M�2RlB�k_���cU�mv ���h��x8��w?��"O_��6��!�[�J��Ϻ�*���O%.R}{xZO ��P�Ns�؎6�֦j��+�(����bM`Oy���>ۈ��p�����:}��|{��o�{��s�a՗�e��@���Q8֕�؝-p��%�-��46��yd�� *%��ĝF �r���=�Φp�$� �.���nХTuw$Q�uAa)ɬ�"9B���v#>�a6�ch/�)�б�#4k�nˆ�g;7 gx0��L�P�V �Ca-��G]e���>�Vy�:�p���@kP���~�,9|d8k�v�q��9����]�n���g3xdi{B�k�v�q�<�N��/D�G��߾�ΣP��Z���d�Q��$�s�b��w����@�ԇ�M����IdD�����tjR�aS�߸��>��$Z��e܃�f���e&V�#��$6\3XB����$�|����SWD!?5&f�Tġ�����	~?r�`Z:$��`k��9���h�N�,m�������L[�����1�sJ����xG���+l*�$Ԙ8L4�D4�9�"B�jj�-ְe���H�Ь���h�uL���K���Q���׎&~Ca"-%BWδ����}�շi;V������?�h����5擓G�y2�Ө��zDO�Df���k�o>l�����fs��_��a�v������� ��vRf�u:�oº��������nEJn����;�0��&c}i�{��놞�\�}�'1��������F���DFᱥ��}�"r"!L�N�o�S8����b�Vj,�z��A�+*�
�/�ɳ9��.:��$��Ȣz���G**  ����K;���Byr�ۋ�� �Z�ϕ]c�6�y������N��� $t�wV�=f�Iė�h}[*���\t�2�禙+7�A]Y�5l��M�onZE�#� �G�9'cC�
�j�3��!%`<��`C�dJ�4x�gv��/C���u��)"��/A#%wOZwy٧(�i4�bY��-?!�٪���ic/(���$�vP�N��h���If��i75%@���	0%ċ�z���1,@]�t���E:pk��%:��^w�z|�d\s�X����]8�7���z:� ��2&e�V7q���q��o�;㚱�1�<�@�b�TTۏd��&<���G��4�
����(%�`[�6c]s�}H��ج�̮ϕ9�d_�s _/�)��Z`�ۇg���(�����$/	 �w�5R��4E���J�D����{����3�<�����(��(�/.�2�cU��,U+Ԉ��p�l�%�"̍*�H<�;��o��mhFKF/qƵ[��4;�0���˨��ɞ�Uz��`>ߴ#h �����'݂����0���ml?V�"cd&��d���w9ixeD@ w*sAn���6�Hr��Kf�kJ%ώcHHHp~�8��/"qԗ��I4�To*���=�y�X#�����O���)���ď&���S�f�Pg��LV�3�(��?h%Rm̍��>��f>j���t��:�w������S͂@��:����'���0�e��PM�B�b�D�݈�2�i�����t��M�NW|�l�c)kQ|hBΰj=�s�`��<w�X�C|}�h��̂4�5J߇7J+:,�q�vPp\�o3h��ό���D�rN�jUp��3HT���"X�S�j�����:�;N]��V2D�b��@��>�)�8Zo����D�M�8θ�҉r��2rz��<�ޤQo�⒕�]����kc2��&e�F�0�،g3�A�5nޣC�$8;���ѻ��-u �c��hE7HعW��������n�c��h�����dϣ�̍����nc!�8��S1�O�.���P��ZP�� �X �$1���8�a���Uq;lO]׺�r�[#����DS�Rt��,�7�Q&p���mbU�8{>���İ�r�L�%�A8�S�����{��@�5�e�x z9���B�j��>{s\y� ���
ehYӨ��O+�̳UM�����m@�Ҋғ�ŕx�j�}<j��myHz�o6}�_�YI����O�F���W���'{� ө�M�o:�8��J�LY�[�B�y/8�XU�����%��g!�q�o��3��U��?5��z	܏��R+&���_����~�ű.��o'A����%�����PD۽A�(��`�|��Q"*���+��;�&cq/;�4��P��I�A
�bm3�T"(�'��s���'^X�~�M5n������x��8s��]4_$0���0��r6��?F���D2f��LyXG���凌��	�0��$&8L�2�VM�UF� ȉ��Q�)�.����Wdզ��҅T����"���R��l�Ȩ���b�pw��נ�6��I-��94̴j:��x��'��`�Q��PQM��xCɆ�
��d��-��+��J��4P�>����=s:J���o��ݦ�$K���c�2w~� K�=8`�~޳;6vW��))��U�<�vxdmd!��ϟ��z!�BA�H��&� %�y�� �%�
O]i�'2���>aq��@�h@~[�7��=P���h��83��֏��KF��՗	�a�`�S�xqi�F׹���V5D��)���NI/���vQj��/2X��7��Qz����y��#���X�p��T%���>�
P�i׺m��C�ޖ�t~��m Td�ƴyP����X���,l�����)�T�+m',k#A���::VR|m1ʁ/�77ȶBW^�Ԫ'iO&d�G�H�aA�}�S&�}p�2,�g���԰{���z�Ȩ"��tZQQ�*��[��E(��8�dC�Hܕ���,�[���n�<�eNR�hR�4���ݲ̑�7aОͶ&�4a�󬑺 ��1Q����k}�k�-�����6��ZUI�U~�?�_�7���vGjj�t�'쬹�IɎ!`�'_�VҊ�CH�w0o��M�s��J���i�g������$Exq��k�ϧK�����ά9�Q�0IKN�������K�3%�;p���b�(�E%Y�](��`�)W�O�K�O0Q�s����>@r�0	�ҚC7�3$�Z���e�*�����
�Xj��_Un6�J1�!�^6�Q��%3��Ib��<>bg��W�PmD����@��<��VN�7Z����M�	�"a#��q��q��Y�rm�Q7��$�IB��$� �ի�9SV�J���$�%W�&�¥i靉%��`�A�&$9EfI�@Q���葬�*�;�mJ
�9�_���K�W����`Z3�&��sw���]7�Vj��*]����"�1�	0��������T4�c�����j��x�[¸�\�������̽ H:��VV���$�_>$<
߅�_I�k|���N�T>73e��fw#s��	=a���mg��ӗN�u��.�2��Y��*���Z��KT��]�E�;d}ҿJӜ�L��#�ђ�Tn���|'��r4�`)�ST)O�ϳ��=���aq�;��
R��9�B��$^��W����H-h[�rZ
�s�O>����t�Ǵ�4O_T�^UF\��25�0K��#V�fB� ��'bl��g���]ͷg���_Q������'��Wi�B��fӧ/$*�v?Qz��~��g��z�W�%��J�3����W�꺅��l���W�D XbZ���q�_�y�D�}_��Fr�W��<V'�h0��$�`��5��2�k�UQO����Z걜)�[A��InmiB�A���gmP�-v}��E�>�=ߜh��Ј2�&�DJ��2�Z���o���a}��4a��8�B �x2f���
'��Ka�+���Ԗ|cGɇ���pZ�g8#��U��-����,�۝|����x<��}�c���rY��x^��>Դ��gW�໋��\n�����{�qXdhc]�+�.�3��g{G[0ؓ�.&�})6��[ԫD�ڿ6 ${�G��&$E&9�y���:���۩�?��t]�gz�� u�H���Ģ~F�\L��t���c��ү��z�����c"V�3��v������K%ݹ��y����՛�	nI��Z�̯+�n�~�F��vY�b�_~]kvM��v�?lw��y%Xy�h�$�+�/���}�du��	��˱O��7�	���>E^i �<`��4�o�O�Ǟa�\�/E2�]_�q��.�`�#4�&�~��u۞o��~;��42����ӕ��lNl�6��*�nC��y���|�>]����O�]���G�
C7��\�з���T.C|G|���W���W3�/ë˿�H�_��YtϿ���5�Z�z[-�y�Q�F��c��p\�}����2�(l��[f�O?�*��kzu��(�ԇ%biJf��i����?�欎�sLg�b��r�Hk�4F�*&=�~S���U�fڒ����W��7}*5wK?�$��6�"�x�>7I_���}Â>i��j�H���zm��6����t�����O��9|)�m?�B�u��fٌ�^�Hq=����P��`��Tg/��6�
��Q�:����q�z�O�Kq��%_����:w���m�
�L�L&��<��'f��Zr�#����߸�}�R�Mʃ<�)�Y[љy�f=���E�"�b|������l��Jz.�t�k�m�����F�X�YgR�i�f�_�(;�����/+��j�O��H�:Z�`�i�>����l3'���O�p�r��x1���듺Vľӭ���W.�l��N���<�T_�ebſ�%�Kݪ�ӟ�:?[�����y���q���o4��#��;:�]%�v͙������s�WKN^������{�3i�_�i�G��ŏ��B�+.���C�\ѽ��{��������"U��Q��?����*�0y�jox���mi�s�zi���[(m�q7Ι?�ྜ�/]�����n,'��c&]+���*��w�2�&.�����.p���܀����I����_����@7���܍d�����
� k$ʴ����/ٿ��<�~�ߊ��;�b��q�(�7{����i��*�RP����DJ|�@6�ܮŶ��bui))���S��;��^��p�x�&M�Ih�p�n��.��]�c�����������->��=<�����{�֢0Ԯ����wx�+�_r�9�5�x�>��ޖ�
x�N��HoO�it��4��s����;,�ly�W	�	wa I����r$H�(��.@�р�a %��(��h G�$��9M�����y�}�N��ު:���:@T�*usO�~�ѵ�,�?��*;�*[x �o�� T6�0Pí� ��������;U��ZÜ�[�,��:��׉.��G�C���Do��Q�G�����R��q�tt� x�;�Pb���\F�B�L��s�;� ��]o^����|�d�c�L���g��'L���� 	 ��:o�^�3넞�����yUN	�Yy�� hE���ĺ|}�ɺ�;3H�roqۅ��bA�)c�yt�.-N;�P�U��[G��kfg��r�ׯ~N'ܡ�����
(�q`��K�2�':��=���p'@��+Z�)f9��Cu$�aQ������?9;=lIa��� ����{RӜ�3)���!����ˬ��"��9)֑�}��I�2Ȇf̭Q)��S�e���[�2+g�W�r�����n|/���v������_��x;�[A�����2dnb�<�a*�<G*`���Э|�F��L
���Tj$�)1����S_�����c7қ���aD�f���]�U�면țh�	���r،�
�����@9b�=2~�4D��j�Qvc!^��N��7�-fh�@5��l��.�b�ܺwRA6�獼-����|Cq��V�e���֒����$1� ��h��w�H��)�%�@�^B(4����k����;�7��"��DK�7��Á���*;~�#.�7����������s[�:Ve�Pn��F~�cH�����
>2�H�n 
��|����ϭ�pS�+���:�Jd��;3}�.M�� }�!q� N�6���w�*�;-_x��{Z���1����gЧۍ�i(�cZ��mc�;M���3�o��ꙋWu%a�g'8?֬y�\{~��lJ�Qi��	�(�/�=N�q��J�/�\�����Y�$�{���<O�Y�*�����.A;��Ytz���9�Kq������o'�����A���sO�$�[O�b���m`���?hTO���P/�S��[����[�ͪJA�*?�rP��T�'5���NtD����w����?�L��e�b+�<��V��дqr	&��r#�C0��3��i�6k����6�ͭ���Ke��.\H�jy;Y	��&p�G�}r�JjB��{����I	�������(V2��A��k�n�s�9��V>��M��ʴ���Iھ�Fa�;��	��6�i�Ň�1����5p�����z��ey�\@��M��q-J�y(�F��c���^a7Z���g��\�ŷl�w>z^�vr(�I0d6=->g�P���n�At.dSұ�GW��=�A̒���U�t��v2ׂb�o�0���?M
�mT��r���~�R�>�!��I+������j�ZY.Vw�Z�h`.��JS۹	�����+�s��]��t+痂Ÿ����\���#%39s0W���}����� G� eٌɱS��
6 D�ӽ?��C�F�tlb�.%B�E���jP��a-��
`����v��v��wʤ\r��/+���R؋��.΍5��c���c�|5�5;�6��K�� �{���!`b8�A��	ŗqc�W�!��3���O+��$Y��o�,~j�a��d�	�'��悩�t�nČ�~�Hu\c�;8��79� ��xU͸�&�g�Ip�I�Ӕ�Hv���m���4�Od�����Y&%�D4�U�*�h��h��z��<��c�hDX ��4.z��(��&�9���$���N_?�� �<kg�_�v�u4��h��r����\��u(d�2{�����;�ݭ� %�ƋAs��;��*�L2�~�5�r2���B��S;�}��0��<�yğ5�z�i��%�)Y.�s�Lh�PxN��8.��_�`�A
i�ދ�����X���o߄Mas��������L�[ɠE�wD�"��5��;x%��v�k`.�d��<�F��"q���2�V�S)��}`F��� �}��:�T����e�-��s>�Y|�̷��`=�Y�7.�6�} Ngf���0M��t�w�t0X��&�ϾZ)�"Ϛ/R�R�z:ő&���-1�Á��r�F��[-�o%���+��ߠ�`s4[������7Szۼ6��љU��Q���+�C�D"�N�Z�h������f(18m���:[��?�<�j.� ec����|P�(a�(���J
(��	��tC�3�[���6S��m3+�ZB��	�A�/Ո���*�#U�-:2l�-���g�qb��C�
tR��E�҄僁�ABU|Z│��i�b�D�����m�+ Y���.}RJ�x>����z�����Rb�4DI�F���?��l��:���`��y�6������8�����7��.�iWwق����ގ޸�K|����ދP��f� ��	Ɉg�K	��F�N�����FU�dYQ�q ��0��?�ѐ�q���<��r�CY3�K#v��S�6(�k2��&���:��F����o��s:ڡ�[a����m�;��rPUJ�mZ2�����m*��.�g>�y���9���dV�թ�����F���kxd.𐝯��G��o�V�7���H����z��="m�W���O��Ok�t��1`��Xs�6T{� �[�X�}]��t��F�s-"��DZ[��8i�>��q�nn|�;(�i!�5�r�n|�ج�TX^�6\��]<��(~U��%��c���LR�Y��MU���ٗ��5zv"z��?ƪڃ�� �~����һ\7�i%��'Ui'���m�iH�:�g)�����Y���7�# ������=�U��ϋ͝$\�^���ެx�گ���"�ZQ��bk�>�r�����@��6���!��3�iÊs�X(RRU��^|�"�=���!we�9�v������t.�xk��bk�Q�z�*?���"�Z��¢*|lE|ޓ_���ά��|���_��QJ�yJ�:׭MM��,�в���"��t�� �n��(i���֋j�b�CA��,I���Vy�A��|i�ib-	��KF>;)w.��ֶ�&��H�4?sۛ�$�Ȩ�����~�wP��?�N)���S�Tbŀ*���e�=g�&LISp�CQ 'ը���j�6��~���/[�������X�=���.q̅�$�>�����ԥ��
vw]����0_�+M:�$���x�t�g)-��c���Z\�1m�[ރ\9�
�h����7����Ag��r��mΨ+}�Y�s��J���Ѥ�	��8L�f�5�a�Y@����ǅ;���hc>Ș22-Ͱ�Z�9�b�u+f<��8 �|#��
[��-�{�h�z�ɒ{��o
�Q����`�V����?y�ކC�v�9?��&� ���p��
�i�7	m\�Ǒ<8���#t���<y�`u�I������8�(����Ҵe?���Y�譣,�)q�C�Zc��"��W����Z�A�A�E���a�K:S��CBd���	�Yo��w4�F��8	���|A���#o�wc�ޡ"��� 4���}JQ�������W|�Z�I���`�^/������za��k(��<][U?H�:�5`��K��������C@b�AZ�˰Lǭ�#�?�:+>pNj�?.��������S����-��f�99��aNK������Jb]��@J���y���\ ��[�a�ʣJGA^�Np3�G
oZ�#��/�3�,��XcF}�Tӕ�z
t�u�_O��Om������p�W;�O���Cd;SR8�[�~Y6BW
AZ-����5���iJ�M����h�����[|&.[��}���Ե+)E���{uh���4��MVJq�W,W�l�x=w���/���F�j�E���+�HH�QT�9`un\��{9Zcjm�]W ��ӗ0sQ5�-97�,
 F�k�l\��=U�"&P�'@�_��8郌���2�䐌x�|�6c6���ˁ�����{�KS	qQ�����t��('�T^P0�°S.T��&"h�55>ϡ˴�Ѳ��j��j+�|��P'WQ��.��O97��V��B �W ��_��/rU�G��2���3�,ɝY������
��)�bNtf�m���\�b��;Ԭ�IU q 4�di��񦣮�����Pv����EF�Y���ncb���څ�=]��0��]������FTN&���>�+�c��7r�TӾc�R�I÷�⛔o��͡�w��0��56��Mb[��i�o��,�$�3kȟY�^��[D뙔��=��ː֩�<�)6*���q��7�f7㮕��X�NxZ�}��������I��[S��+<3�z���La�x��&�wy촻�V�K|�!)����A�A�FQп�}�u	���V�y&��� AbS�y`���$���z� �P{����ܛ�O�C`�G�IW^Ć����C�E����V
�Ӻa��$�&���Ȳ�~%� z@,������(��G�z�I�S[Y&��.w�7�$���~�jY�=���t��h �EP|�g�6�5
C�#�B�g۾?12}����K �*b��9�����]:�ty��"��{�W�l�\b.�l��Z/�Y5��Ż"jf.w�����C'���靕h���)��蝄�Ût�+�z�D;�(��˛�j�X���Ȝ���c���
��|Q�t.�/���]����9
��I��lX$p#��l��:�f���*ķ�0���\�ֶ1����xT���c�t��(����Ǒ�_6����JUwz"U�g�ޞ"�r<B:*���b�Ý~�7V�)]U����ƏF��#X�b&&-`Z�Š�����克�p�2[���j�����`�LrMԲ��+/O6'���t�.9�A�] ����2Uv>���n;���XI�h[E�_7<��	���$̣T~	PF��"�Pv�� @�C#���-��l�A>�`m4b|��I��T�ZBKH���E��<s�pʷ�+�uLfg
�hz}�G�5C1�Cn��9?���N�m���$�n���ST<�̍j�!ΗsR�����H�t� ��Xnsb�{��BPyԾ��le�;�0H���p�g�T���>te �.TauδxFR��gq��X��b|N���**e捊����E�b��4F]:Ɨ7�tk�Q����r>��Ƕ�'B� %:��_M�Y,=���+�yWE�j�m5��<B(��K{��	u�2���Cb�<�QJ`�M  l��e����x��.��m���K)��˭a�F���}ݵ?�}g߽������'��ӊ�K�f����/�"�A��V�����ZϬ|��y3�T9�;Q[WY�v��V[P��Q�9}�?��tc-���I�jhlUFWڱ�|��GWP �turZ�b�+@e�����#�tn%��Q0�H$�#W�n��O�MhBH@��a�]"�ߒ���L2��㝏2�އ�VqS��1�EaŘ�SA�][�Fy�|$����B�h�Y�a��� �qk�q�ڣV�w���g�@�s�ܪ��3�N�~��4�	�k`e&�j���y�%P��
�r�e��u	����%�ǩM'T���ŌV���xz�ʅ5�L�*��ހ�tCVG�t3O��N��ZOb1Te�k5&�3����G���of��`<i �-.�9�mk�B�r ����
�U$��?8��ip�"���N��R�*V�ھ5�k���wS6>�-�k����3Qk\s4Y�/�a[W��1z��M�
w�.�{[��>�<�L���9��Z�G>{�������̇�&��Ε��߅� $��Kj6z��x�LT�,vd�nG��T�弾�-���O�k��.�n}PA�-Y��{;�V
�[xԡЎj�ۿ�(�݊ �]^���Ox�Z�44#�ё��Trb%̟�ڣ���?�k��k�+���T�;���F/	-���o�kY)w�z[^Q��HS|o����|E=j � �2(Ot�la�X�*�Q�K�!*�+���ՊX	pʢ
_ N^�9$=1O�`��l����tZ�U(Z���a��)�<}��z�ud�34FK�f�Ǜ�:��͍�`��x:B1w��Mq�K�mm����V ���<�2�?%����\�����<Z���#��'%�A��5P�o������/�BW���p���9����c)��A���咼D��皩Ϗ:ax�F����2_����3��I4�yi�rP��OpblW��/�p�|�(E��1�`�S�Nv'�g�EZ)��j2޼
�%@��sR�*��6�j��)t�A�h���;��f� Qy�N��z�i<'ds$���8������p4�hi܉ M��[RC���(�!�G��<��zƢ+m.�×�MN3�������z��Z�:��)/�GL8׺��\��{��m_j��c
�]3�S�}M@#��M�oޙn����~5AO�Qs����[j54eՕ#��+M�x���Dᕝz�|(�����Ö籧��
����}�����
j_.�_����WS�b��6ɵ���g��Q�E��΂MT	�]z`�@�>���F��#L&��BBg�V�P�׀TF-ע�/ݶ^xE���&j���~�����z"Tw������ m�x,��<���agN}k'�s~I�kc����2tŭ$���<,@�^4X��gsm��ڴ���6ir2Ci(�cy�]Y=���4,59M�s!M&�u�j��į�"e�˒��E�s�y3z��[g����JW�f�<�$Ԋ�P�O"����i �g�����d7�=G@�3�S��8-*��nQ㓔��j���H.���E�'cs�a�1��z�	%��:N�@7|����S���qP)2"N	۰��'���T+���D��P�W������j�!���V�#m��P��.i���Y����)����]�e����2'/�2QX���uTr�^�B_���l���|CGZ�o���(���9�t��4ڌ��KkA�0�\:��J�5�[����(�2�R��g�����k��we)OH̉Z�eT5n�V����\���܀����&�5�`y ����k�� ���/uG�l_�$޿ڙt؄}#tk��3�JFX�/�������Hxx83���&��,��9�"@c��đ�#�QCPT@��ϋO
���[@S�����g��r�
�:M���_Vv�* �q-U�hk��U���}U�����:�*����'��JrkG�),����p���OPHXC�� ��?��?�&>d<+}Ғ��,�r�}N����������$hz(��d�8�a��p9����3;4j{�l�N؄N�� "��[���n�6`�nV�����uq�k�����I�j�ZOc^Г+z�y�=w�خ�63/>�DN~@*���0��
�b>�:��i����/#o�yJ�ƻ���X�R
s�)�}a��Wl�?o��ZF��7=��E����T���
��!���ܾ̩���;~��<Q Ϭ�������B���cdq3f#_��yt�q-�A�3�[�� &�@,���Е��釾���<+�4�0F��ǤrZ׉'j{�|�6˖Nz3��;Y�ؤ�6���~�x�*<+1�>kW}�x���� ��;��* �QZ��!�
�ퟎAVg�}?�_�3}��}�o�k,k�����:���<�6�|y���^�D�G���i!zWv:����}Igޥ��޻��߻Ln�;V%�AW6M�=P�T��e1o�r�t�H�0���F˩��8�ƞ���}e���l�es`�����N4~"��~D3�p����i�r����Wֻe I;ɛ#�?�3h���`��B�<��xG靾�Y��i��S���t������������Ç��#��on\۸=ul�
���V�^yn�Υ��N�E�<�jN(}�����Z��|#�Iۉ��G�d�`P�|ƣKf��&&��m,E9 ���q�s�i�OB���})�f����ܓ�Y��¦~� �L���=kZdk��I̾E"p)�G&Eg�/u�Dr�r��o�2~�$���k�SY�,�X?��s<�����T�:�S9����~hzϖ��/t�2T�0��H0)�r<`���BT7���΄-J~h/���|Z��)X:��)� F~s��Q?� �j�E��pg�>\V������f�$�-"�AWj��ܒg{�5:!�굺CS����@�k�B{}���ͧ��uh]Do����;��	���[�k��꺱����,3O�U�y���Qh��p�"��bOvl@4��U�����^+MܾS���`8��L�NeI��D�&~!�ɺ"�_05��GcC���/�L��&J�~�����-?�S�o>���8|��] ������k+N��w0�׷�g��j�f�90(�:�0��T�Iқ�}:�lP���B4�_�wh�g�����Xv��� �Sw�8P���ߴ���}�����H�L�\)�O�Õ%���?��-�,���LH����ɥ��?h>��KxWc=���-����|�h�����c�z��X��W'�C��G\�!)kwFg4ɻ-є�,��-KQ�o��$�ۺd����{�`�όv����ȃ(1h��ӿ�"(&�7$����YH��=	�&�Z�k{Km=�ki�A�I�nY�y'gﲵ��P�.Y:�r�(C73�2V�(��Y��6Ֆ���M�) @BC�l�fySO����R��L�
w\�P�x���j>�ܫ�� �Su��*�/��ˡ�|�ȧx:��_�v��������g �}?��$*̽���df�&�p�fk���1.���ߡ��g���e.��-�'�F�e��xa�U G�&��{��e�Y��#O�F�����+?��l�x�ч�P|�O[~iWmj�d1�X
����:d��Y�W��#0�����u��}��������j�xZZ���a��LL���x�����/o�5� �N��sa#��濥} ���b;iM��2Y|�j�h9��ՠ�;�v7����9���F�ŋ�FP�ňM�"�X`��J�v��eh���E���2N��oޞ���|���l5�s�e̾�9�N�>~l����{�Sq��ktT�ڲ]�O�_�-uXw@Eҝ�n{'�
�;A�����sE�V
�ei0i��*��1䶢�cxM����E�x�* q���l"��Sϒ6�!�v~�d�\kҗ��F�Y@;L�.�����\"k獊�����o͕@�����]aVi��Ȱ%}P�:��v��#s�ҵ���%�{So;D�I:���W�b�M�
�@��� o� (��STF�s�#U/㺸g�6��n�B�}>a�����tF�Ү���"law6��Z���q �t�m���D0C�^�� �	��Լc= VF�D'c���?:b�ݓ�FU���8}H �;A'�	c��1|t 5VȔ�d��:�j� MTj�u*�qu��V�z�5sU%Ū�>�f�`����-g��\1T�F��K����{Yk˦E3y���@��V�V^XE�̓xw��ؠo����qH�"�����1�X#��Bȕ���?'��,%'&�,�e�S �MN��S�5�B2��Y$[��ϱ����������fpʿ��v�~��� ����h2UV���z��UQ�u#Y�k5��4yи �U�վ�8�R|U1� R�իrn�3v��qq��#���Q)+<�P�O�Ԡl@��׊��$X����}�
�*�X�J�+��;7�!�W��r����|��?wd�:��XB���X=� �Y��׵��EUW�NQ���\TX{`���ʺ��3*���v��j-_�Y�^���՘�|���e�<=�$�x��F�O7�͎'��:}�kE� �Ӭ�J�_�+�G����>���@�V;��� ��	e�k���PD��}�{�`K�%Co���N�=�YZ���E/��PJ���3�S���D�DF*|� �ל�u�����At������pb�u�T�s Fݲ�T���躴t�z��R�P���o:�����`�i�Ykؓ�S���x�L�����Z�2�f7J+��i�#S䷎�&��ǃ{ZP�L� ��$=��S���J�wc��{,�N�D]I����n�p��Ϋ���m<Vf��/^4��C<$�NR����i2b��J�� ��[J*��l�@���@�S����f)�ߒ�H.T��j: �f۾:�g���U�|e����:��瞾���e�%���ST��ݞ>�ڝ��?���y�ם��;a��������_�P3]?4T �8����OvC��R%�yr����U���x*�<�������!�,����m�,ѓ����d�[��.k5��J�/$�]��Ld|Ʋ���F! #	�����.�rφ��"�ӕsd㻟�j�k�N��tg�j�=M{�kS�޻���"�R��.�;'F�Ā�t�1VUKƥe��k�� `��W���0i��b$�nYZ��_���{ s�=�Ǿ�E�d�/�4��V=� �35��Rx����e�EȈ��(ŗަJS?f����~������_� .̛\�j���#d�t=�t@"���dO|TC�T]�b�"Kg�5��ŏ{4c�p���mb�;0Y�n҇v��JS+5�Ӽ�>k	���@���V)�� Y�c�'�Fl�I�S��07��1;�!#���~�'����FxB2�~��|~�����/�#	o��н@ad;�7K���?$��3�������;ܾ۠ ����a̾�F��P6�}�v�&
�7�mZ^ϻ�I��H�'!�3��S�O����gR`���E�9�?�A�"4�O��Gn������2LGC�5�n� ����fw���2�Q��"r.����Y�x��rVCr��(v1��&��H3°'�~�-�g;r��8�_ȕ���ڸ�Y�G�����bc�ul6S��l�:�h���~b���Ъ� )_v,��s4�S�� ���(G[IP%�|R�H��W���C+��f �Z��݋}t��!P���ꇹ�����x��@�˚�d{��z>�Ĵ����T�9�VL�Xp��+3�~����L�F����0�~l�G���� $��:��5��[�ڙ��%��>�1�ꜯ\x�hp�8u�F���R�1��͘�Ud�r
����𤃊R��s��ks0��%�6���p�L����d��CNU$��ڙiT�P������)�k�ݫ�ɖg'��8
	9��Sm�3�Ͻ&�+h�rL~�T�W�M���/�c�A12�%�!�U�s~��Nߢ�u,��"�>�Ƅ�h��ߖ۔�I`�؀��[�q�����Dm�r,��g�� @��W]*+�s;�����/�9ܲ��qI��k?{���A('I��u�_~[>�n��jP�}d��KP�62����8I�'Ȓņ�lɛ���y�AH�;ߜ1������F9��N�\������P���^7�}��-�p����4�jD�zM�A��A���|��c��d��U�C2c�4�CU3�y˵���.I��Ԇ	aJys��~�ct�F�R%�]&����)���Zo�5Kn�������L��z���3���מ�'�M\_&�.z\��)��%siÕNUc�d#�yS�Ut/E �ۗ�k�d�%��@4��X�i=��$�x��8E�*�$�ק���T�춄r*H&�v���l�&�?���Y���?��ťC��7�:Y�W�b��S�=��7�AO
�z�ZMƋj�����wܝE��1ݤӏ���\�ƾ�'GEJ���^��?�2���c`{P��ŧk�mh\�*�����1���ϛϜp-��_/���a�e�{7�5dc:dF
��&JiL�>�+<F`�|�F�;^�5Ӱ�a�!m����0�%h]�B9�Y|��w�TY2�27����"���Vf;���,��ǡ�f0��luhۍ�kXǀ�j&_��CC������g���E���$�8��KM��;6E��Ӏg�C��p1Z!�l��]���4�~.@����~�4�	�%�3}�h��aas���Ճq�u�x�U�6�N5q)��������,'N�rAG�=3�}K�ouQ���ں�0������n�v��+��h(8�+3�i�cjv�_��mȭ���LhL�6}��Nl��me��A�H������
Ŧ�]��­2ܪ��3Aˆ^�%����n<��F
�6w��F9�;Ц�����!�z����x�t�:�=G&>�,N������o�L��w�%��OAx��S�+�/��a���x	^7��t(W�k�_N`[<{���.w�ѥ��0�'�kᆬ�>Կ�'��z1�g��C= Pc��s��^���6GT�C���緖�۶&�v2�-%T6��y{A#^p���� �.��GU3�=��z��%l�Y�6[�h�f|�}׌i�B�^q�����,}�yB��G�mi�D��"����3\��><.�(-

)}mkn�]WD+��;6v�C�=�C���G�t:��& �ڝQ�`�����bgP)�_$.�n�-�;�ۗ�?��g�`g-�ץ���չ�\�{�Yit�a�Rn\ PX��9v�M��W.p`��-�2��C��a|m����2�*8P��,��N��s5�Y�Y��4��G헻 	OgI�T�#8�d��,`>mhY��; ���$�#����.��*���i��f�5������kT]k>JV�h��3���	 S��Y�{^�
��}��:tsm��ͤ8�0=f?C���n�L
0BǢ:Ty�b]:�X�0���CxZ��>{��%�vvܧ�s SŞs����)�!���y-�x�Uq���C�}O+s�':�t��w8J?��.�*.��Fu=tMM�r�yC�p�*С��"�(�B)O�{�b�߇o9�]�6z�]�� �N ������OA)��:9��e̺�"6a#@���^U��&ɛ7����=���,mk	HU	�u|�H-'��'uac?�D6(My�2�v�����<4.'8��, �Qm�u�h�� 8<u&�r1�_��������Y���U�農X͢�����=��A��z��6��<n����f 	p�� ��L��N��D	������i]48�C�]eh?�]_�uTi�X�����_�wE�j�}tm˜=���&�-�o7�`�AOE�T��k����h�	�~�}���`AO�h�꺁��S�f�֒ �����݄>tI%j���s�i[�Y�铷q	�%�U#��������.����ã��[W��l���@�
��t|B#�L���w���,���"\��]�?e�*'��޾�.����x>���p��]'6�3�#�z�
iA�;�Gχ;0�4��t@��|�]{zs1Vg)z���xق�X4G%�(��B\�#��q32g�C��Aͻy5���m#��BL��4t��?j*�%�	w`^d=F�XY�����m>�� �4ӊԸ�؆Ǐk{$����D�����Ro�NS��:RO]ݫt�����@5��h��)2��  ���jv3�������]�U#�k[�x� ��.za�E��ѣ�q�T3�A��^%�*(�;���vD�o��X�eI�ɪ� �tWQl����Zw�R�Py�%hQ�Ovs�ݠA>�K�P=�{�+{��Ɔ���۲���$ ��9���A�Ჷ�����	z�pdH�v�C����OǯD��=����Z��� >�\"\��0�X��"d2��*=�򫸂��ZM��2��^.�������TR� xI�ŗT����T���>���	��~����)�|��Ho9�4v�WW������T���(��z�\�����K��{�B �V�����.�j��B����JM	��<D9{���ă�b���Ϋ�?�s�7@��f;3&�OW�8�uJE	�Ԣ���ro�a��J��h��+�a-���o9e,\VOu�^�"�Ǿ��1��,�VW���ۃ���8�U����7��_�k�qޭq�ؘ�w�2�jzxh �v9�9��dǚ"[M�[�<0p�^��^w�������?��v�`�9R�?Z��Z��bC4��+���������S�F������K�9�cɀff^+"]��Ž5	���D3���c������¸L�u�/��E��!M�W���W	��_w�{�ǔ1$:�� ���k_x��v�4�8�v�ȅh9�n���������m]�z���Ɠ�ڋ��-ZI��L���T����L�1�1sk�W&�U������+��G+�q����1�B�N�ӵ�H�˜��Xt	�.@�]�4�2<J��Ƈ�l���U ��o�l{�?t��o�aW������?"��;Q1�Yx���� �$�FM�E�1:��
��S�� >�D��t�E{/~���.I'�C����j���'������\��]�"��!�A�V�M���[Um��5@$��u[a�1�j����e^-�,4!��1N#<���\C	���.���|]���fC�I^0���.��}���/g䪱%.U��Q�p��v���V.�:��:��J,ݣEn��6��}/5 uN�7rW�.�"��z��M�����ޅ|f�>XJ]��2�s���c�Cpo��2��6����>I���>�|�;�#zR���X�K����'$������1�B��$ŵ�&��3t��(�K�8S���q�������ޅ�ܕ��c�T��8B?̾Y��y�{���f|�,z}��8��M�"��Eq�>ݞ��z�~�gh�v���ͼ-tF�ZD�t�n
�g�$��U���c���Gy�l�zӢ�`��t�w7:�r{k ��8��W��>�s2����9h����%���M�ъ��F_��m$L��-�e˳�����z)��H��Q\A\��,�g?ǜ�7�i��s�(�etܒ�5�����)���l��F�DC5�{}��������1,�J��2���RG)j݌+x�F�0C�8;�)��+xn��p��(�Y��*��3x��,�]��A�'흝����O���(s��¿OV�W|�x�&��A.��ˡ��v?�1	7��s���'Q	wc=��LN��_���B�}�r�g�2Sz"a��͠��<�3Q�4[E�d3�hk��osO��Ϋ�A��ߓyQ1sx��~)z�������w�Y��ȧ���H���?tt�/@�(�@�oekH��N�`�4�4��
�Y
��;(g�O�Sy���j�����ST�!h���\	��H��gv�C���/��ǧL��#\A<	 ��Q9��%�d1�7 �%�wJyz��`�E|�o�� h����,��C�?1{Pb��
i�d��po�~���p; �s~��z�]\W� �]��owe�bmf��j��H��u�tu��X�ZҶ�Ƥ�Y0�Nj �]/T��}���`(G���C�_L�Ŀ�A���}B�T�]�Ʌ+Pl��lx��$��L�`�.fS1�^.��Ό�?�̍ρG\�^L��K==o4+(��W�`�]e�?��� � �'���\n=Xu��WO�M����(��`B��ms�!a�����a���GU�d]H�?�xk������7޹�o�6Mt���h��W��Z�e�/�7���v��&�n�&�£;4�sR�� �� �Z�Z4�:3�{��I������i�p"���c�# Z��W���9��P��D	�Z5�>)�1j�R�o��_�mi�>V�T�IJO�����o;���_�8��9�*�;�J���?��#�I�Yx�|ޠ��aqU�e�Qv���Zq �����0�Uz<�a2�j7��R��*~V�.��@�se�|J�5*����}*|��x�����'�R����ePs��̌���ypPo2����uj47+�#� �Ճ.'oG����~E���K����x{���(�L�9y��3 �ܾ��e���g��+>��l��m�[��U�����/bf��R���P�yI��1v�򵰏V�/1�v�slDB8�C��:�j�]*Ǜ�q�pK'z�҇�r�k��䵇�}ȟc)W��;��i缍[�l1�NG0��K��LF�[��pxi8���eEK;[���� �Jq{}�j�Ja����Ըt/&/�);��[	��-7��烓��@�G�G��j��`@�J�z'$M*d��YBW���߉���*���a�'�D��_�k���D'�h����ݨ;�����b�2�РNWp��,5�o�1՛}B({Ӿ��l����D��e�ш<|
�V�8@=yfk��$�'�S��
'�Y��WJ��s��P���jo���*��i��@r:�Ќ��O�<��t��� w��8vQ�X�4�� @�N���1�ZG�T���#��j���p-#O�[�q�I�3$�*�D�KuS��;qU�%��6�	 Vh�������U�.�R�`Kv��ҵ�#��^>#]:W�F�E�������b���0���x�Zw�oǋ�Wh�ӻhx����o F�s��H�����,��"�=ZwKR��C�\v%��� Y"8��-����M�E�ȾN6��E�T�2�I--�Dm�"s�*soЩYe������#�, �����Y������諫�ρ�-�Z�|�2�26*[X��5Y���@R�5�v֝��0���vj�h��eZAL��T�5�NRsZ����U�����1���%@��ꐹIe^Vr�+}W@�G�nV	.�NbwV]Ѭ�'e�=��  �$:���5~��7�LŬ��1"f ��y���h][;��w`G�>�� ��v�x�Y�d@�8r�H!��7��`}'��5s�g�;�q?��l�)��h���׊����7��W��ʷ�J��
�n%�1/�o��1q��[�����]W��v��M�{��O�ς`t�P�3����?�����tGP���'��rxz��o㥝���bx����x��|Q��M3y�� ��>��� o�?i?����C������ �^f�m��N�*�H6�_�0����,��2�H�-M��J�~A�\�M#�6z�!����,��?�ॹ�0�m0(@�Ö���{҆�E��2�k� a ׯE�0�����oA7����1��P)�&�&/vڰR���@�4L.���pW��+o��Q�	�=��Qu2�C�8������ȩ����l	�߇�u���O��+^�#.~b���	�80�����k����Q�w!���ʵ��PC�{(<r�e�5i����w��澋��f����#B�WA�����/��4�ek�&E�rzJv}�8n2��>��m���ڣ�.e�%^����BQ:�Ig5j�Hm�Y.קdz��ރ���%F��l�E|���3x/:?���?�A��L<�k1�)�_����C�!%�Ex;�L]��>{�z��V��k<L�~L��2$6JdӲ�	F�^�\|BrJ�p��M��[]`˴G�bA���U�"�M�Buq�N)�SO!� ���!�)�x�a5�x�̎_C�#�q���?�� �P{�YV�6o����!�s�t��RH��0\i8�;��u+ȕ�=(K�zyGM���9Rf�$=��I@�rm�ZԺTLJu�!~LWɶ�ӄ:F���!ɋ��C<����)P�������MȌ�	�U���A�@�N�����NlaBl�9�*7�k�Ϛ����.�k�^��׀��>D�x�I2_d7��lr�#�(M��m-���թ���ܓ}�z8�Q�@7bl4�5Fu�kQU�];ݟ=��0�H��b{��N"g���!{|���'*{Q�T�A<��J!Df Ou1�p�����;.��`m4߯�sy����{�B�PZ�Kl��d�]R�g�F\�T��y��I������@	�ѯ�����%���
g��;�g�:-G*�͸�t��&���� ����~l[~"���XN�pDHW6�M��x��?S(R�*��
��|��<��G��I���(��^��1��R���X�x@��W0�l~����+���w ��d?vɕ�j�R_8R���"���ú�������D,�0�$��	�,a�0D��T�nH�֖Ѹ�LQ��"�we�����)�Q	�lql�����BIr*zك��5�`3�( ���-"�z�/�1���L�7^d��O��&��B��j���p���FV��Ld� qP�k+��@Ԉ�Hę�������.�`�`&'�|�] HL/��h�cL
�ꈊ�+�AX��A=�'Z�`
N�9�����$��Iz0Vg(+V5�;ޏ]_�#��k���X�H X��8�ߑ�����Ü5n��i榞�ѐ��Iju��_��=X�EĀ�O��S+S�;��IȹX�H0�����~�J����.+��t�Px-���-�����n�z�ɔ��TJ�sl(�\�8�?/�\��ᶝ A!�Ny�� �q�Q�K�G�Y�XNOW_�kA9Y�^��^�g"��3��ް�uw�-K��w;���*m���C�ͩ���[oԄ�A�����|�Aj9)=yN&O�^��+��it:�8y��4�lM�|��uB��>���'/b�%@2���ς�~�����K��G�����/��v�R���~�e����3�^#.\Q�"=r�c>Y�2(������L�)�RZP��ӁY 5��]�QS�:�Ƞ�9��H��;�����K����P��iXF���ݍK��	�QY?���2���h�i��&.6�K<6?ę�R]9v� �!#X`e�鄘Y�-��"m����.�_��E��L]y T��Wn����M����J!B�� �}Ϛ}���e�ʒ*�ؗc0�dg$�m�[���{�,���ߙ�<���<�{�{R�Y�W�'�e`��_3ƨ2T�#��{Y�A�8G�8�(ѥW�}S>�<	?oJ���K��g������kod���}��'/g���O�.�"@������9V[�5`��M���2 �̄�e�\��Xߑn��r�O�n�o��R}�}4��n�g&+*j�3�\m\� .Ȋ�;x�P�'�M�������F=��*P���Y�)�L((�	�� ;!�l�b�+�W 4v9����1���;M��f:=74�XNw*�{X��?uC�U��$�GrobH]C1�Gw~Gf=��h�!�G�(>�n�>}�J#&4�2�o��v��,]�8d�S�?L�r\��gCլ�_�����S��:��h׋��	��e����v��S@V��C�}�������o-�U�W%�'T����v�юO�UĬ��_��E)��ۻG,^���g�w��6�y�	PL���6le_��R������"�w�)s�'i��kb��a��﬉��`���f�c��0������
�
qHD��Gt�M��.�k����3w�{�3�:��K1��.�2�ك�:B��z`�m�rS�(@:�0+����W�lI����n� ��>��u�S����5�t�k˟g��eÚo�]�,��ה7,�o�����zA:�(.<h�3��墣�E�_�>�������g��]�ډ[ty��_#S����my.�& i=` kh�\ս���BnۦO ]8	�IF<qg��还<-��VS8]c	����?�^����	0�� q2 $ׄ����Nx�ó~�Sp�O�9q�����h�_<gW�|�Bp{��%tbn�N�ȡ[�]�@Г����&'�u��D����������f�Dz;���O��<d6���~��1��T`��ob%���h�S�f�*��Y��̀@l��qn}	�?����?�t��'���1�n a�7����+o�N<�M��1苒!`���V-��o��՛o�T��캫8b!�n��6=���?V��0�*P	\c j��*���g�\5X�V|l0S��$��]:߹`E�������E}I�R�(4(������[��-c�y���"(�X҅�����E^î(�ѻK��+��_��������Lx��~�rk��N�0�䭁��;��6�_�/�< ^Ȗ��:|yK���Y��`Axp��&�?ua��4�pJQ�����	��@�p˺z-s�?-/���egt]�}�+��wf��Y�Mp!vg�/�jj�J6�15	1zg�����-�ٽ�<	b�?i�4�5^���U����`<�fy|��mP��U���6�0�	n׫Q�x��a�����1A����A
�H���B<Th'e�ډ;�t�?��GН/	ӿA;_sh����݇�;?}�[4��{'��k�1:z��
�"e�7�m���@D3�T���{�H�`
k
^՝� �'y�4<rwpu~Յ�`2{ uee���hg��|t�\�t����2�C�Ԑt�b
��^�D	�!y�.��p�{
��.g�R�cU�-������ۑ�y�#?�KM�Z2�駘��Z@J)V�\��=�{0(�ï�*�������Q���z�t���|�.?��ea]��p(�	�3[��:�Hh���	�[��(	�~�^�ⅴ��������Lg�H�6�a��kW��Ar5�-Y��L��y���FPp���f�nhɱ����T�Z��o��~^-!��Z�S��`UP�ϭ9�֡���K�&�������1���@xѮm1�n?�s����h;��� �J.�ܖ�O�l �z�5Y�8�u������0�?��Z�etN���i$�\�	�Nm����6�8x׉�BM�w�JѰ1`0�KW�:H4�Nlm7W~E{70�}O����0��	!in-�O��;�)	o��J�f�LR}z	/����4ޣ����(Eð6`'��E�0�S�㒥�]k��.��<�+_�$2�Mg����A��:K�+�x�@��G���q��-�'���%z:�t�(�>@ eiZ��nd���|j�8��z_g�/�i+Cr����4�(���<�&�3� �p!��kp>t]�P��#Q�
@Iç&�,k��p�T=�cP�=H*Y�$���P!�����U$s~�5e1e�Q&���Y���͙4����럿<��x���s5��O����G}9��{�����''�+����>����W��Y;'�&�8?��B��mɈ1��|7�P�p�_"C�6;���_{{��w����:N+Z���>L�?>�q�j�e=���a�z̴p�|�|�~��1>�g���>�xtr��	tu�S��?����:�P�k�|��l�c9�kS��I�;��dA-�n�>=i�=od��z�,�͖�1�j���\��8U�s��>��p��^�Ì!��:��|&t�LV�!\���ӴP�8��q�L��7,l4{���S��p9W4=k�WR7F����: t���Um�8y�뾧���0-߫u�9�jb�㏤®�M�A!)�"�i}���ۏ��x�&�i�38G�q㫨:�
�|�Ęf��q���О�*��AT��I�!��Όxbg٧~�l\ �|6{�@>!c{jpJ�U`=o7ae�'~��PPdx��@���� ��oo���L�
�D;����D5gٱ3��A�ί'�z�J} �FL{�9�)#cB�-i���E��AY��O��W�����������gB�s�mm88���a.�f̺��1<\_L����5���y�Q�������1�tl�9�q��� �%�:}f:��3(F�*.��i����;�Omr��M���LI-�� l�	���v_�C�N�u��B��0l�����O-��U��Ni�֛I�嚴#��c���>f�u��E^�>?��J��ar��o��"�QS'��Qm,�~��?c��D�~SU�C�eO��\1��Iiȟ��䞏�M=rVrȮ #q���������ͦ�M^���M�F���_gb��Ͼ��Tj�p��+��_�{@l���Gڥn��e;<�W͘O�����4��z"?�C��P�cU����ZgĜ/�����[�^�V�˶<[�X�<7T����Q���:�|��d��i	��Z�î�#��}f��=��9n��������{Fz�9Jg�����	�U�h���W��N��d�T_�x��jd&�̨-W����Ji�3i�%g��9�1�����6e<����t[I���,σ�n�釅@tY�co�˗���)�YL����yǢ�5i��Bx��@|+����'+ +#�̕�Yd7Z�*�Hg��L�د3+Ε��AH-�*��C9C_�t�cj�UB��'����1�=�% %�� �^��퐳\�_����M�}����T�]���+�"V��ES�$'���;*fB8���	�7|��:~M-V�������VN��O�!#+l��2�f�������:�a���,,r&{~a��b��gw��ȉ՞�z���z���@������%O�N� ��}�/�	D�! �M�d�/��~eǙ�Z�q�i�3�?�Ƕ�ݼ����V��U����@b��(�W�w/�/{�o"t���=�IQ���*8��+�
�-���#5$���oVlu3����U�����h��ح~�������gߊ�iٗq��ᩯ�5��jo|��4Y�}�e���L�t���M`�/�UѼ��N�<	f	��!�1 Fq�I���IK����:VXY��~u�v+?�&����V�.�נ��l
F=��i�5"M��/b� \)�+����S{�n�O���k�~�bZ&Y�����x]�o���۫?����Tbh��`�kZ*�@���4б���"��}�X��U��Y(���a�K�vU��8����X~��ɡ�:|�2�AV:�.�)�KJ�����+��QǘX��j��ט��B0�v�%ݔX����zI�����1�>I�*v��N:�T�S�>��}Fc��~�G�d��Q�U�,�m�O�,\ɯ}A>�My�r	4X��M�|��}�.~������䳎�UA\�/�>ԑ��w�v\��3$�֥%�3�Fa�%��tII�2��a�b��6���,�=?㱬r�-"22�#%�����m�.4�_�2���|e"����\_@/��������C�d��C���ȴ$�۵��{�8���Z��dx>����9����ۼ�;��2ۖb��HǬg����Mj��#���(lE�^pm_6��шL*�(40�W�ǯ�=�/�"K^����?Ȏ�Q}�i�rQ���r�Ja��pJ(E(�O�èˤ���?j��tɻ*1�3CQ�ǙV�f�Xe�7����4X�M��zm��N�;1A$��X��=�L����h$^'hB�j
 A���+%I�X��£}D/dl�,�j[tPRHB�N��u�9�l�����1����4�_����ev�o�D���P$�PXL���ZiJQL����Tr|�;���1Ӫ�e.�-�d��7�S�6�Tj�s#u`�a^Y	��o��va��<�5�~��Г�	�L�E�\�a�W�D���ݶ�M�g��P\c�,-�أX�ƚ)��`��!/\#���wC��Ċ ����eb=��<*�-cp
td�u?ɕvO�N���v�1�jgEmyE(���\��a��G�Ω_�Hˇ�v�
�X
n9�hj9�I��5Q�z�l��5���>�j��A}Q�0�j+�O��PjȆ����Ga�����#֑��s�5��$�7}C�"b&�Ol��'
�DՏC1�� �j��C�l�uGd��{����8x� ��z6	��nTc�ρ qr�k��ZJ�5X��A%�=)���}����ȩ� p�c�rn[�v�8n�j^�@���`^Y�3pxe}��ez�1����Bmi�֛q6���)�я�g���G�+j�}!���aixW 1�Vj��m��z��Ї���,)i�1��k�JdW�
;&��m�Ѯ�l_6KE���yX��x�v�����2�p�\�A潸��P�\˩��G}ɳ�Qli��m'��p�E��хGNj��f��e�j���1�fim�� �T8��O�E����˿�6П���B��q�='��������
!Q7E�4h�b��e�Qf�Sb��D	�� �J�m�hj�Ciq�����\�t�3���6��H�l�� V�c�m�DK���:�]�i>G�L��^��_Cy����v�L.�L~t�K��Ӈ�g�t�C2��!g��sdK�*j=3/�*1;L��<��=:�|��)m���4@�����"W\'h����-���{���c�y.�9��d��緋wTeM^H��Ik�m"{�����ph=Ym��ǩ~���yD���L#9Z[}�z�����y�W&CE��u�O����-�.�pð�/�N���HG��N�~�$r������%2 ��0o����C�B�|+ef���8��L�J ��7Yq���t��om^6�K}�>wO�X�jq�_(�z�X<�@"�C|5��d*�rl�E��[��ֵ����$���:C3��X�z�F��d�<Gy^'���L���
]]3Ɨ`1��GTo���2���w�e�hY�>/��^&����CGHA��1��&��9�.�e���B?mZ�cnS�����P��,ʮx�Gm�yMh���%��n�d�Q�,����/��h<q�ʹ�+nbO������1�L��e�-��|<4��a������@3�n5^w��o��PQ���f���ōt�?�s�:HKvf��y�2��M�1�$���ǝq2��qg����W��'lфTӇ���Ss�x��v9�cL>r��/S���W?��Ƕ��C�#�_=�G��;�=(&V�>={#�E¼�=Zb_�L}���UB��j��x��$����6A~�Q��K��ݩg[�dU�Si�9���w,4s�"�������D&�k�μ!�-�'����\ӾE%�.� FG*&�r?o6?��Jv��ު�3A����x��k��{4P?�ߝlm�T��.bF"��:F�L2�:�st�Q]���T)w���@S�T��u*H���//߁^�Ψ�@�b<�e1�>���F5�U��=C����p����+A5���bk���*��⯳�pn��H]۵���N"�;7��dq+Rܫ�6gM*���M�9�s�,�$�A�+�fW�_�-<�?���P��t�C�N�=�a��|�6i���׽�u�m�0>"["͔������Wvg�P=ƽC�L%�%7��G��Z�=��v��v�h�;;)�٤��0�T��C֬������᱁ý]ب�y���_�ɱ�ԯ͒�{�����[+=	���p�%�)����Q{��b{���F����c��&n6w��� AXZ9�]�ܝ^�p�}C}���.���}�$/BE��͊d�� �5ȟ7.ܩ��� Hʼ,��[��[C�-�(�P����QQ�)�G�#�UpqJų��s�����k9mI�^_�]�b�l�iz%h��]���)�BYH�[�X�ZɄ�o�Ou���/�"�"�����3��,��}'�����{`�u5��H}��"�ӽ���%��||��	.�C��	�3?��h`B>� "�5O�;4�����A�iiE��)D1|@�i�=�p�^_������̓[L-4��5�@��F�)���ZKm|3Pf�"�ƟR�q��8��!�V�*�� 9#���G}XQМ>��$j�^K��B�xh}b�g��B=���A�.�����Hi��������_�`���Fk�,��@�#w��c�m��ڴ�7}�2l�׽l�!eفY��$Z�>a��S�w B�nY!禱IY�qNw���c��HM�r��#S{�M��ų�Xj5�t�������Ƹ*��$"���B ��C�#-D��s��߉��h��0h� ��>�R�����>�Ǧ/ u�o+�%C��.�dD6�����ѕ��G��H�(�ٿ*��v�b����l�+R���W7�e�\���OC�>"���([j�|תM��+BN�յy�#�2�Nc���+S��q��0�3oS>�Wz�Ω��'�A�A�K�k��G�����6dۢ�_ H��n�W0�U��<�Ed���@�[��WJ![P����ق-=�����X���U�qd�X�Cg�؞a�}oӾ�;��ˀ7.��
v�t�v|_.�@�=b̆v_LJD:U�����mg��&�O�(��2S��UEEA��n�|���ǳ?I-ͯ/����ۘ}��ez״�ќ�����N4}�J&VH��f���jB���i%�a���4\5�����Y"[E*�V��v�Tr���36��/�����DB������P0�a?Ud	;U�%^��U���d���m�� ~��?i�&d��k��IHĩf���31t�P΀����[�Mb���ČeS�3�ڵ�~�}�4�xa��GbS���Դ��~��b\����QAվ;��Q�5Cu���9o��ۇ���C�~�5G'[����m�H�A���6�瘫!���ؿ�Z&ܸ��?-�B�ߧ���g��>9@���BJ}/3����D/�2�e����U3�f��Z��1^au�gO�i�B.:���[~
��;#�9i�Q!YN��ъ�U(�����K�r�/T�^���)��<���������V��[�����P�$^R�Z�{I@��p��jc1D�t�r�!i�8v�*�y������ït.u�;���!�� ��N�P�"vIqo=_f���qE�wZNI{�$�FP�C��[���y�l�K{=mտ�I���9J�"���G?z��}���Ї
v��2�F��\F�Л�9Ax�l �� ��Dñgg<�KwK���wv_@����n� �HL�c�]3���"���뭂�)}�bEHDo)��[�Ib$����X�uGsbg����<!rd����q�)u0��]w3�8��(�@����#�(w;��9v���Bz����X2;�8��7�6�� ��r n��T7-�˷�
��"U��Gdn,�x�ch"f��{3�>�Y��*}P�3�%���)Q'��JG�*ʢ`�/������M)�K; S,ӿ �a�[�����qo�>��x�A��K�gV��z��G
ެe9�_L>,���E�#����n��o���I�]h���ta}����Y�i�_5� %�ώI��Oj>�8G�=��6����_��C�By-D�6DoY�P��u�`��QԀ�'r��mE)��1����jn;����9|��@�b����3����M�,|�K1N�Gm~s�R�'2^�{�&�Ɋ>���&Z�0�k��t������C�g���G���QŗE�*v*!���ߟP8a�];H�<����섾^;�:$W+K�CzQ�!ȱGn�ʗ݄�vi�����}@�Ї)bh*1�h�����]#��p��1r`O"F�0K�b��ΠfHi2G|�Y�A�D��	Pg��p�����>�]-�Y�~��A����HI�t�9������}�Wq[gS	p�"/J,�k;�u/a��<.���������`1���� ՆNh����<�ne�\���D��C��
J����ں�N�/�v��AoL��LA�|]�R��ϋ�,�JK�j?�N���R�N�:���}W�h�- ye�������< ��m�$'+UYJj�e�=���ߨg��2�A7��R�����G��U ,b4:��A�+A�n� ]���W@S~Hi^�2�
�"��N�hS��2���"NAh4>�u�aS}˺�s:Z�XDN�7�$sq�w��
�Č0ƪ��;EB��"�oD[���leB�c̑�[�:�"�[��������ي8[F��ɐ�����٣mx�d���L����J�_�g�����1Ǆ������LG_-!:#}m"�+i�C��RMx�o5���=�'E�C(�.|�1�yDD6��Z0�����h!k��Mo�"��Q��Fj߷�������9�+�D��}�����e�^2dH�/�q�XW�U�횐�Q��:A�}���ŋBAp��$\���n�X����k�k�1y����"�s�"	�����	%���1�[y��@⛪�v�`�:�s*� �:J�\��s(�IF٪Э�1�#���Dg�1��x�KǄ�g��ԙ��	�I�b�	�-��2<�d�qu���J��ߧ;B�4\����،�!;���g7g�xa���%�_@[��w`^���
��Whji<�U�&#�m�5�&���Y���˼�tH�����!��w�(�뭢
.n����D(@�c�M~����z�c�>�$q��h�� ��	��a�gw�f/hy����$�B]��V����P$�����-_��)���b~��BYȬ�Q&��b�Ɲfs��R)�l�gg�^�����@����~S��=n�I�t[H���ǴP�R���-6K�#ᒋ-��S�i��v|4,~k;���M��6�Y����ce�rip�kT�����2�I���?�~���p2�}��^�Q���N�1-��s�Y늆��e@��{>��|���hN�"�E�bapH��NaL���:V�C�_x�U�^�$�'��!nw$�ЇQ7�J�a͞OJ��4���7���Dy�I�Slc�c�z�	��"�)�DԀl�]��'�����b?֤��O�*Iv�8	:}��\�&[&X�f<0�N���Y\��+��술VWip.�d�9�$��� 2��m9I_��ֲ8T"U��H�Yv��}���n��ͺ�č���$�������
��5b�_���aq)x�W�	���[�;�W[۶�a����(������t��-�
��:#��㡍�$���o�*�{��%�;'���i�V4��>&�h��������	-��e&�Xd�7?[R�V&1��!Z ��Ic5ez�f�u��	�R���j2�]lK#Я	=!\��Q���e~�����T�-\��!U�nף�}�y�qX)T�l��.X�V�4�@YI��4Ў�R+�nuqг�*�@��<V�1�a�KJP`Q�
�cyj>�k=�����~dC����.�A ٴ'���Ss5� �+C�˧r[����9�=�3힕�٘D ��κ�1���j6��ٚc�a�0��2(	1!K�g+ ��èYc�����q�"F6NBʎ�#�h�B�,!�[%/|+/)n[��ɿdAF����j���Xw��]�԰�Q��"|)*����L_��[t��p)�?o6kH��W	���1���ٖ���MS����|���B�QQ9�,R�|��j�g''����_C�m8��˿�Ėm�(튓��m����+�Ti��> ~7q�`0c��]1v��_fz�o���x��9CeT���W&�*���wc�ب�n�e�$f��2]�5���)]K�8�OX�7�r��xh@5q��&j1l����PR<�=O���_k q��B�����Ҋ/���J��q�=coC���kX�4h���0���U�CyK/�5I".vfr�p�X��V6��]��ʷt��|_h�/h[�%�	��آѢ�'�
�	����9���TP!}cU�r?g�B�RY �9�WR����!��i��������'�o��ٿ:��g�0,�,0����~���|N	�yC9{�*�ԝ��w��ƙ����l?yX\��y��H�vA�����`G��o$���a��)g�������^�pZX���+z�q�g�� ����۱ק+���u7����]ö�{�B�X>2bܑ�q>$?]e�<�<g������I�����ߊT��2�+�oj�(�}�����z\R����������K��q�=�A�I�~��*���s���ǪE��}2}����H��#��٧���/�W�r�)��6̵���}V�q�����% �����CJ{��RV��(X����b@#ʏ����F9�:�t����s��W�Ӏ����Y��HG��o��`E �Zz
��pɁqL؁H�ed���D>��򼅡�D�<Gkc��"��*~Η�k^�GI��J�VȂ��H���,����xO�}��������c m�%:6`7����Q6��BA����߃5v�C�~	8��7}i�F+��o�zI�vB�ڜo�XQ�=�;u:m���ӗ�'[�F	X�^�GL1�E���}�>>k~����M�W�2ϵ�tE���đ�Hz�i�:��ev@0HK��qiY��MP��Tx�c�I�ŀ���oǊ��n|_�ϩ�e"�".;�\(S-<m�!�$���h�DG�J�*����nY��K�N���3}͡0��=��D����)�Z��2�%eq�`��>�]0�Q��"���Sp�*��ZŘ��,F�'�ڙ�^i��b^����!,, X���] ��Y�S�;r��n���̵��B&��@jW�.���1�Y�i{��1ot#�~N�>gA��,Y|�k��ޣ�A�F�f�:i�Е���:�:�q߳ϣ�K�5�3�[:D��t��������������vC
擔L�%Z����-���N'�_�♟�Z\�S�� ?�P���	hb�i��������sdd������;���L�j(���gDT�d�%�q	-�����Ľ �1�vΥBS��T�/}{Hy]c�n��=��v#���%����6[>58#�  ڵ~B"�n��g��� �܄c�r,����
C/�pR:�L�V�j��p��V �=V�Ozɺ��C/?��Q��By�\��|ؑ��_R�rYk���b���GS�u����J�_�����_Ĥ�K=�����:ǃƶ��{[��-������Vgق���d��w �$m'�(�����P��d&�*�+ŵ.t���^I�ZUü��5�!�*�A>�U���>�ƅ��U�vLCh�G��)�הּ����9_�۝�8�_�@��u�ݚ���s�}�&�0�k�w��#E�4���_�� ����.w�K*���?��޽=S�aϽ�#�(�թe���Uآ������|~u��ؓ��F(��+0�����a�F�o��cJ^�ǳ�N te�;�g9(��� ��R�b�N.��u?�7�N���C��T���F�k|�r�X1���_�?��"�L�P��*/|,[d%������#p�s��k��D�s�rSÔ�(����7a�Q���לk��%$N,�Ś�r�Gw��!/�Y�i�>��Oճal-��h��\ާnG���#��qk���2s%��;kg��y~�R��&d�+��n�������;~D�6�\0���Gɧ`���ʴ,�����2�A�����9Z�,>��{��w� ���Uh�mK6�P�v�[�Bg�cS<���K{�j,�4/�}��0������cbJ�6q˓"����^/�i;�m�%B�[\� C�XD�a\�݉d�NUܱ2��4یM�ݵ�L���P0��jD�F���Bht���s�0'��v�bwp�qẵ��o�*��Fd���|c�H�u�uF�rvzW�5�YSp#�Z�qXM��?	0V�>Hx��;]Q���A�(��R�~�5^��I�6J"���Ä ���> u'x�Re�[I�C���Z��P��՘�*Ҕ��2�u-y�7ETR��D�����b!
�}�a:�9���@
�D���m���=yM�^�0>�lϽul���^�B�ږ��iC]��wE�Uz��Q��5�S�g�������n^���)��"b�N��cY͊�
0��k��/o�̉�9Y�L3��L�W�|}��I9�-Ő�������M>�n� �
L�y�O�d����e�Pt��S`����>��F�	��*'v`%�k���#<Y(e T��:!.]��{�v���굜��|�\{��	m.��$�1Y�e3r
򢏶�N�Z�t����0²���%G#f�v��_�*�$.ޞ�s����ZMŔ���f�l�?6�{?��p�U0����B3�#TUD��l�>����� ���s (�8.��%
YZ���4z̟�=��-it��`���ANA���J������Z�!�^G�|E>�J{�q%�F=�sX��a�3���ǯ DWT��}h2����8C�f�X�g���A`��=l��8�ȫH�����L������Z������@��ǆ)�,K�E�zU��
���r�f�WP���Mڅ�*�9����t5��#�t���X�� ;7�oӶ�j��B����#��7�ƃ�X݂���(B~CVR�����=����JnFO��?/y� �=�W����I��)hu�4�[�K�m��r�{Z�HM�$����$���e��.s�\˰��Z_@Y7@�����-�(�,�Ro���ۼ��T+��G�{d���]�xzv����8Q�A��}cX>�H��OO�Ee�6E"�67���	Nw�~�ٵYKG޶���iA�ǬU���e��\�b�?�X!5�VFl�S��_p;8�O=IK���l2\-#V��Tƥ�:�rtb�^q \�l��s�0C^�Z��J{� ?�"�$=���7��77Zo�U�I��+ϮC�M��a�k�6J�������-�,u>�"pE�	�H�۠¥h�,���v�qG��`�iU�~î�"��s�ۦ�8ϕB�5X�Z'����jϞ����J@S���"��S�������@ˌ������[ȋLg�:M��u��a��d�Kk���6`]��3����	X�Ut�_���]X�����7�4��#:��n98L(j�Ű���M��5�����Z�w�A��bh��5�!	o��yެ(m�� �1�S�8�$�1UB�(� G@�ܫ�ո0��;��,�h�dT+>J�L!���C6�ѭ>K�*r��`���b%�<I�\�/�����s�'NQ� �3z�38��=ӣ���oM�%?l��+��Kڏ=,ԗ�fls0l��g�lw��_ �v��
"�Zy��b���,��r�6q�p�n��� q#�Ǧ�xWeӱ,`����aRt���z�Ei�w�1!e(V P�t�Z;�ah��Ҽo5~FL��l�P
���Z��t�W6�$/㈶3��D���Y��`2��r��|���=J(�f��i�m�B���ew�+p-xN����4y\��+kV1��(��6l�*��+��Z��6;X�H��Kx�<G!n�B��2aW1]�v�1]q[�a�D5G��Ɉ�9��ĥ6�{��)�˺�� �����'<a������>f�i!D�L+��®��ԝt(/�Gsn� �'���7� B�3��e��2���uu�o��Ob�pki���CQ�Od�b�viN�ͺ�;�/+��;�_Z���u�H���܀��]���Q��#�f�j�[�3����8U˸�u�'S�
o�7�� xӻS�}��G��"q}�O���_<�,D��Łg�踞蘾���k�]E����*pbE>PZ &�bF�����<��FN�8M7�`u��hX�N�r���xpp�Yaǯ�=�Il{{o��cS�k�)öp��>��:�)�<�Vo4�s^A�!&n����{��AR.���b��94��/�
�w���յy@��B����^ML� ��kN3N?���0I<�L䖡��pc�+ ��k�W\m��еelE��Z^IP�XWoPRr�������#ׅ?�f���v�'����B�q�Y����7��W'���@;�w��.'G�s�j�E��4T���mi���[�d�1e[���~�j(K`W'�����?�j�@��!T��]d���gk�E��I]F���MJ:��o�`Ϧ+M�WQDg�7H��� +{v�i�8��]z��QE�b��ם�E�~x�[ �q��<�=���L�fY�7���}�t 
A�:A�-h����RM�B8�����}̔�%R���<��"Vܯ$x�1t�@ē^d`6��L�7|~W�V^���Ěݎ?Nu�� W�b�����"��
�g/����W����_?��Z���<��+���xqR-��v�����*aZ<N ��|VM+�w�� �Z;�Xc�%>����d�yu�k�|��/������3ٛ����=�g�GD����KB'l��y������d��^p!v��9��c���y��Y�
�&�=�RaGr�"$=׃S:ғ����>
L_�)�U1�W�m�<n����1'��%����$�������c�M�J�G�L�IOF]S�s�Վ�ή�C_����Z��NH�	� ,Y}�~.�w>
�haς-U�_ۣ�E׼a��3��P��D]dz������	<��W-�}O���ٺ�ū�����v;���.��M�j�G��z��p���vKH�����̈́6!H��rt��g����>e��!�{n=�jj	����Y�z�ќ_�Ni���l��I�w>6���f�޶�a	Y��{@��ݖ���oK���w������h�<~-ZZ'~��Ǐ#�1�r\˥7E%�]�r0�۹M���Y����r� N�z_Z���՘�*�+��!��M�u�.�fԿ��G�U\d�p�P�r'��������O���9�Z{�p8�u7��x���0���5�ϰ�B�ݿ���wuH)�6�a������٢G�mԨ.�kB���J,e`	�5�,�;z#0^�G%�YX��)��]�����vAX�Y��e�0��F�V22c�Pq�:Kg��+2�����#���G�O��'���?F�8�G*)Pn����%�qv>�-�lz�ױ�u��9v�h���tٍ��C߉�r�[�������v�\��35HB;
����>�ȹ {�kŁ�7d�>d��T	��T��$]ϓ۩�;/��p��WæWS�zm�"�$S>Q%B���_Ѵ�9��C"%Z� w`�ԡ�o�ߗ�&E�岅��	��2��JZ���*_�����;^���"�.�Vr�ʛ��"���>�	��8������P�@o���O�#:��!�7,t�ΣL�Đ*(�Q&*�����j�1?�/����t��<�`����`�!9]���E���y�G��oDy��xJ>�v{%�c���`3RZ�����c#{Q+��]�~��%ܒ�v��ݏ��n�T�B�^���p3�
K��2�v��V��d�)&���ծpA==�G?�
�sC��i��T��F>Z��NΆاr�=W[3���m��:a9vň�E�i�0�Mc��u[����ʽP�*�XM:�Pk�-���_�8E"w\��B�F*�n���b�!w�l�=�����w*b�ekD�B��|[��ey�E|M)8��7�G*�BDʨ��ĭ<���?�
F���p�*��k+�)St�U��t:|(�6��m)�O��E��Q+��o�H���\�����a]vkv.���W��n�危S��>�B�����F�%5�*��j�v�˳G�(��$E��P��0+{�Z��H�~5dϖ,��V@Tv?�v9}��UK�~�X�F�H�0��V���2Yb��*�#��@�:�_�Rx��^��7t������j��0|[��:���BC�evxʦ�D�r��� 6���kR��k"�ބ�M�������E�ŧk2��8Ŭ���6���\N.e6�D���[������u�\|E+�>��*o�V�k#s�8��WQ;�i�}h���j��\����s�UX*MT�ԿVm�rσ��1h���|�R�lz�G�F0��R]��ȴ��U#� sM�l����ل�2�~Z1�w0��T_��2g���8���(Ε;* *��_�.�jhR���D	��Ƌ��SX4����!�݈�=�c��#���y��S��k�}[�`O�>����!�=��W`N?��h��H/��V�Q�����Z"�ҥA �%/�|����A�x=�Y���^Z�zB��ZQE���d�#n��L~S����*T1t�ȼ��^��,��r,>?3q�ݧ4@����1���C�Ae��q�^����z>���~֛@�A�t��?�
DM�_ԙ�G�\�P��u�dg��m���óS��"��+d@��j?5�������˝������I��=�5a��2n��E��L�I��]u�W1�&m�ބQ���ա��R�Ϩ0���{�Ǭ$>(!��Я�Ɂt�O�<���.ZN�ui�5�::4LƆ���M/6i�`��s�u>��,ۯ����M:�N��W�`v!�К�8���Kat�ϣ� ,Z�~Ls�P��Dj��T�$��U��*}�As.���dI��hP�0�nx̝�V��$�bi��i�'�,�H@\�2��BhC��9�QjW[nqA�g������Ꝇ����m���Ra���y�":Ʉ�����3�a�y�ʽ�X/Q�n��b�sxD�P#�H4p�_���?��Ը�W���9����˭�)�T{�Q��N�4.x|�� �����Z�m14�炦�3 �J]�����(CŰ�=��]�V��;
�'΍���L��aE��(�ě��5?������j]fTk]�׸�M���N�����霿�X~�H�]�b��P�Y���$SP|�r4�2�[V�Q��[��܃|�7���P-������3��V�%�I�[0r�"-py�0�Gh�?Sm�(Ug ��1����þ���P�8S|I"��N��tS��:�j��{ R�~+K��]�n�ވ������7��Y���8O��"ﱘ��#u�<��Dܳ[�.���mmQ�;���\r�@B!��8�rV��[�|��|"�����5e؂s�S�m��	��܅j'�u��� 0�mo2.�l?���Q0��ћ/��rў��|�f�ݘgg)����~r�'h���kv�/��>����Rn^w'lL�:�G�ێ�g
��0)p�ͣǒ��ۼ:a!ʵw��M�<���$`��̻���ǜ�DfQ��Z@b4���焪�]y/���6�~᷅��0����Y����.�������aM�q�0���� AB���Fi%�%���"�5L@EEZ@@@B�ѣk�tw�Rb�6z4�k����7�q�Rw���'��y�, �A�'�d� 0��Euef3�ۏT��5x+�2_S�7�X�}77Wv�+���ϣ��8� ;TZ�r[�!�D�ʠ= �Q�����߂p'�޲BZ.�bCG�30ۖӖ9�ؚEb�j��F��	Z'ʅEG�8V{r7�O�W��We�Ǎ�O屚����p'Un�7Xi�u���Q(���
�n��&�}����b���h�?Ka�N��a��ɲ�5U~'Z��׻����M%��`L����見�pt#����ʏ����;�:�׈�Z��'��fO���1֨d������,�/��E��䷟cq���9�8�N���,��,�����7l���:�.P�f�S��ɗ��Hl=����G\	�x��a[�����?*#E]G��.�l���4�� �C��W����Z��y��G��.��.I�olZ�H����p�N#�c4QX���7(������P��667Q);4�I2�h���f(Z��5N����OI�f[y�����/m/]Z�"d7��4��$�7�E�<W�!o����G&�Y��]Eڣ�H���7�����2��+�V|�|N{(c]I'[GL��)���4l7��F}Ĳ|s���ϟɸ���7|�o��m�njT�ʋ��<$�xs�� K�2�{YIe�Η��r\PJ��G�t0�0i���\��%kv�9����b%��c b9�،ryA'{����͚-��[�N����R��]'�@f�vK��b��Ǥ�2о����ą	^�e	+����nE�v��$�6���V�����E����ƼT�У.��4�u���:[1�������C�㐛[^|�!H�)'G�E$�D.�����Yo������'�hRq(�.����鱣�q���\[6 H5/��Z{���6���@���PP�ˮ�~��Nt^̈���/���=�n��Y��L����ו�*yͥ�;�p�y��6��}��45�²�O�����]w�}����x6�Fk�����0+�L��i���h�}L?��4�i���V]ǀ|I���� Y����&&���noQ�)��x.]��ktj\K�:�g3�%�v( �~[��#y��	!�z/i�u-(7;��d8��8������;�׮_�c@9t��k��au~  ��_�~�&�/���F+�C�c _3��JqG��x���߻ͼ2���H/|y�	qy��zM�ʬ�	Er
k�e��N�'�iZu��S҄R�ٵI;\m����\�-����}(@%dc�R%��u�B����2Gj���/��O��R�2=����7�Q<�l��d>��n��I��[�� O�u�P]_bh34�N�s�'����w�Ls��a�Z�M.+�*�qV
1a��:�܉4��
@��jpWN����e������{Y.�I������ķ��@ꉓ���\j�N�ЩsKg�$[b�L*��P�����Q*�
ͩ�+�G�,�V�[WkU�F����z �Y�I��1E_$���X�9^�S��gRW� �%�H%dw�NG�,���O
��/g�2���y���h�P8�(��7�me���<����P�/ܽ�_�o54ЧW3n��������)R�߈!�CFA���X7N�5~
>2���/]A�N�Gw�m\����}ƙ�Hż���M9�mE��<Ù���%�n���]�z
�y�?d��u)N����p&�H/������a���;�o@��m�^0=���\`G
 �|hN�o� \3YQ,6��8�s�c$脸���@ƥ01I��^�0hԜ�X( í{�y�t�g��d_q��e����M�:�- �K�`�s��-N �d���Yp���]�����j��%>z�۔�@�_�&y��}��o��k֌���(���L&Q:���b��0�A���r���
��o�o��`s+�B�2�ʬH4���}�Υ����z!�e�����[�[��"���1����o蚵[I�N�R۝�n��e�R�Ӷ�X�tY1�ת�nf.҅%��v?����$^��L �� &@�̐�����*o��<�cJ�$�C��<�sA��`ho��)�ad��(B����-Z�13�> dv�_<Ox�OpA�
��3��]�a-�&��1%nya���\v���m��r�kYe�M��0�y\�ύ��=> ^��	hMO���z|��&�oIsV���>� 4$�FJR4��x̴8an�×�s6��AfO��Aqg������9:��z�T�$P�u��t9Ώ��i���Օ������a<]��ZW���K�L_s>����n,i��M��ҁ�[g_EB�_~&0�ˬqZצּjM�W����Fꦻo��~�:��ښ̳GF�C-{��A��?����X��xI
����2�K��ޱ/#�8+��B3�NB�4d�{��HU�C����z��	!��v�E@�(_{7q}��}nӷV��^��7�|�Lז-��4AML��3b��f�1V���s��Լ��d���,+�S1�I�p^_����+�c6X����GI���W ��c�71Z��q�|�0h�G�lÛBY����4^.e]����z��,�='��5Kb֢E���+~�Q�b�)�|Ҕ! 
�*6#��<=��X��i��9H��d��T�Q�����9����*��N�e��U`~��L�+������*t�x5l����]R�l��@Z�+�M����#%GW x��Բ������� ֽ$��"]���]0nkd����qYDcn�Ƃ��q��\ ����)�YUs���	��ly��^w�3Δ4�j�T�&�s'�L�f<5����,Ǿl���i�Ahn�[�ڭ)����.L�H[��5�/tfveo��Z��rqq�C���/2����3�:lv��!ɘ?��:C�
�t��d#76��'TCUR�N��Q��ܺ���餙R�6�֔17��ַ���P�%�M���inO���{�ي���'���	��3#����1V������0����2	��������O��˼(|�犙]F�m�ǖ�+���9�B��/�e��Y�.夏Q�vɯ����<�VwҒs�!�z� �]�ԯo�x�h-�[^a-q�4˚�on�ѧ����P�t�5��Z��&��g�Vb�G�FO̙��nY�v�Z�.�_�������q[]�%ճ���O-:� 43M�b�'����/4�%	��cc:��WF�i*H�п
�Rn�����?UX�I��S$%&��ݚ������<��;Ah�"� ْ��9�ka��ܠvw�)3{p�~�B�1�t���lI(`<���_m�Xr&2$:��-�A�zG�k֓0�<�Қ7G8N�%��lW`�ޙX(��H@�6�kP�j8��wRdtZ�ʺ�i��������%!R��idM��g�r{fۊ%1P�[�����V��c�VZݭ�e�����r0Г��y�hٽ����?t9<>��������GV��A8&0�[����`�j����볇<"�p{I�J ���g3�u&��������G�L��	��JV瀄�$zT�5��ޤ�E;�����K@�ON��`���AzP��q�c���}�W|���_|Z�1 �]���S�LFV�vT.J��o+����V�c�������-J}� ��2���-$?&�I� ܬ\���>�B�}�I�N���۽po�y�h��-��V��Qn��꜅R�#�+�ݠ���En��#b��K�����Zw�f��}cWrK�/D7k�(���[ķ���c���#��$��8:�N�X�LB��b�D`r�=�_�4=���̍�����w�\��].�100�E�i��J󅹢^Ӣ�c����=�,��m%��Vp(��xR��֒���OzY̋b�O�K+��|����t'4���*n� ��=n!���0�����(.Sq�S/���ˇ|�PXZ�d�k&��[�oہ-�5�~%��sY��� ��đ1�Wn9�F/t�j��F�����R�i���s-���0,��2�V��6�-Fiq��_����m5sE\g�D�eךq[�r��`MG��X�}#P����*��ԅ�Sr���*W�i��Cӳ� z�_`�}�PC�I�h��`.tz+�|��|��3?�F\/�(���}��������
jfQ	(%e�*�m��?(��@�$��Om�g�7j��u
��Gz.=�ta|2.P��v�Ί��::����"� �01�]g���R<����f�i�}+� ��W�	?3ӜXny�	�n�v�<��R$�"[<���x�W߲)�7����ʼN��7'L��H�]OY��;�Q�$hm�~�o��R�n/ǩb���]KD����%�~���ߐ��^��~��j%��Y���ڙ�ė^�Jѩ��A��Z�L#�$��w�C�;�$��8���x�h�-C�	Cͻ�����4> ����ٿ�����Y��म��e�󻓔I��i�8z�~��f_tLzϗb a�v��+���]��1+�s��6V���V@Q�-��<�ԣl]�|P��������B&[��%M+X:;;��O�<��E�z�,Eʿ�O<,��w�\(Π�[=�� �[�m�?����Y���k����n�G�}( aK�?���,2�Md�/
�o��&6,��X����(l�L�SYэ��h#�S��&}%B.漐�ч� ��O�[��ԯ2Q���OS��,���J�A�&�'+p�BbR(�>� ����|��$�\�m��x
�Q�,;ܷ�������j��c0d�l &�eg����l�s�^�l�d!��(�����5��U;2�H�FT��F�!O���-�WʝA#G�d��H�����B�WY����4�.��`=�d�="�y�*����$~<�Vd:ώLV�!��xb,��Mn������1'L��Q=L�9�דϱڑ�n*ja�a&=�_+4�.P$L��1%�	���5 
+��Y�l?2&�J]����ղ�;H��2wR�l�����X���� �������U� ��]�K�b��j�R� �O�fP�BHsJ��
˫p}*��C?d%���ߚ41��v
��w��	��B0� ����[5�V�)T-��
�w��K�eOG��$7�JT�ʚ�
J�YQ��ٹ�>���ϧ��]��q���}]�0�S�&ѽW���Ʀ�ye��DJ*7�a��߹݉�	��G����(�0�դ˖+/�@s*:���o)�X�'���bo�=�e]z֜�h�]����ų�R�Ν [y�F�pO�í;������;*6&r)X]6\�~��"&��ɭ[�f���ZsK1@��\$�٣%��t.��S��-�P5��*D������|�q5��z���<Lq���ۿ1Z2����?{��??��?��?m�3���?��&�O���w09go���vU����Z�4@1��^8���C�kd�M�hosJzdԴ�h��פ�v��"���8u#~I�'���7ˣ���Q�وl8w\�Q�	Wb�kk�q*�*�IqR�Å�O�8�i��w
��"�z ���t�E���zᵄ�BiW�|T�l\*S�����^|zv`�)�I:D��lF�Ccc��FY�D	���N���7~�a�¼��P�|
#`H��y/I���g�&��/�1O؇%��{��&󌢓dqO��wjaX�2.+���q�u c>��}��MGHOO���B^���	�F]�6��?P~���ˏ�}������������ū�/���*̈j��N�;��S5��Wi�U�h�I����%��)o$�X�'����x�^�Nj����6�Nw�;���wڼ�o�!�e�R	R�/�	zY�P��3<�Mi��5?v����J@o�\����&���n���K]��yi�w�s��Gȩ�����xj�n:	����Q�������!�ĽB���e�WuL��C����ֈ�M���Z�ư�H4�@�b�hg���g8ū��~7�V��^-#������Y#��J����q�$�:5�'z��nyL�yV�s���.�����<!�MW�I�q�g}%^�l_�65?!m)&t��=�5�^�ЉH���|9z8}��!Y��i||����㥕�+>����
�|��Ǭ��Fg���$ŉ��M��d�Kj��(���d�	�_��߇�+��xi]�5��������'h����mi/����;+E:����;d6}�s�XB���X���ǅm'�2�ʘ��5"��>�2��5�]S]k��V
�ʖ����G��<n�?{�z}6H��m����^!�v:�r^z��6kz��o{f����������Z��uf}�{�n�eXn&wSg�ɬ�-�����ߛ�U�m�Bb� �q��VW���0���)���_B����Q�l��_W6��B���^�\�@ؘ)�-���TM����]5a��g���¢�?�������4F�g4����;�3�s�2�F��0�M29���p��g���d#	L0
�ZJ�z�v�(�m-�](I�(]d��I?�y�ڨ�s+������r}J/��`
_�Fڳ���Ò�C��9'OFݪ:_O.�u�w����k��Ĉ�wk�B�n��j]�`܍�移����(������JF�\i���1Lպ/j'�G�H� �R�jXu�G�pPP��x�&U3Y�/��~�Y3	�Ǩ�.��5@���}n�RQR=�X5"���M���afzz�*G�^<�me��w�dWݎސ�C|�;�����F'Ů{�0��w�O����?l+��ZcËC�mO��Ƕi>���A�mY!��^c%Y���C����;�S��پen�\	��H�閑�;Y_J2�X���E��TG��#\������V[D���a-�&�m5g���u�O����
ɓ�x�y��N��Y�Ě%��n�|��ɕ(��� ?���*&Щ�>c��N}���~%>~�A�vy�i�	�L5�������'����YbM���\��XEe0�@�銕�I�Y���"�$<ݵ"F0 ��_����R�
�tEFDn>��f�M�L=M=�_�'į�@u���"���vv;+�&�`��Q���/�h�>!�7���Ք��ƣ*�����s�Qq<��%�U���1];2?����s=3ٻr�qn�(;���n��DH���m��"�:L=�0������w61"�-�����Jt����������8��d;<����~��i�Kn9Ϟ�[[~�ͻ��@Y�:it���D����'�:N6kw���
� P-
����w���io<�� DD��s�J�n���,��R�A?">n�����w.��9��?�S�/H��Y;Eo��ڌ���H �	���'��%��*++M���`=��`o���u��TF㶐0���Vꑗ���9)U�C�^ 㝰�ۢ35�W����9Hk�d�AO�B/��s�n=m�/j��mc��/�M�2u�\]���N��R=�Y�h?}��&v<�����x�N�.���hJ5f�/o�Z=� ���BM����z!J51i;!ȎeQ+���zi�CާGĒ�(F2���4D`�t˱!���З���|�3SU4B�t���w��K� d�nVڣ/�.{i��5	��K:���H�u4�x�n􎽛����O<��Y����=|�Ϧ|+���
��O��b�gC���-�9@��U7I�R�Y(� �^����!��䯺P�e�y\S�%�x�G<��8�zlydtnEd�&�4��T53 k�e5'>䓥�>�c����ǈ��e��V������m������^P�M���_f�a��1�ⰶ_�Ny]��L6r���ن<G;?|ć� n�`nЍ�~�頋�I.�+C���l��R�pPf�������g��<5'I2'
�c�)an�Ӝ����pW�b��~YV�<��2O��z&?��S�єQC-�CL�N�W[LXf`
����߈��>��&�N�ƒ�"�*�HD��%4���'-��o"��yOޢ���@��2qj����Ù�Bi�h�Zb6Y�sB�	@�����U���,���dW�R6Ά��P��7T��;�,=�I'�ꏭgl'3��ݺ�����WHYs��[��a��@��Eܼ4��{c�	�+�M��cN'��y�&u�%-�����Y�{ߊ�Y�{k����8^�o�=�A6�CT�d���P�7:s���
!��	���1ʐxu���X���9��wyו��*�6~������꟝�.s��G�\1:0� ��E�	��Ց$�	�0�2�����ɔX���6x�q����	UF��%�8������W�Wq.-W�Y����>�g�P���] w��>,��.�v�RU9�_��{��� �x`P���Bwc���P!_^R���]��k!�nrSD��*�=���.O>��߉�Ъ�6�L���۴BJ�-�%�m� �Z�T�5R���P��݈NU
P�T䇄>�	ںR@H"zq�^�č� \�>����^e�1+c��XK��#}� iXR��G3�V
MO�f��z�T'u��Ub�U��ah����bdp�D�b��@��'��R����C�O�5s���۾��|�c��}��j��6(�q)BT��+�+ �:�^V}S���7��$�G��ɞ�7�n��W�z�7j_��@(�6K{w�|�M��B�u��Tc+�d��v����r�<U�$�Di�׾��
����[��z�\��7i#3k�2|u�7� �@:��[wI�D�N�Ƿ(��ijNq�v�s�vh������W-����}�+׋ee�T���8�=y:�wFgFw�yK#�-�F����ǋO|�~��V�[,Õ!\�U�;/֙�@eWg� �}u���|���T0A]�����I�3��SE�n����b ���@�N/��Rq���A����^��j��8��H�1j���ݕd�fę�!^�H�%������a!,�#4ޏ`=��v���IW���[��|��4M�%�+S�թ	���7���>�H��z�'�7T�z�����-�(}F�N=��1��r�����-O��t<���v��p�LH0&�'��rמ����Z3�)�Qٻ���x��ʟ��q�d�K�>�i�5kO<�ȯ6u���{|�a��R�Nl��n�S+��@�N���� ��� ���Pҝ���ϐsX^yJEJw���.<�V3�:<a-C���U�Yȹ�S��י��vׯF�����<�N���W|�+��^P�J�����8{���r������ZAI-3��#<C��`r�tsep��O�p����)�BvFi�# q�H���i��h8YŠ��@?,ئ����_h4���u18h���d��r�)(e��8lU�9Z�H�}�WOl@=��|��������z!"ǳ�2t���P�T�k�v�B~��Y�ϗ����������(z��g�<�K�Od3��%�E��d��*_˜(���J��&Օ�OL����+���}�Le&��^��M��a� u Y7�����ȉ%U��W� R$�����-8�0���~d1ډ�X���.O�SQM{���}�CeH�ih�\���+����L;���g/�į�D��ao_�f�aK���������;m	<W"L���Vl��eK���[%iA�^��c#�4��B5f�L�r�� ���Xa�
���>��z��6_�r��hT%?�w.(��+�����[,�b~�Qf/�S��2{�l���XP������s�lQ9��ʿ���b���Uk�<>A͐hߕAٺ�3���X�V15OK��v�e�|7l��!���]Q��e��q�#��h/I�(
�ʳ��v8h7�&뾵��M��m��ҩ[O��%>�}c6)\���ڇ�o(�� J��ԇ�[��i��;P0���������fa�t����������z>�H*xĳ�
v�}����t�U1�ʛ(r���ؙg��2��<�4���w��C ��4������ظ?h�v��{6����q�t� �v�>��=o������pB��V�L�(Q��0���-m
�!T����<��K�M�3�s*_����ٽYI��+�h�-��>e"���!�
H�+$>$�G�*��$�2�3mJD�	P*z�D+��~wSs(2Ll\�Ob��o%����T��^�[N����):�#t&rC�k�y8��l�!i�,X���jl�p�:���/⥬W�֕&�]92�WH���С�������ʯ��1��fz��Gt�a���d���td<w'SN�-e��쫓��+c���0�?�́�?u�B���6Iv~�)<�b(.\���7}G��J$x�Q�4���͌+�v|��A����l���<1͸}�T�2��F�ke
 � �"���6��W�r�V�����~,�vZA���T���㇃?��գ%y��+V^>�-����H���Iq��a6���i׈8���rDs.Q f"Av�~�9�b��Y��R���� �D�d�i����^6�ꇜ_�Ĵ(��V�V]!���ʀ\�M�n
�<,��w#aBs��"�Sd�V���۫��<��!j��D���Uuԭ�k�:ϖ�F����]�Qv�/ʎ��Y��е_����'�d���p�ԕ���� -���}��RR1�r��z	���WH�!nᬺV��E$��sd��t2�����	$ͧ�'�����O���y��N���q�YߍY�&r���*�	��;�Hx�����XH�1�h��=��74��D=\����ưNȄ0K�Uu�$%�g��_)�T�fci8�E*�m��:��c,�^�PhLa���l��W9?�?�����2�8.?������ WNX�:E�W#2�Iyf��-`���8�Q���(��"'d;�.��ʍ�	�R'�P-Dq��7���6�ֲg|�t�����:.k�������z����"ɉ��S�u�5���^Z�Ffĩ���^�./��ҷ��M��H.�h|��0v/����F�j�.�����E���G�#����M"��J���B���qj��r�[�谄������'�5F�]�����>d���wo��6��u��z�M�@K��9�s�f����\D̘hqg*x�ü��Nd��P�n&��`�<�
��+Xq:�zY��U�؄GX�ˡߑ�+߈h���,J���f�1'F�Gx�H�Y��r���3������_�qs�t��o���RǠ�����G����Xm7�)���ߡA9M�h	,c���	4~�8���2��y��� `PV#���ZE �E����_�M#Mhq�1݈�����i~��$�,�!�j�����9_� ������y_�h�FG]�~Y�3�0J�=�7�q �'Y���W$������8�q%�0=�fPV�P����&��>��̚�iɛ|�W 'f�%/��V��0�g� �C��u1]P��ЗC���&�|ǹd�	w��Ɍ��xc'ٷ�>�0|z0*;sXu�������GXPX�8�e�i�]>9Rm�>(3!���{(UB�VJVMh��|��Ç
���7�����ml'��F���Ѷ�7�mT�"ؙ��p��O=�"�-�H���&��ec#��������?خ6�^F��6�9��4b&-	��>�$M�<����=rCf�P�FW�������p�c�����K�|	�}C?�"����y��PR�u"����?C�?C0
҉�d����un����{�-	�x�����o������%���9�q�p�9�i��'k��҂�s ]��H��% �چ�嗨��i*:�[��O��z��H}��a&�L%]iIW�*i`���]��Po��W)r�R�����d�a�}iO1��])E�����ϴf:�H�ry�iY�PԼ�gm���T�H-�z}�)�LW�Bv���4E��	@��"�*��_�.�����Y�aL���#��.f��9 �􎶰�T5q���! ���̵�U��Ab��: a�N={8G�Ӳ���*����e#��E���{}P~2x�}d/�4�-�,g;ԨR��]z��H�^�O�[C9s��N�}u��J�}Cƨ��UqiO%j� :f���0ᨤ�I�f��.)��%	e+m�i�Co�R~�涍s�8�S���dj�v�����Θ����W�N������D&�2v�Y�8�;�2{&63
�I�D���2��儐�,>�_G��9�z�k_F>�Q�.jk6T�,?��>c(���L�8
�E�b��ρe��/��;L�6w�15� �l����d��h��Glh/%:���;�k]Pk�eq�\|�'f�֦��iS0�����Ę�F� F�BT{����C����k�����і:��o�~.��\����0(���)<<:�UBڼ���C8�#v|u��h&6ˁ)�S�śo2���6����� Z}�r��mc��__	���G�_dN���cX�+'kj�B�ڹ�qҐ��C�p*�W���wM�*z?gWV� c�mm�Z�5:
8�`9�(�:B^Nc��]�C�Z��/e,S{�S�$f��oq��t'��Y@OǨgY֦�;�N﷟1�-3�+`<?5ew5���f{Y`�u]?}�*D٤7j2{����4�p_ٟ�^�T3������
�����b6뙏Y��LJ��E����?�*�ݰI�.��>|gӹ���3,b���A��"�W��?�l��nuў?�9�i���?i=��8kM黤`%�4�
� ѐ��#
���v���O㏗���L�,��lM�A�����>sIU��@!�*N)�j�6�(��Pl�I��į�u������̚:���A���K|��nj4����׾�����~��?��r�,8����Ė�%ę�R�v�����#�k�]�Z	����ᙡ5ΓP����D�ӧK��ok,|���#@oӎ 'X�Ϛ���t;�T�̗���l��$�#�+=�0�f6H��U�R�e# �������tm���q��X��v8c.�0�Q����Y�)&�*��i�XFY17ђW(�Z��{���Ͽ"f[{Qa����^4����V?�D�Tu���l�S�U��A���=#D~J�,��ĝ*���uL�'v�5{�1v8�'E �й2�<�)"b�m��ܲ;A�M6��Ӄ���u�d��b8��$A���P�u�$Rg�/z��Qy��sx���� t3�X4W��@ar.@넕-�G��o����N�+$��W��Ye;\O��`ɨ8���{�6V
�{���8��V�� E��8��4p��䥯*���CV�x���ȏ@�}pn�|�9��u?I�&]�BElCc΋Qb�Ү�u�{ŭDa�7�`@��������λ
 )���,��_
*7�����5�b-���ں�qGEO"#��h ���Zό��{��딕��.��5���kVg4x_!��$E�v.]v��
�+y��
����g����k$�e���Ws5���k���K��4x�P�ə�<�H��Gbq*zZ�9<ľՋqTW�ШBN}12Z�G|��k {�wՇK� �KC�m(V�/�7�n��ns�q.���d���x�=-��hd]�����d��h�B�zl����ߴ����8�Ei������ͭ,GR�)e�xU�N�mnOx�FoۮM�02�ڋWr�'�4��Īg��ǟ%rnZ��`�I�C��E7�9a͇���2����b/��ل+�~�Ò���"�}1���HB��U'�تP*56���d(��r��&�q'8/#u�\���g�$�D=�AD4�&57�3���s���w5o}S�90����P��*%�m�k||��&��L��|G����x묦���}��tz-ũ��oT�@�1�<0=�2u�S>�,�	4-���辚��%��,G�Q�(���t}�*&��P뗑�I���ȅ���u$���p< g��[&8�,� �O��7#�{u��)yr���\��C0>����{om����*��
���+�%߉��'�8���-+�]= z7R����ɑ?z�}h��n�k�^�u+gHeϳ�J��jL�ρR�&w����}9>���)��9'ǽ�Υ�R��>S���,/��q嶭l����ݭ���f�����
{8��?#����{�d_pŨm��S>V] ������"�J��cb���d��O���ΚAIra�a�E���犉^�.HS���7�+���*�p�;��ʦ�g�Z�j���',�T�K|ީ�|A�2�I�y��OVYV�o"y��X[�IQ���c0%��U2�����N%7M$�����j�9$��Ӳ���J�1I��\� JC*~'p&�"\:2�L=}�l����o�Wxޕc7��+�}j	�����g�W�9z�)�M�c?��.�� 7����.Cw����LO�|�����ܹ�*78�;(��=��;0�I���d�@��d�X���Aꮌ.�.j2�%ŖQOCC�Քr����� ����0�׺,����F�t��'�:�Qa�li��|H=[�v�T�9^F�Y����jH`sV�zye�c���*L�{K���zh�a��y�b�xpHg����ͨ[�{F�,��խ��S��P�X����j.�b :ޕ�φYj�� u[#\���]5�ȑ���n���<�绘��g3z��ң��
i�
�H����^��w.ֻ.��/��G����p �U����$�ϡ�W��`�+SoDdݴ�q�����᫰b�����{�,\���_�>ջ�\�4Wյ���[@Iߡ�2](y��+�kiڴ�:�Z/�?��gW��;��T�6���I�Cl^������X�x����E 7#*Y&�OZ��U[��$��·gd,m��C3�8��:n��hEѠzfh/,+>>Y��c��Gyk���z��q\`5���7]Wt�=L�]��%��@N�!����=� �J����^�Q����صci�����X�xE��m���2��TRt����hK~�S~��UMܯ�]����螺����NWO~8��u�{��o��BX�zf���%�J���6�����_�p�W��#w5.h�}���������j�XtWᄍv���n�ᱵ}��E_��?15��>4��������V�M8JKS������m��O�]TN��C�'��s>��M"�b��������ꌖ�e=7����-��5+4�1��}<f��`��n$�B��l�^�X�PYR�g
�6U���Do��5���W��ڼ�w&�U>� A��~J�g��H���%ʳ(+�l3�ҝ��y.�P���F���2S�sk�����W���J]㓜jL�*���+oM���O&]F?�|ĕ:8d�g�hQV����FU��m�tE{�gB�?ݾ�Jį�Uf���i
��;N�v��̥���YN�x����s�ak��[['��}_��z+z����wu��SD|.��<]p���/��It_,@��̕��l��`&Α��a"O���m�}arj�@7a�����)!Q�]��M�M(*�����k CtE�z'�(v|�]�-�(%b{�U�T�aCA#/���7��+����%�lĸ�ɍ�v��_������.
���^~�f��7��_�����J�(�/�ư����Bw�����2 K��_���bF�F^x���\�({~ȩ��7
��)�66�o���W	7��NU��
��^Z�Fr���e��]Y�^Y����:��F	HWW��Z$Tu�kVV��dn�xG�r�LL�=���K�f9&��䝏p?2;\�d���d�Z,���EiJ�$��+�E���-z�鳍�	=��+����f��;�W���W��j��=��Pe�"�ᔯ�F~R48e$�����*_QO���4j �iG�UΨy�7e�� ��]��d�*F
�C��\.ZY����3���[53W廬�0��8�Α��쵤w�"= �'�Q�n@�h�p���Y,W����G��z�L!ȫ���t.�Ͽ���!�k. :E��U�7_ T�����P��6�ࡤ�b�W~CI���K�������t��X�K<��\54U ��ި�{:;�T��X�,g�d"{!��O���^R#M��}�W�
YN� T��R�4'��2��d<�O8U;Fz��(=Pp���`L7��{K�{���[V��c<��/Z��L�s+{/v�_T)���T�X�Fl�:Y�z��sX��O*�ϼ��
�a/.s�R�@�����X��#�;)��<x���~��qg�"�:W�Ȱ��x���pB����� � 0��>%ӧc��������/�3���X���D^�-T�t��/�t���U���ڵ@��,gzj��W��O�unE��k2:9��(-y��p'�{͆�4J���_�^�Yn���I�vԳ�����Kb�)8�ȗٱ:�f"<+,d��Q���iL8AF֍˾c	x��O}�ʥ���j��K��o�Z�=�s#��]Ȫ�j��ײ?ǻ�o��������S�giy��T��.2lmfze��Q�涚��F+���X�.�*�|��T_G��X2[�n?��U�����F-�'�fz0���=Q ��ͦ�E�R9/���u�~&���2	*���q}���)���ȅ�sx
\ Ns�8vVU��6@��oa�]J邭l��)#�8�$�����.M9Jۅ�IH�o���\~��+/~��Y����ta�j���ҳTn'���8y�d�x�ռ����,uu`t��F��`�R��ZM[gSN*'al�#��]g���rj��ϕqS5~��MK�4;�:�;Px��Ƥ��L��z�L>)�����,���R7Ss}�z��R��͝B˒�6@wP�+��������0N�eb��#dK`�M��I}E��Lvgm����*Yz���?�Y�py�
�{ź�u��/O�*�ܢ>k��+�#�PA�wLyJ@5��,�|KWc5��V�-��{��z�LO�N�Ֆ��T=�{��l�����מ�\Y��K�O4>U�^�V�N����<^�-	,�������K&6�<2�+�zL�1\/jM~��ܩ��0��Y������y�������z�2y�����M�em�6�Z����GU1MK��U�Jx7m���u��3����@���`q�_}�BI
����U+p��Kb�R6rY��^#�v�͞��8`7��7�Կ�.����L�e�ߥ7��땂�n�f�UR��*s��pu?�ω������)����`T�WOS���}?QoөM�X��G�[GE�}o��VP)��RRQD	AZ:�c�!UDA@��D�T��n��y� ���]�Z�Z,�?��s�~���}�9wR�W�,�ˠۛ��&����G�"`�P� �>�Cw����>�[���^36���W����y����F�afRO�i����Xj�3I�o��lu����0��{`ڋ�zj��>�I�͑EN��+���7�&��Iw�Nɉ�B��~�o�|t�-_?戄�v��e��HH��d�e�U_����ӕwB�U�eH\�tU����D%v�0�EH������,��7=g_X}0�n�	[��C�B����S�'�{�2
A0"-h��]v�����m����E�6�Q���p�U��	���a���������r�1�ₖP�l�;�y���1~�bI�b��Z�X+��­~�M���%�t]��iv���v/���?|�ǲ�k��}0}�/����&O '�u�œ�<�l�#�R�G7����y���_Σ_����#�LCi��ܕe1K�Fl�5��3�*��L27���9QZ��+�L�RŁ�>��0�:�5��4��6-I^W2�I��"���+�/�1�%߿���c�G�������!�x���N�f��Q��ؙ��=��/<��b�-!5����.�p0�~p���*-�C��V`��8���`�C����Γ�������z��_�A������.��K���޳�V�w
�A��Vя*���p���2�s�%�6�a�ز�ӡw�~�WÄ�����?*5)�7<1?������d�P���x����dw(��T�� ��,X���$}���~�<�?�q=�7�Ӆ�/�IN��09,�_�?���߁�9�@�A����U�^�Zr�}����E��G1�n���@�'�;�8�o�!�����_ʃD�͋�@V]iߔ:DZ�-͆�v��b� L�8�$K��:j�;�Tȭ�R����9���?muH�
�"~�[��"4���Hq;�82J� p���ڶC���P�$�}k^'���ݓ��<5}"�W��W2��uf�^Uq��|�N��4=�&�gp��h�+Vo��V9�ٵ(�I���+�];�)��?]*���'�_\�Y�<�K[�}w�F���(��A����%�b�3���ʠ$��;�5�"_*A�(���Ε�[q-�%zS�Xe���P�o5}�o�7�crq�;��D���`���)Ef�o�kt�������:T��?���%6j��LP;u�WVB��q��K��9ȭ�Y��\?�J)M���c%�{�],"Pl�M��n,�%V'�z��OTU��_W�V���H�?rH��'
�T8#��3qq5T�{���ͫٞ"d�A�t�����*N�QS�Hc~�n��\���	� ���X=�1��xg}F����(��.��;;�DrXBz�u8@z(0<���̓:y�H���9Kf��>���~���r	h���[�*�~�����(�J��J戛�
��������&94����Nڪ}����Z.:��7x�pd�9:��zX��0dDKz���~C�˚�G��U�GȽo���Q�g�?v�&��[R�}x�����s���̵��c�/�{��������ݚ���1����v��_&"�|���+5I����_�-J��i����2��Ǉp�	V9}xO�5=�X5��pl�}"����|�)p�(f�{cX��/��5_|s����N�-�[�ooa�v:�;!�I{\#[�N�P��LoSm�0@/)/'�I	��Ȥ܏����:�*�Я�j��L}��@cM1��1��S�FK@/��&X@W,�œ#j�{.�"�$�Jɰ#r��omy�/���	+u׆�:ҋ�?��5蔿^S���
fJ���Ͼ��s��*Y�b�b�0m,T�S 5�����N
���@ORG�XO��9i���0���G΂*�7">,����֑v��������@�����r5����}��K���ͨ�?,��[Y�0|*�z��s��u��O�{H�^�e������ �5l"��\,���e-=qa�7��|�]��+����J��XL�0a����R�n���-�C(.2J)�� �7m������>c��g�^�'n�b"׼s�ɚ�c��3��7]P����=ZyȌ{F��/ɧu�S�We@ڝĚ�i52��'�=Q��maQߙ$x�Xo}_yK�dW�v|��o"ν�_���jE��ܠ�Q��GZ���:�pc�,�]����BRJ�I��B謄ui�s��F4�
v�������0z(�4��rқk��"�:A��I ��YI?�-8\��c����YH �27+yL�z�|�h��7��z�rD������_��S#Dɓ=�{�4Y�u��?������*�j����w A���w�
YG������g�¸8_؇��{+��P�w̐3�Iq��k'5��چ�W��CW^�1��rP2CP:�Q��X&:���Q�G�<U~I�_�K���������E�<pzs��S��<a�m6,&������U	������RM1�ֽ8a�8��q8^M�xh�D�CR5�$W~��W���?!��V���fy5*��)�~L�KuSRn�Oؓ����R��H�t~Z=AnW��)��S&i�d�6sk��h���1N�'#Vë��$�54��WƵ���(Т��M#����w�{��Ί�����Q�OO��z������e><���x(�H<0C^nT@�k>}��`�l�@�����V {tKQ �VQ`z�X缦��-ߢ�ҷ����M�>�p���:,HۻF�;y*�1<����B���޽��g"b>Y���0<?Y��{N��"�U��y������O�2M�Gu�V��)�����~}d����:[��7(?	�T��C��R��@�t���ڰ������}��́2�2�|�[_�+��~���5��8$��M謎��Qe�;�q����!��1b��r��O�F(}��}xeܟE�d�y���/QV�$6a�=�����_yxU���ە��bz�.G�tBi���
�W�XݴGߤ[�"`�EB8�~J��k�h�?��ghX�Q��!Ng�3��Nٱ��U.���U~Y�fO���з�:��h�!Xg�5_�1P�LA<�}�˩�!���F/�uL����`�gI���S��X�j�����5ź{ ��HC V�ȓ�ޥ�N�hǥ�h,� ���Y?�Ey�^������ۍ�	���lZ��u��S��zӛ^�8�v��:�_ƽ���@Sb�oNWRA����i|�蕎x�7����W��R2+�]����@����Bɶ���x1k�*�������x�:v���'�Nw{k��j����:���	�R~���K� ����1k0(z�!,D�)��w���<��"�7��J\׊�L~����s��B����@p��I��uL�63�T�h�+�"��h�I*'i���kR�s����xo�a�R`Q|�&���V�)�41��l>5A�yޜw/R:�F�1�S����N�vR�HC��t\��y��VE|[��
|t�����o[���#=�)PKh��,��&F���� �Μ�f��O��(9�'��[Oz�����5'��C3_�d��f��eߝJ%�����Z�Xެ˸�R�����@�x���Q���
0dkS`ޑf���ݾm�S�s��%A^g�c��2�1�meV�"�1�qf�v����j,�f���F�%b��)���8<���HS+CLVoC���_f�Mo�74���T$�ݛUxR����;$w�mx���\v��C��G�3?�v�#3��A. �x)t��_$Z�@3c0 ������9�������4���A'�@���܀dz��}�Y�7�*7��L7Ĩ"�;�e�J��F�:Eg�4�v���S+��Q�T,x��tv+��,��Ӊ��[�f���9\n��Ŗ�����DG��W�0����f��<���O:�F�J�p�$G0�:lM�	�M!��r�JzY��wAῥ���<�ڼ���"~A	��u:�VB*}���m껨�g�	/�Go4��ՉG��E\�?`��wd4V
�C)-���x�0I��K�eB<Ü�#���$��ώ������?_�w3`��Ƕ�(%�&���=K<��������h٫��/vew��_�u�|7���Yb��-�<|�a4�1�)�m�
��/���f�x[������p��
�ı�]������_�y��0�)3Jx���C?6�[��ޑ�q��
����n[Z��8��o��:�	��h����ȏ��K��ֶf,o�W����5J/��ٛ��u�?^���p!�,_-T�@~�N;/pK��>��^���l�BtP��[O1���(�v���,��9����y��9:1r2?=��[�)�'��+uٜ1��e�2C�{la�v�ߟX��Z�y-�YT�󺺇�[x�q�珠=���b����)�a6���j�R���
T��e��C�F5�9�Vw�NQ�ɪ���1.Ƽұ��Y�B<v>����q��S/�(�����}�~c&��;��"�O��� �g�~p�l��X�"y�Jü�^`�w��4�p��M�N���AI~��#s\ڸ"c�m~z����H���"E$e=w{����dQ���Cl��[qm��ݥXI��W�����X�VuI�X�V�u��m[�9�&�e��;W�?&>���h��?��_�*I�78=e>�|���s�	�B�8�9�� 1�g�s�u5�Aѡk���j�#��N	^��.���L�P����c�+�:#�6K,��^ޖڮO��"�"��[���1��Z6�s�0����"��:m'͇�j2�/68b����`�����](�9�#�#s4ڸ�UX'�����ee��qE~�zc��网cP-�����}>ъVn���N�`i41�n���.ԹXW�H�+��0>�O���_Iܵ��k�,�.���9cp�o�׬y�Z��V>]NlexE�
�X�}bW�O-YB���a�-�L�P���V�+�󭎩�!@�����=���U�����*�]`jM����ў
��wu��ĢR�H�j>���ʛ{3�Q��;֦�w�8Jo���:5�ɖ�k+�]�7��9�p��5��ŗyYQ��7�xe���J��*+��T�)�1���U�/G�{:iE�YJ/�3�V����e�5Y��C/a3"�,����%�ߐ3>m�BM�D�wD~��[�IG{��������[Smd~1��E��T�07/&�kS@#}��Ӄ����ra������f�O����i���K�AuÓ5�2�^�V>�����������F-�!�G6g�|������EG��jP�1mPTӞ�&,���y�{���94�Ԡ�jl?����s7�|�v'緈���掃4���9YRj��)��_E1�%���g��eTd65W��~�	W���]���͜窩>�rvg1˖�V��ޭ> @�]�B[]�Z�S3�O}�� -��7�\?��q�'G{4Ѝ ��y���>W��6��#ϧ�J�(��� �`�I��*h!P���ޙJ!��p��;)��Wk>��eЇ��W^�apn�l���D�{�ܜl\���fP_�h��Vsy-j��"X���_�L�Z� �h�9�{=VP��@T�2=�s��}��wz����Hg�������Z���2M�����9~�
��U����4�ߘH*0�'H���0����Y3ܴB1W�!��^�÷��砒�1����e�3ы-��OmS�C8�[�~�p-�Z�RR��wϡ�����rǡ%�G������|Z�=@>�e�����6��ig�0�[�c��RT��fw%���,P>�+����^[7V9�R��UIP`�}�x2�=Vbu\չ�}���*`���Xh�~`m�b,�
z���''.��>oh�;��Wϥf�XpzbR<�������\Z�D ��,��c�����l�3#��y�N�g5�.�y�vqE� XmT�M���9Yb�ƌ�;��h�HJ|E"�y�Z���$b[qr2z�5)�$`���x�wWk%����&���é�9 �0~�/}�(X+��gh#�P5��di�@����5�Oy��8����f����t���Rb�rKcѷ� ����>�hؤ���jȥA��+~U��<*g'Ն��0���*�6��NB�]���.���_,��5��}�� �'z�l_xu�ָ�-MY�������W��PH�h�����>5b?@sf��]����ٗ�i�J=AM�N�S�>n�$ӡ$�R(���ICąs`nwL����*��R�:c/^82�gaA��O��:MqM�eA�.$��J�P����0�K���z���`f�� r��˿d�u��	L��f� ^���a�e�#
�u%��>phYYBGU�&V�
ڢ�n?���u�nP)Ծ�yI��|}���Sy�l�)��8�u�毲/A�O!�Z_��-v�a�FI'�R�fڭ���:D�{>x���������Z3}д���3��wNab�i������_]ޅ-��:[ʮj�c!{��Q�L�A��zs�۷lc��D������Wա��(Ekh�p�Εq������:�� �N}�Ӽ�%GW��ق&��F�J`Z2��Y+s�pu��|�R����\i3�?jD�d%1s�&���O� �7ۨ�m'�U;�ټ���%�4�D���64ّ^�g�e�E���T�����{�L�^�3c��S������'Cb�2����d@���rdC�fx�����e,w�|	��Y���.Io��9Xp<)�lp��wb�r��n�Gl`�e<X��n)����-� 龜ص�w2�_qF����K4�7N�x�� ��b���8��8�C�'���H/�� =�m��k����Ӌ{s�? ��_��S��ヨ՞�í��n��TQZ��:�~�3��>c�=	H_����}o��q��҅*^+ٰ��U�ܱDl�y>��O��g��UlC1�ݱ��e�ZgM�&�H4L�x>�嚛5��ѿ��4�S`�����nl��S*��f�>}��wt��]���36�"#�yO�fsk!!�6ٗ�*��h�=9��[��-���^,7E�������������&�H�z�������,��|tr,2�]kŦ����R��<^���U�!�x@̲I��I�3YQ߬Q��5x�:ܰ�m����^HJΝU�ȘO�# �G);�]|����Z��L���-E[m�v�A��w	��v���EI&�V���^b�1��+)�g3)޷Um�Ӂ-=�E�+>3�.o��B�o-i�޵E!k吵� ż��y^da����~�2��f)���Z����������s�KN�e����w��s �Z�0�X,*(A@�y�����u��&�����)h���<�p���*�`u�,OM�X(�-�{���D8�D��jS#L2I�a��$�?r� ��Ԑv�l�H��;t�ϓ<�����^(l�;D�����@�2���Li�"���L��
*ڡ��~z"�)��b�Ƒ���%G��].P������&a<<kM���}�5cЎ}g�1��*�%6��>q#R�5��)���!�����E$t+i���k�p���7�o�}�*AݻQ'��'�G���K�j���9���Z3[̚I�X<�=�XA�����-�����_>���K�D�S����?��[�*�5s=����&~�IFW
��j�{��p��s�����Q ���Lγ\QrZ������{ Tb�K�y�ɴѡI.,��F�VxdbY%�t'�����]���ED ��1A~��)��QG���ϯ�-*�'��e%vJQ��ԡ�! 
�k�'x����/���š�FQ̒����(���3�@�?{��0���w�����Y���am[y(�8,w�#8�|�:Ȁ&�g�Vv���pr��i��5"�� ��_��P>W���&D���G���:��H:�|�/�4g:�/F)���K�v�����l֜ĭ!T
��W�9�٬�!>O.��|�;���׼Oz��.�d�"��:S�{�g+Tv�@{s�Sĭmoq�*U�\�� %)Gb���^?��e��!,g)��=��¯K�#�5T@P� %]�I��-پ3`3����2�|^��7�a�}��Jܡ�Y���!׀�دL�R���jU��lG��2�����N�F��u�|Ľ�@n|̷>V�y���L_��^Uh��X���j(��:�n}�d{�)��t<���l��H�#�g�z���ţ�V�{�B�/�Gݖ�j�uB���!�r���Xl��~�ֱ��=_ג�8V�,n���?���Xֳ�?MF'���t,�o��'80��-�u�1ԑ����SzF���1��M�2�;E��|�2�5B�2���L$�D��LOh��Wb���N��C!�b((�0>Oy�mH���5��L;���^D��_�����c���h�%���ύ���1h/򺇦���`zc�v�PѦ�{��Y2��C��|d�5e2�� M4h��!�fy3>�Mq���q�֑v�mގe�=��VV;/�sH�rBr����:�$!�Y��~�Z��h�TO(�1���a�wov��x������_����zI�	ڋ,�=-V�v]L�̄�zl(`��Y�C���Rנ��<��0qS�!-����db�r�ҫ�G���
Tc�Zׄ���j}�3�m@����vr�.buK�8� ��@���')�ΉI�C�_83��f�D�يN��|�E�
$T�;ʾ;�z��B��aߙF�R:Y�����F�2)x�|�I;�����kc^qR�$�~4x�ZKj���a�Q�6�����$�����x=���fT�'�����r�p 8�ݞ���X�'�At\|��$��7c��F��`�����lk8���6����U��v�&X��-q�4(k�I_&
�g?�~�W:��e�|��g���1?���^��"���]��9϶�U0>��ؾ���F�@v�k���Ov����^��b�Za�����@�e��ۑ�/��cD��G���%Yc��T#�h+�ͲA���3fƀ�ĉ%�@O2�f�(�U��v��ZL9��n��vNy�Bl@�M��I�ݽ�ޓIIr��3;��3��bD0HS��ط�N��6�(���P{�\������fj+}Le�զY�����k\�����uZ5'z4�<�[R`�o��t5�B����᳭��M�Y�>u$D+�L$�-*rB�G�O�H��	���o�O�#)R�Œ}����]m2Kf����
[�W�j�g�Vn)ۧ�8�\���؍
�(	�A��kٞQ8�  ��zt���%n�RQm^v�݄O��#QBd/��w�K��.�	�e9{��Dz<w�S<�%�_�Ր�	�v���C_�+/A�A��t����/���:NLd��+:���W�<S?NN|����ʄ�}c=��31vS-���[�e,��K֖�V6-��Jgk�b��sF0�x� hΓ��Uo�Ks���n�Bd�Ϲ%:6������W�Dh�Rx+�4X0\^�T<XL�l� u�}��[�,Y�E[r`(��,X:��N_�p���ɳ�a��O��ݻ>��.-����,o���L������Y��=.l�\��>^F}��D�tq�`���%$���ΩPQ��Z��]��E��1�"�7SDi|��UH�|�GY�:P(	�0N���\<�gip��t��b��E-`3��X���g*1G�I[�Ү�9'��E��!�pSX�j����f�h���`��� �������BU�tK�0-��`'{��G*�so03^�E���_�ꆮ��>ڕ�����TP��?q�?�X�JQ��F$a�h�#�Η��.����8F��_��3p����SK�Qʈ��C׭�my K�0I�=V�0��_�� �F�����Y N��Fov����K5����jF�U�m|,���	�pse�Ԩ?�z���Q���h���0����<,�|��=�4��mٳy��SG�����щi �`b�3s4�L�R����:��!k�2���)^D�si�%�]��9?%�u�?�@ �6���o�ke�����gȭ�6��h�?�0E���$E<`��0vy�B��] ��ۇ�M�>�Fh-※�Ia�a�zO�-8�(}���/����#�F�tS��X�)����J)A��y:p:� �1��)F5�7I���
���������g�ptíTE��{h'Í�T�Po����<O��{Y􉂑h�脳�dA���kZk�{��e}VH
|_^-�t�|uR,q>�(4{i�e�/�&�=K�:<�v�܅�U%N$^P��x�S1�F�Q4OvϻϨ!�Ake#��U�b�c���&�3+)�F����e;�s��j�[/ZX���ܵZU]�9żF�����nc�Ջ�'���[�J�g�&�"ZO��ٕV�WfτM�L�Z��uܮ�e_6�U2fqu}��Cz�&���K�hy�r���k�E�		ے5+Lh�MÑ��e��Y =�;�$��Q�?������?��|��49 \�m{V6ʮߨ���~$�%R�o�����o��Y��P���ӕ@����T��zC��f��Ͻ/����5-P��X�dBf~>��u�~w{\�s��P�½Rђ�yQ����IЩG�Y��|�7'����e3Ǟ4Q�T/
�ݚ��F����i �
0�ʣƳ�nqϑσ�d�1�%t��/���7��]��i8�b<�X+k �4z3g��'�Ɍ�E�����Y�Q�$�_]�`����2��꣹��˷�<���b a�mi��Qm'�A�����b��a�Ϗ��w�g��QqXr��T��s_ �����c/ஃ!=�W�ܼ\�"70vy��3���0�g�ٸ$���������d�Sϛ�:��-c�Uf�,���C�:����������|W;I��{�i{�������g�n���$~�/�G�?Eo�������ˮ��tg"@��^JHyEY�]���K�*��\��5����l�}[-�ϖ<l��J\>05�/�\k��-�����؝���䠐Թ�]�s�4�5Ņ�kh;=+¡��^�G��nu��N�D�T��~��~����7�z.�dF�qL&j���R�
��,T���k7�KG#:2@g���}&�z�5�x�U�m�i�	&`�l
����efa������+�]Y��1a�qiIv��^��7��u��$H�¡�xʁ7�;�8)E�V�E+������T�i�^�
βŻ^�&K�b&ׅ,r�$U_�`=�Q\�S��=KM�>6��h�EnB_����{ұ��W�uԡ��~��\��d�u%�Fz�v��v�HU���?�`��Y������ƁQP��F�������S��W��#qe����\/�����D}n�����*�37d7�ʕ�x�uj����ݤ|�P���O�ub_���[Q���r�n��Õ���]B��jH�;ގ>ߪ�L6�y��i}��s����f�G�Y��{���6�'�T�q��çvo ~��\:;y����cqEd��f�bz�B�p1��U���{Y�}YZ,)�M�H�y�7�cRo���sD�q��"��z�q�x�� ���?����h�V��{�]4���D*��G��������) ��e�Ϋ	�ل*ɒ����ؿ+Y�*L1�H�/�Q�O�9�_�@{U���1�޳\��&�����a����}0���� `������4�LX��#<E��EK{he��(-�S2Wj��B���[��>�#l���ߔJVB��ׅ]V�)�FD4j���ጾ���T��^��kw$d���4�:���_��	�83�4�5B<Z�up����,���1�9LQ(r�^MV�WY�)P�j���>b��;d�[���T65�� 2JV�K�3���8<��H]>���r�1/ ?n�O�ر.�����Nzt����R���O����W�Pn3S����m��]]���w�&��?���3*������%�5@��ñ�Pe�%���a���Z�5���� "��O����5C�E�B_a ��-rZ'��zMuH*Ƶ�=+�:K����j�y��g�o+��у=����iB��I�a@s����hϏ��Ƥ4��v<Ky��Θwۻ꧓��z�Fp����|Y>"������zn-Y���WIw��+�c�g\ _Ť�rLY�k{���8�B�����������d�z�Kc?�$��[R(Z��9R=zz��Bww6�B^l�\�!��U�� �;�y�O��w˛�?��<H�e�W�v8�K��BZ�A�wtf�;�@eem�����_�O9�.}01�*
�RÌ�,Wj�sJ�YJ��К���)��]L�~��]=�����w�}���Ώ�O�FW�}-���L�����\rpH�2��ր��+�O&����y7zC��> +ȃ���g�&��V�HV{������p�'yU'Q}�k�t�r?�}T7|[&���P��$�$��>L�'�<��
�(_��߯�S��KS_z)�ȇ�GP%FOߴ"�PF ��_�H3l�K��[�I��p{�%�n��.2��p�����١8� �t��E����c��"��ú(�mhW���--�TԎB�@j�����0�W1	�����x�:���n�-� 1�U͡��!�iYЮ$���ڱM0���X�����h=�
@�~�{�jf3}�w]"1��j�((��D�~#n^�R�|Oڠ�=C��9���Qꌕ0��+"�z����'3sd}��Xb���?����I9�u0[̸z ����d�����������өP�i��ux��R�a��O�[��
�񾺖�w*�z�
�?%v�qL�Ƕ�DP������B�,i��E���>����k�Y"q����?Kó4���E��5��I^�8���^��.2��ho<���ʞ|�Q�r8�hem�7M�zͬ��zl	u�������M�ǳ�u�d+V1���"*��ec�p$�����d8�348eyH��J����J5<ֽ�jrk����<�Ӓ�	��U[�t���M���Tߺɖ��A���k���(2�p(<�	@�ee��I�M+�����(���_F�,���0�p84з�R�e�t��)6a��3|yK�y�o�J����b��#����,����@�?�k�2lО�_�O���-��w�բ��u��$.-��⾓&a�o>C�/���>0��p�o� +*i�F��ҍ�"�0��B�~m��i���+*�#n<uc��&��ߗ�楒����//�A�wXR0��w��c܄��=�Q͇
�A�����A��w�XcX���+������������V<�n�t���7 ����X����s2=���BK�,y����h�l�0�sզW�����C��Ä���/�t�R��+0g��lar�gկ��eiӽ����O�q�mk���v�<�<�%�<�hy*-�}Mk��!�V��0�!��ֻ������k� A�eM����<�?�!�>3��Gg�.��X�&Pr���l�'l#U"vt�Ɍ���^(]�N�`)�����oJ_ѝ�����`�Bn��{�9j��c��T24x��L���-FX3R<���^�C_������0�Ӕ[���9�f�Gy�78�2��7�k!4�Z��酆�Gi�Ҝ�e?��/� ���޽����`��y�(-����h�ٟ)�L<��0��]�8]��f��U@�J��˦�~�d���o��ԟa��)T ���}a�w-��3���F��L�A��]�yo�Q~Cl���Y#��x��S��h�\%�ً;+r:,d4�*
X�tM�
�tP�Қ�\)�
��d��l���Ʀ���/k@a�<���p<_�l�NV�l�B[�
%J�����
�x�tz��n�o4�`��FϚX�)ZʶO�34֮��
=�~�e��t��r�u?.Epܣ�خ�P���U��Q��<�N���;w�\�ą��a������A�~�������NaTW���T��p�샳Ǡ�a��6�/�gI?(yf�yOV�ZD}����Cy��ݜ�I�����5n����e(����*V��ѹRɐ��2�rFg�s��ߤ?q)�	g�;���0�2a��&'�g>>�ٯ��S������C����(�;��=�ҡ����~./]�r/�'td(���^~�y�a��$6���!'���(x��n�8נ�������m���8␝"kje��Q�z�$���UR8��L?���}U;u�f�|��'�	5��,>ڒFy�L�{��hIJGu%E�06t	/Y'0�]���ݻ���D?Q�Lhu���=�g�8����<��ey4�3���B*����	��d.�[��������66l+��������-D��j�}���h;��X^��3㽹�#c$6����͔��U��<��~쵘~��ߤ��C���q�q��q
�l{�%l#�������猻�R؁�ԩb��~F�¨�A_@֯JOK�6"AZ�m���'�q��u�Ou��Z��?^�>�l�=(6���Ƚ��S�#/���F-�qȚ˰��/� ��w�,��{~�,�Z;�!�����(s�K�pv��� �?wI�A(n�1��8�M��d��\���P����v�W�G���0ه���jyz���fF{�I�M�dB�p�/�����"+2.��L�ͳ������{#����t�φ!<�cl�w�T0��X���h~��-��n\1nM �t�]p�~ YTgs�F�1�b�'������h�J�<za �0}�� �-dru}��e(Mw$l��M��F�:��$�|���qQ(�`�v�Fӏ�'L�O�ʣ�����p����mh)��ign��<�7��٫ҌF�Z_�4"Lb�,��
C�����u����3��9:t�Z�BP��h���Õ�2	�=h�Y^F�R��5�޲�	�ݫ�l�<���Mҥʻ���|�O��cK�!���sUe�T�_@w��
�H��G7c��V;r�7GЇ�PH����(��T�
��E#��"��7/4P)"��;E��q\H��z��K�e��u(���ti����Y��b��?�ɸ�c4g��\��o�ބ���L�n[4�<l���(=J��B��Z#���	��>�<[V���QY��9e�x\_�h
�_�8�ФzO�{�\>&k\7�ǥ�8/�FK�=:.�%�?0l����=N�/|��s�,��F���kZ���拫-���1�Ay��Y��ppT��G{��)ǭ�2O��w���'$�����D��u0�Ro��F���`���5{G�c���}�|�F��s"C��S���	#גs�R��Y��	9E䲲--��������38a�&����;�e �#���L݀�� ��j��n1�g�s~(`�
���L�>,��ѷ��E�'G��}��!��!`��;'o���_��]λ����Z嗵�5@��ſκ���.�NGLt�g��ͼT�`iݍ�=��xٚK�T�-�	d$�Rv��������`�W�J�����+R�~N��o�]n�<Z���g�����x����@�r�fe���̉I	ј�it�Y6���Y6_cOy��`��Q�����1�f���ᎏq/(��$1P>vc���O�����C��p�.Ӱ4���Pŀ ����"�#�in���F<�ү<����H�m�����}\�������
߅�H��Wq��kx�N�3O�t�i��6<��7���r���/O� ��5H����D������vS��M�Iq�y��P���l�9d�����p���,)�Xޤ�ﱡ�s��c<�I�Po)]Pk���
L�J��{�^t�y7*Yv�#u/��(��_|U�N!%�)KJ� ��g�UZ�{A�j��M12�_�8%�?f
��ԗ8S&c�D�i�@�*�Z��M��V�b��_'�7S����PY�3ӛ0�ú�I�;m���!�f
e��S���#�x5��%�~��P ��� +>&�oX�\_M�L4��{
	ޒ�Eܲ��� -���sV��V����N��j�g������[��X��s^���o���ը���{sw� �<��(ǉ<F5;" `c)V��`a-��pZ	C�fyWD=@װ���� U��9�&�x�OR�|��*�!~틄�s/�Ү���4�g3�
��9-ұ�F�-����h�B�v]�g�)�v��Ȫ���3���}��)�L�h�L��K��_g�{'�8w�{��q�}hR�?���Y�H�����VC����+M���I�vߡ;�ɭ�2l����|�rХ�|6T�J	���2�!i��w��������b�pqC�BU�2q�x�/����~2��N��Ca�3����S}�� q��{��,�����0f��B+1��Q�<��*�N f��1�U�yj��>���sl$z�@�*������i�h5�}��m��<�x�/u��h���)t��9����
�t���b���d�3EF9$S���c�ISxR4E�pH9n�����2ʑ��8r�PK\�����<�aխ[�E�9��� -|�1�&J��p_C5Lԟwh�ݙ�X����i���8axS^��k��]���`c#�Fp����'�VΈ&���>��b O������㱝��OdƎk�[l�����q��O���?駶�k��`�#H����p�o�������-�S��HDa�`=��S�����]�zw��l��;�p�JL���,Lwr�(���X������LЍ��O���3��ih�t��%BM���L����{"�ຍ�z
�~��OKʊ|5���+��Z��}��[�b������^�zz8��WREF=ػi�`}�q|]�|�����"�w�cO��E�o@�����7�c�S��}�73���_F0q����.�(��ge�}^�U�+|�Jn�v��rZ��!8ꟹ�Da�ގ��p�ΪD���;�I<������1�"��v�T�L���qM��.J����x���:<����^M�]�q���QaT�� �HA�n�HWi�T�5���
"MzJ�JP)�Ez�$@�B�=�2����޵d-��$'���{�'�	M�_XM(1>�� =T:�{3��m3������$���G�v������2E�����0c�-�[�C#�rӅ�R�_�[���/��I5٪�x!�d�&�Ύ)ah��M ;H�ޑ���Sۡ���/-\����߈�9�R�p}-R�1P2�[��%u�p�C�#�D��J~��B+��VMf�(�H��s|{0����/�.�m2W��3#f^H=?=qH0o<Ua��L��[������⻌��*�f}��<h��.����$n�M��5��T�QL��]�����}p��և�K<Z�ɼ�&��]�J�اT����^7���qz7Π��\]R�C��D�#K���p��I{���2H��<BG	߃��á)�:�����aIó��j���|�zh��ղ��R�v#���4��o���|�9��'�.�d�`�a��D�h�۩)�������[6�ߖ��}Ѯ�^�%]+�� �+O���=�����o�X��v��?|�ƪ�)�����!���S!�oFo+��&]u5_$>�׷�}ߓ��`o����i�^d��4y{ڜS��y�
$����G���ѓ&�C�Bg�3
e9�el�L�:_l��>����^�5�?��q��f� ��$�_a�ߞ��n�5)��~c�>�Ѫ'��U��J����ѥ;q􊐎;5vhR�J�by	�N�4(\X���`��I;�I�]@܂%Md���T�3�2jE�ij2����/��pV����!v)�O%"��eRA�É��e�iu0F���HW�U��M�7|Kܩ�G*���+�����5�����^:{	0NY�qC&
?qyo|���׈GWb�iAsz��=����臙�����T���F�i5�W!�y�mr�> ᤿sa�g�M�me�&��V���N�I��y���W�%�zG������?E3_k�ܙ�J-%�Җ[��[{��Y0T�E�2�3P�┌U�i�C�9�|, �;��_�n&}G��S|��`�w�i���p3ǭ)T7R��MUuB߃���c��6E�?H������B������_�x[h
�Ȑ)I�Ǩ
P��U��xz��s*|��ы���m:#>���/>���T���}5*ݧN�L\��|�C���%�0��))*/w�Yt����#���B��B�2�=u�G�v��T,�0�D����?bN�?��O�CG޸'?>
�˭�жh$[�Y�4:Zr�B��_`�EDi׹���ѝ����/_Np�LŊJ�M�h;�]�������o�Ve��6������H�'Ӿ�B�#����[zw��4�j|��У�� V�F�P`�H��R�i���s��lg�ZM6�0D5��Yp�0l�rv�咫z�0�E��W�?�Ƴ�V���8{\��n<歅u�.�<�]]w�H�)\�"���@U�?���!��x*1e34�K��V�R�z�-P�j��������Z�g�܇��}���52|P�3[Vj���G;6���h��[��{�-%%m���ΓIߕ?ԃ�fr�Bj�]���C��-���@��e��j���4d����b��߆RGK�_l�}��٠YN��^6����؍��I��'����������{.�F�g�3/��{;\��Ү�C��(�x+���N3��z�;��e� �x��^� �T�k5�~"b�D]i�'W�&�y�c��5��ª�O��[wbǆ��0+�kꝄ�F*"
,�W1ˠ�NxX��v��0��:*4#�UU1F~��<ǂh7=�A�zh1%"��3;���ݦ��i�#���W23���3�oy���d�f
��և
�E�F�
�/�/P��Q�����Ƀ(jBQ~�̔�`����h��f�2�gx�O\�s��Ja��RK��򊳒��	01Qѡ#�#u`b*db�+�_ͨ�t������C�
�H@fu�B����eYv�*s��kNn�t]������G(���%e�	���[owE��6R������R�`gz�9���ֹ�w8	Ɂoi�+�����?�#�p$H]w� s�{o:@-,�W V��W?��SF6��5c99���	���C2�	�@�>���2u5ժ�ϼɲ��8^�W�݈�On��=46TZ�Dg9)�Ε�Ӑ���#M���Z(���`5lTK˟���m������s�)�<��y#��.�:q�':kD'�ų�%�=p�:�B:]���������?�V���5�	4O�9W�a7�ﹹ9�e _���ɂ�����W���J��t˄8��b��n�=_���g4�yMK�W���DdZ�]��Qnntr�����A�T��f��	
�>��3Tga�hܷ
��o˴Z�� ���@�k���Ew�}|Z����l)��FJ��7H]�o�`�/�]zM���([zJ���d�����1\�E���7�H��DB�h���ϫ��{�֩ސ}�
����M	����Ѣ|�Й3h��NF��؛���YW���ɯg5���썢��
���V�Ţ|� |!�o�K��ؾL��ה�}�ᢵ_&�������dR��)��Y�h` ��f,�	w_t �T�J�PT�T&�b�I�g�X�,<����_+쌨�R(�5?a���o@v��
��u���r]�bG4���G"=F�]K[��28^r�k�X�V�bۭ��2���^�@��#�(J�eڀ%5��[�륍.ҩ��l^�!k_/[�^*Ȫ���x�1�݇��9�����?�!���20�͗�\�V�\�'m��WIώd�KS�I�uN?�x��u2�aXf[�FY�`���'�8ot,^BL��xɿ���\#~�K���n�Vj�E�!g��Ɠ�L�j�S�^E�^y������~k�.(C�y)���.��A">��ލ�(��,�3P�}�v���o@��W]��U9���ۦ�Uf�I�0[W�:--��W�9�g�>��!a(�<~���xR.K��M����2������ʇ�G}5���;����C{Z�~�G����t��%ԋ�
��rzߍ�t2�
��Q b��<�t��.ˍFD?�}�gzW�����٥��f��f^D��9R�:I���Jo�4h�n��'�S�,�����1�� ���$g�-��w"��`'Ҥ�ٸݝC�{�IUS=�\H�P.,4v���$�EE� �{�4E�������I�pL�����h��5��@?A�֋��xx�І�s���J������+!�o�t�K`+١ӣ�^t:�%$�3����^��z��Nwy3|:f�\Y�2�Yh�y2a�f؁�y���-Y��VJ��J�-����X}���EN]�g�[�7��K�>R������� ��Run��m�E�+�uN���7�	�24�zM�{Jڅ�<s�0Ev�-�V(G�4�t��`���n7K��HN=8^�S�ZE*����"��̕��}��N�O�A+B:֌nC�/�A	��������h_�Bgcц�E-͙�hkG*#/Ln�t=(��Q//:PnTN��S4���$Y��L1���y�.�0�_���X
ʞ��H�/��'�����v=�H���p|q�GP��jD��Z=��Ym;t���`~;��qH��z�ߗ-!?�Z1�0bS��2�J��v��9��>�P~�#�0�6�&�#��4jav��Yg�!k�7���$�t�Zy����羫��t�0!���M?�7���*��h����A����L|-�3&)�z���!Ǹ���֮�fC��AA�^A!,Y<В�"�R[h�6�M�� ���{�$�9cCy�f�߈�<x`ad�ꏞ���>f}e�;9��0�e<2�~w���K�>�V��L0�dC{u%�4���FU:2/����S��-�-*�i�]��<�u��[J���#Lj���aX���9q�(�
���`|�P�����ށ�ε�J���(I�e��Vg�ԞS9�x>�h�L�,3�u�|.�'�-'�vE�Á��<\uCU��<���%E8�4։��k9V4�,�3�.C��&�����Bڝ�S}���}�f���V�w/_^����q|��~�����Vm�o����8�Dp�z�o�x�:4u=umبb�߮Wq�� Uf#&�a9o۶�/��^JD�*;�ӽ���̈́ݰ�4�;�z�g��@@�;��"z�w�HK�@9����Ex�~9f��R.b�ژ'������ca����f���u�wN�BF����J|�J�w��M�+��#�Bh��/�4_��mESa�G� �_RT��T�"��&�e��|���F�I�����N����902S���[ƣ\��x� 2*��\�|�	/���n,�lkʰ;�S��e!=�m+��e떚��%���N�1�]����2@m��P����Ҩu�Y*�h����e^\��vL���r�b�Z�CA��j����{�/��7��4}Yar� GzASg�c3��^�Ϣ����Iq���
M����]�~90�4K<�yT�����4��nz���d��I��	���\���I�uӘ�߁���g��	3O\^�g֪�T��RB
�c:�A���`+`~��.�WɆ>���=pO�Z��k�gM�)0۸T
�WB�Hx��ݗ�1���M��AH˰!�xM{���]|o�*��Te��O����IlG�R��f	�l���)`̞k������KxY��SI���6��@~M��e��� �	�z㩘������7�_��1U��g ���8P�{IӽQh��.��%W=����A's�d`��_^�$�ἴ1��*�@�>Ogj��l��� ��yx�r�E5�z��3�����3.����������l�R�������4�m�n�{��tw�R��hb�i)�1-3/���(�H��λ��q�������U=�m���p�s�3���f;+[�_��qH��� n��q�:���e@��쎺 )GUj�՗tq���%>H��f9H�R��:7�����̌tNT�=�9���aer�IϿ�����Y>� �����o��@�4i.8/<�/�N%|�4����k�*�d!��[���\��d�V�>��~_MZ�i��{K�=��;9CD]�V]��M�|��N���,��`��9�\��rF��lk��
��BL��� #o����nW2D#v���#��Lm���Qf�ќt��qP��X��K\kQ� ��f�h�g8�|�@�]�W���v�q���|r�"��f烒
43�JGZ��َA�>�J��N�>oqWih�+s��Q���`uY��xg�(љE�� ��3l*f�9j�=G�J�w����66Yij�a�t���zs�dcl��;%���d��c':�G"�M��:(y�������͍/~�x�8f[SI@�[�8��دr��3O��Κ<0T��,�Gq7�)=�;�  ܩ`�V�X3��(իK
%��0f��2ᬾS�oP��>��^ܑ�U4,�	-ዼ�-��r�u]����b[[G/��6�b�E��MA�K$m�O؄�lc��)	�?J���X皀�BAO��E��o��;����b�Ө(ic�hW�3��u�_��4������<����w�Za�9C�}<��1COo��W�uZ�C_������cF?=�Z;OˤMwH`���EL1ui�"|Q M�Nк�Υr�i����S�C�A� 	�{o3�ݺ��bl����E�F��p~��h+��=���0��i&,�S37���X��mEN0���M:�b2�28@���� �չ���M!9�7��ϕ.W�;��#,-��et� ������h��\��يv��@H3�������ϱ�f.2��"3����)e�[W��D�H�`�<�e0���JDE^��`9ϱ�Jt$#%� �~��q��`�6&���=�k�V&G�tf�b� -�o�[Y@[�_^�}l�C�
i�-��}���X��g���gm�.�K m��l��]#k�W�.@�A�|�N������`��s>c��N�>�G��oF����@�� ��3٢�R�&E
b#?�[��[����� h,��f5G���� �9��y����9��b�SG���B�۸J1��Ui'�(׼=�ӥpn���r�Μ{M�y ����1��}�����4**bx8�*����%`��~hb`�Xz�� >^C��� ?����n^��@��~ ��ϭ���|�ix�~�����є�L�+Bjxa�b`ty�I�����萺�)yp5͋�����Z��̱k����_��}�T�'���5�3,ɤ���/I<c��|4��V�ݿ�ecK[ӈ����@�Te���L)�$)Zz;��D�:r���u)�ݾD�1�2)���}+��Dɴ e��{Q��e_�|m�̦|Nx8�U�r�B�5'E���˵��뎣0ѐ�o�Ѧ�#��p��m�vG���I���?MF� k��~��0���\s��4� �:"�-��i00� ������ ��vb^�����������(qW@�O�!��쪁v��m9\��S�]��e����0j�.�\ߤ�����֕� �zp</+�������$1�`���q�ps����+o��Z��߀	�c��@9#'c�8���i\ۮ 捾+$�P�-�Y��p~�E
�ݮ��mE�}�Z���.���J�ɀ�{IY���G&'������>{̕��@�{��P�Ց8����0[���0�C5��A�nd�Em����J�3ٞΧ�Hefui�)��K�˕� 򃛉�!���ݎ������88$��$P�������v�i(��$�r�(tE�d	�_��F�\����Phow.e)4�
���+����.����լ�2uvI�]F-' ]�����0��&�r�y'#������� E_��b����Ũ���� �� �ؠ[�����}�Ϙ�J�ĳ����]X���Į]%�@%=��w6�ץ�B~�Ěf6m�O�!�1��G"w�2���( �Q�6j�{���F�\ls|� K=�~f��T�s�;��27�(�uQm� ��l�]����}��q�@�h���\�$E�%�L�5G��)�&"��W���,l�5���pSz�(�252�@��]+�ny�!�Q��{֫�B�Xs��Ԗ�,��x[�x�hIk9�'0V��̬H�I[�&�I��.22g}
�ccL��M��l�/[a�0C�H��̎�}[W�����;-/��^�y��h�mM��$&�! #o�H���w��5�J����X_����!��ii�Lo4���¾<S���A��z:|�i�M3lz��49v�TL�J��{˝Q���?fS�b��Lإ��Q�h<���6�W��h�R<�+�%�\
ۉ�|5p�o����Ӈ7n���NsԨ6?؅z3N�J���<0�+���wVC����҇�©u%9Qs8׿�!I@�twl����5�Ԛ@����6���?��x�Ixcɓ)��n�Ɂ�����@���3h%���(^,�VL������x�UHl��PBkBƑ��a�sb�OM�P�5H�8=ݩ|Ҹ��R1V��\�S��6�Y����hP-�tѢ9|���X��I���C
4��I⯗	y�莩,��$���ߪ�&s�7�=�!OL��ݠ�v�S�Y�ň�.�f)��EL��,N�3��u���gij�����+�ʎp��yd�QU8�+��=����<��H�f'���@��6ZdT�^t¾z9P_RH�[*\�+CA]��9�>����x\jfwy%p����eͣy�UYam>���r'L|����Կ�,�d��7��d� ��X�G��;����t�V`'�����i��ȉ�Rb㘬ѫwo��!��h�wmT����R�$�@�+�6�������MŅ�؁3x���/����6SA��;vu����F)�p�Hb<�r��0�O~�S�d�U���H����J����{3�TfZ�i�
(l�Bv^w��2m�yۏ���� :׊�h�����d��bYLgju��k�6֜����G�U��L;:�W�M��}�*��FMlP�4*��U��eD��Ao��^��Vڱ��?�&?����!�����i����̙^�rY7d1$u���h�J	T��@-0�jn)�۪;�����V	�s�s )^?|+�h���N���W�Q�ٻ`�v�H��N�`T^�����v�i.�ÓJ��E�"~`:L�0��:��n�@��a&6�p�s�u��ڠ7�j�a��[��bGٺ�9���� ܈8���E�e����q�k��{�B�o P}�׾QgEN=c�"\⡺(��(3�V�b=���[�|+�8{p�h���m���*m�N��0w��0�UL=��f�^ی�9����!�9/9��m�'�[�p��u@���{]w�Uo���9��8�}��1�r��K�?�z�N�0b)��B+�z�M~����3k�{�z���tg��gŅT���T����L��HX�]���Đ�NJ0�<��Ɣ6��j4�	�ȋS���?�^��[.�]�g���� \�P%XX���V�	6�E0`pP��`���#�j
�L��4���x�Z���lgB�,9[l��w�f#xN��`LI��s��9�ڽ��'�C�����1d��y�m)gXr���ǫ.�I1���-��.�=�	���4�-E���:�+�,�<�V��Kq^�-��|��)~���=>E��~��P�.������M]�$�qd��ӯ�O�!w�_����E�"z������,���L��ϣ"h��w�J��ï��D)�dJ����e��uo|[<v֛>��0J�#���k�?dC�T��%wB��C/G1i�=w��3�d�;[�p��I���U78D�]�[�,�t��k���*M������ Fgef���c�1'�^]�����u����7��;w�˹�� ���'����BOy�������p���	�%)�w2�<t�#g*6�+�h�?>{냯ϸ�1�m��f�i�@cë���E������0v�6(ɔ�l4>U:Q���{�H���|!%Ui�����ks���n��4�_�L��'-�����B�QO�eۼEA��*kk�/<���yϽ�
�P\�
fm�yϋSr+�e%�z�rJ!���u�O2��QUP����{+��5x�-]�����~�'h`�2E�5T>��HX���Jq��3Tc@f}�\R���6�̒��`�E���J�`�w żyvA��H�\(.��zF��S\{����� ���fx߷��G���%�x�+�V�D�v��MX�� !y�2�$j��rr�[ )��SR�����6�2g��vC���[����B�+��]��C�'��:�����;��S��7� E�x+�oP��R�ߎjw_�Tќ����8��K�x+;J�r���lv�}_��!t�
6l����3Q�@"�v�Q�@���U�E��{<vr�˒���`?��/���_�m��`Ñ�FG���OIh����D�_ ��gP����[�<�4׽���^�]Ҹ	�žbd�:G�^z�m-m�.���������Ƣ|����%#r�ZCPq�	�X�@��Ѡ�������K���1v.�����!p��S)@�^w�����H��O6x����J�V���70�l)�R�[����cP� ư�,��&n����>�,܆���3�:O>����G�W��.5���(ے �,r�v�
NX�a�QZE|q�W��?�.Zڇnl���l�O�\e��SSe7� /�zGb���[�8��8�a)��	 �A��/�*N^�]}��zOiw!�<�W����$�#��|��]ï���'d���s�dN�Q4�v Wj��*yMM'<5\�6a� E�Gq���0���Ygl��<�©w�Z�°,�\.�BQ&������S�����5���7�/5h"��S�drO�=������7Վ=�z?yc�p,D�_õ~%�H�)�ͺ��U���B3� ��ƻ�^�P���{�P�Z����Rg}c��j"^�Op[%M-��L�v⮻�^+j�7.S�9Q�����}��ݏ�څĦ�.��@�e��g������I��VHг���Ȋ��rk����.�ԟ��b�jDN�ښ�3���X�?�&w���g�Db�Q��Lt�ju�2F������M���"����Ӛٻ	��@v�Al�2�"���7�+�*0Nq�=��-�f2�b�`���ޜ6H����
���'��]�u��O����\t��?YE!c.E�lIH�OM�{��X��Q!���%�p���l���ZS
���ۀF�9�WtlS̴�^��lL%)gp�kU����u���(�x���fYE��k��T�����l�A��r"���*~�'Csz}�)�<48g�ĥ�E!��g��E��e�����f�<�6�Vgژ�L��I���c�K�:W�YV���n�uo�������.���i,]�'��	�>ϥ����&��>0���"�b+Pp9=wt�F�`����-�k*��wQ��S+"sW?��ɥ���V�'yAqƊI��lM�,2���l����h�c���ʧ��p)�Ť��~��~�d��w`����)Ƴ������)~���5N?h6����o�Z=�a�WY��k����,��5�˰��ɑ�����gI=�vB];��<EARb��ō`��1�٭��
Y猨�-U�D��>��̜m� �M��ܾ<�r��J�����Bv4"��� �$���
a_A�̦̳S�L���HA��k�f�%�h���yn�T���G����^�chc��I0��SLc��6	��i�wz=�Zơ#��&-9JR��:@�V;��S$�?�0J1�0՞�u�i��WO�߇�E����hKjд�&w��e%Bf}����j�Sm[oyl#V�{�	�#�Q�;}��VC����I���<i	T�E%e��f[�����傑�J��(�U���)|ޘ
��{ "���n\����[�����!+a�b�:����RH2ä��7�]�� ��DX�V�&��Ɣ�:��e2�9���!��ȿ2��&y)v`D?�4�Z*��\ccm��B^@��x��!0�����я1BڌX���Ff�<Z�CcQ���gu�沬	���\uB������p�칑�����)�W�^�����W
�i�VO���U�ec�ٝI=��C��X��1Қ�G���J'a1����ŵ��A<~�$<L�ř��r�c����_�����t��QR�S֋���2-踹gaI�EH��&d�����l+���	߮���a��x���ͅ�๿�~:�G��_G�Ck.ZA_H�~��@��x��G�QY�Q<:L��΢�<�)�~�T�!ݼTu���:i�3���R�@�6�@�k)融�iX���ik���V0��=?,5в2\��Êc�הbV�H�=���zb�ϭm�A�奢��b��������8g�Ҹ�����)`=ᔢ&�Y��EM�w�6W�`i#�K��<�l��|�0.�����1>�	���J"��kTs��[p}�Z��T�B>n��}�.A�M�E��?!�4�)�H�^pߠ��d�N�H���H6�VM���#�gP����.E���ڝ�]ħ>E�u@�m��pX7D !n��3S�Z\#Ӹ+" *L�����s��\/VR��x� ��"�R�C����C%7@������gt��ʜ��Y�/�͟�%�����:I������ǀK#��&$�]����"�m{/Oas���Q��7!�l~�lKYԁ�_oOތt-�&dY�!و���L�^��8q6�Ǔ�+�/�1�V�FF$�������y^����:���E˚�[@k��� ��7�1 �r<�0�jl��AYqr���f�L�sP���UJɋ�R�)0G%I����3+�f0��� ִPI,2?x���O7�Ht�"ĬgQw�ND�n̖�O���1�X`���l���y�d�Im�)K3Ӷ�
1C����Ff�@Z���v����
Xyh��C5"S-���d����7�p�h�릵��C���Ӷ��`�u�B�r5-�Xͥ7��xN,1�Aӛk������o�5��j
w�E��nW�|f�:�$��%�C D+gF�ӻ�S�,�3��B��?0 ,����.�as�چ-���
9������.��d.�`�yBb�,����䳌B��z������Ŋ���FF�?��5&�N�Z�Ī;��EC���p&� !���D��IGM0��u�[�h!�q\��̀�T���[
�Y��W�܏ XZZzK'e~�jW���E��5i��j�Y����@
()&D���G�E����iӛ����BI���r@�j?KKԷ�k�Rz@vC�-�Ƶ�	��ǧk��Voy� �����y�� &8I"�qk�ύ�����z�q1!Lo�l[��l�'jƚԘJV|5�*ԙ�ؽ�䆱K��4��q3Ԑ�G�Ǳ��f�x�����F;�E��t�6.�u_PS܋rwe�c��rq�-���¼�����ߥ��:��&S��e���%ʴmt��X)6^�7�5q���S*�BW`��;2;7������ ��K���I�9����<��YKZM6�N(�$�l��-����G�d�Hvu��+a���(�G&u�9��^,B2��i�rM�JЅ_͋T�����5%K��D�����NH��{)DN<JY�J��� �]���$�Ku��vsa� �m���J��|Mdw��'v���u���iW����4�g������䞂�����l)݈k�I��pcC�6���&T�k�hWEV/�,�4���Ո(�Mm���~���\z�L�i_*%[�:�!����a�pg)�y/`�@���	�8~�&0�QiR�G�_$F-�xIFh2�����/��nY�x�Y'ֆe�_��������h���k�=�Ƒ���\����;���N�Bo`m��D�F���	<t�ݚ�5U�]${��m����kl0v;��v�O͸MΩ	�j��D���&�O����!�S�l��Y�Ԗ�q|�%���˄��VAw�KY<f2=9z�~n����z	!�"l����m�QQ��ޠ�+4ù.���_�L�Gٯ;�E4�;�`�9''A�"�$ݿ%[Ppi�QXx�s�U��	+˜S�GBr⺚��;��-Z�m��֊A�}���`���'���a��~]q6���Y�VRzI�b�&L�#g�K�� ��u˵�C�d�Ǥ?�ZK�mR�H7��Z\M��%�śQ?�H*�yJ�a��"&!"�g,�Z�ӓz2�g�������&3���GN���n�7�.�P��v%{�A���/u�kU���y9�� 76}>x�����	��]��v�ô�m�Ȇ,�ֶ5��6����fu����Gt�\ϋN%�B��b���{�j��ݼ_(,�)6����]�&��bp�},߅�N���#ؐ��������c����qQ+8���a��PŃ�s��؋��1ѩܤ,�Ȗ?A��#z����\�
�.[sg�Buv�������D˿},����c�5��f��1{M�0Y]`X�X1ݪ��*Ks�Bڧ�UD�/<�miHh#��*�T",��fjz��(4�70�|���TE�D�����m��h�}����F�,FcE%����F�/r� �e�Nd�h��0ę6�J���L�7���}��=�Cs*��,�C�F���G<��m�xh��%CE�|J`C�Uu���{�M���Q�m$?H������RSMp:--�3�b�¹A=7O}���'����������u��.
�,
]͵�'�̿{
�l_Q�b���f<TZ��4�y�]�F&���Ĵ�<eAQ��p�S2����r�k��q3�*��3[t���93ٗܖaxu}�y�$��>�c�y��ٍm��c(�^rxXC�ޛv�ʛP��k�`�0㚑�M(�Ƌ�����+�"�೵ZT^a8�쬏3l�x����aYb�*�����=���FD���"sB]��z��p�|�L+c���W�<��@GyJ�ڎe������OU��&QNƤ�Z>*��'����lp��ڃ�ԫ�(�LN2�g����L����_u���/������V[tbs-�����8tS&���&ͼ!����s���P�Q�i����������sǏZ�N����mep������m��͙,�K��﹪��($�2���^�}�ìbc����ɨ��\���G�e.�b�M��FZ�Sf�r������>��S�0ӯ";��M�v��ڀ#���#��;A)�/��6�]'�D����!�Qwv�����mYzn+Gs̝�J�u�,,Kpj�I��^9:(�[��`pin���{֑�*�nIC�5	n��1m��O��U���B���i�Z���ք(���Ֆ8��Q�ַ�!M��jV5�0�ײ}뇧iuŠ$+Նb��=��g�P�v9�'s���^��{�W�{�
�#�#�:Y��-]X������Es��u�e����I��(/�86��D��$�cRo��a�B�a�����D��7��1bի�aꏧ;�O�dSPU����6��6�������u�j���j����8W17���}���և�:n�R�fTG�d
�t�w��d�åֳ���ܱ
eڭ�.���r^�7���}ϊ�vb�!O|g�'�hJmլ�0M��:��,�}��QB�_�'m;�[�<8y�{=9�L��_�<�^4�Z�u�2�K1^Ȭ|�e"n^1�ΠOA?�Ro����n�WnFL�]>�bU�1�Ǻu͋��U/KRh��u+���(��l:����o̘�_9�����˛H�O�6��3K�0�M�tOi��n�PzJ�XhޜҀ�[���g�۫��=5u����c'�2}�:���f�x�;�7#\���}�j����zV6��n��y7�|��ʽIί���j��I��3b��U��z�:I�&�jO,!S�p�Q���n��ξ}h�=�>:3�,]�,IRYRA��<�usч�wC6�
#�
����
�W�����vi�����I#�Y��w�_�g����G�U�.�ޘF3{Z�^����Hߨ' Sw'm���Ч:�z9v0��>��ѥ�$��
=K�X7B[G��g�+6팷�����fw����L[>��2?��l9�B�^�����_?�i���������O������4M���'h���ץ���ژ�����8�������o?����E.�sџ��\��?��u�qj�����yY���=���_�����ϫ�W?�~^���y�����ϫ�W?�~^���y����ݫ�g���#��!����2Ō"��XrBvL�R��������z7�a�M{�C'9;?qg����y���V@�$t��<Ӿ��W�����Ϣ��j�Vz�>	i��y�鸖Ք���_1?��'k"���xc�۫�c.���qC��"��lj\��foN��>�ܯ���g��?_����^:�"�p�+k��=^c|�]�}�(�-��/[[(�gԢE��|��MȀ>WϿ���ԓ��Z��{�T�U���_"o�@�<j�7*���3��";������+�]f�p'�����7��0Ȭ}Gv�/��>j�Ӹ��N�����h2A5�f(��Ɔ*M��싽��F��^\9{d���ǎ<�S��G��h�ʌ��G{��e��d���9�,t�E�恻D�ŉ�4�B��%H!��hK��/�A�5�ۑ���ص!<�Բ#uO]����tt�h�ڷ��O��/+�h�Z�D"�q�4�� (��X���4v
����.D���i6�:�3{����?�����������@�_S���^���x� �B�m!@�e��xt���:k�����{7g�)A~�ٳ���7	<z��q:�?O��n\�eǎ�+����{(T��ީ/|�x���6t/,W���2�-�.��?����C��,��b��]��---r�hn�����蹑�hw<�5� �NЦ��v�W���!���f�NP��~@Ӝ�@�d�-������4Fkg�Ǐ�w�	ٗ�欣C��y1���#B�_w�h���O-�s�����3���3��P<ǃ���SU�B��h^o�ױ����B�\0�+�x"z�2��˗�hz� �Wn�&!�ko�st�T�ϓ+6���_��иi�6@K4WJ������N�����ʀ��˖����K �6����u���
��˗v��n}�L.����V-��B���4c7$׳�	�S�$Mss���_h~�w9�(X~�J�
�wo_�^:���v5��׉9����~��I炔���0p��#ݣl@2n±\���]�9j�r� `��΁^����v�D^^^�8}m7�pH��(mY���e��������I�srr*�oC���=+z�`^��h>���N��ksw�<�<��0z1���9���o{Fgc��F��^������2wss�s����G�Nt�,���{�N��Jhؕ*��!�����֓�k���SGg�ę$��tws��=�+.*�z�Ҟ���ny��E�wWrfff�i(o�eO��g��~w�ݺkԇQ�P�&�?0��p��.�l����w���Ԏ� 剿����u�S .�=V�W\H@����야]����(�u��^8��f���w�%��C�'
�m܀ҾVt7�n;���f0�����py�n_��+ X��A���ce:���s0 ���O�7Q��-�O?�ض�7�<6,چ��L�]t�h���	qC�nn>C�}u�ޫ%|���Z*���ސ��ׇ���S�Q���>3�AF;(�A1Vc5��(����3�m.[�YG��J���=���0E�|�� ���n^|K�r]{A��Ƌ/��������-,��*�$���YK%�8ǲ��hS t,��R�Z�:x�eb�@N�x�h��1�P`���;2zg������_�j5{��U1#��G	ͼ셯@q�|E[���ŵ�.D��9�'i@Z\BV	ьf�_���.���HÞҥ�4|�G���3@y񽯢o�8���պk�:/r�1��k�c�Pn���4-������ U�\����\'�K���{:b�I2W�I�p����ݹ��
t�Z��"�!���.�:u�!�k��s{�S�\�L�q�7`�GN'��v� �����׼nFiM�%�u$d�Tb��;��{��� U3V\B��AB}�?%�
�;z����Tj0d�K��d�U�l9S�L�X*+��z�4����{*�K�
�!���ج���t�-^<��=4>;��0�R�6>�� `�Zϵ����Зhܕ��\k	L���s�S�bF�QpppG�c��^�����f�+g�K����xUcOU��q͢6�t�����斁�
� ��+GUx������s���+�!I5;{�) ��W���F+>?���)��b�E�����.�Ɏ�G3:j�_��ɪ*�h е��Ȫ�D> y�w#/������z�6�ubIXԣ=3���bdx1ۅ@��Q�x9$iה!�مSuuzR���}�h����P�J8~�� X�!^�K���~�����):LG�|�W�/�IY\8����@�[���忴U�?ީ@�{cq�ͨ��*���)�^�yv��[����0ὠT��wC��@����D�!r��M�Rs;�%"�7�#��:XZ�CszΞ�� ����>2���H롍4m��y�� ���(U^�@����{�W� f�������Rjg�q�ǽ�����&��&�L~����+x�T:!�ڹ���(���O���|�Dc���2ю����:r�Hi��f	9�+h�\��s�`�{ (��� K:�h��h=��]QW��?FFcfgeݦB�w�4��C<�s��o��?(߀�N�נ���u4u}���V۪��VPQ�PG�BZQ	(���� dD�Rdoٴ�+��(�� ��^��B
2�)�Y"���G��O�ͽ��9�s�}�����Ԏ�:s|'�u |0�+/��P�@���b�t
�!a�O֞H��+y���kB��*�H���y��CCC��}
��h�#��NC5'	?t'b�<q��Tx���UM���K����!��5�J�QBg��2b���߉l���4�	��K����d��=i�B�脄�{wQ����U^)�6��:?�~P^�~��KM�18a1l<-c��s��B�֢M��`�O08�4k4%����'{�҃��<�&Ҁ��$�G�E����Bm��0M�byP�}�s���چ��5����/�Y���$�j��A-�c�87>�yP��ƉT0�W�b��ZJv�K�zB8ʽE-�̂�$����j	0}8yqee��<�S^�ްu��ya�k�v�� ��t��,��~9���љ����|�;Z�=7�{%�\��lI:�cVou�K�r�NP�z�:}!�8@lM�P�ߏ~�����TȓC�sK���(~�ܢ���zU�6C(������8ޫH�*�(=���hɿ�h9<\gH���&������S|lG"��_����z�,�׏/�{�f�`�Do�G��3��sIr8gOI�����LR?�C�XqvZZZ���|XY��a&��1�_㿑��c�G|v�0����̷^��! ��b�6P�LD��p{q��p�j���p���]v66��(�7��E�A������JRD]�>j*`��Z|Y���ZA�����:�e� ,[q��l����˗/�f*�H�������]{���D�۷og*��C-��Dݘ�
4��,����շbB�������1~JT!G�4��Ign�~(UsI*\�Z��>��sn���z�~p'��O�)mo��:b�w�Yd9K�A�uY�
������i�/c�/��P�z�s$�r���k�Vj%+yi�qC=A�V� ӕ	�˩��_K�mS<�n����	]L��_���r����Y�w=��s�^Z�'.���(ԣ�l��q$"�Z�ɞ��s]tՋ؊Y��,XK,��~��]������8P�&��g�*\�{�KjU�˚�E>4� ����/ 
��٭?�eu��h���/�����_9A�b>-|�;�zӥ��Q�b�)m���]��k��L�ݺu+��n�}�&�t�9�j楫O�2P�|~��
ग़��{�z��(��fR@���Ʊ6 7���Q�s�����v,�b���ήH��Gm�Rh�gP3�%�Ɨ@ܿ��Xp��^*fE��)�g�b�Og,BQ*c�V�a]V�}�ZT��
௮|���{aQ�H�7
s�Q�=�kOӏ���Nī�B�$2�e$O�"�#�J$�5�ķ.�SKR�J]�IQ�:�+m���ŽHZg��^��sS�ǗJ�>���*�F����Y�? ����)S�:����&E�����Vdu�-��u��`��8��7��DD݉��EB�,
Th`�~JK����#&�k���C�c��IE�Y^�S�n�Yȿ��1���"�B��ɉ�٭���R�{\�PW׮�@m��h�B��2������g<@6t����p>QVշ�k�{Rs�1;!ٲ힕Up�cL�����>�X_�#����m=�O��,�L��y?�qh�D ����x�Ȣ���J4^7���$2�3��y�� ��.Sf�s�*�^Ut��T�|	�$� Ԓ�H��Pd�U��k{{@�Yi6 �%��]q�Q�c���R��ϝ(#e撰������	���������ڴ���1z�r���=U��dH���ێ�>�	s�@���!��-���3+Zِ$�a��bQ���i�ROR50�]]],}���ϻ����ފ[��W%:��M��u�]��f@�~]V��m��#��;��y���J���i���mE�#65}�WQZ���!�F�JD52p�������*}���M�H��h6 f�u�rnh�K��Q�T���Ce��R��/gK� ����Ku���s��}��(�Q�˵�"O�t�O(o�&��;��E�] /;��ٝ�%A]�V(Z���ǇN���é��l$0|,��pL��GD��Jzv�FE]����YV��i5^UUe�N&��-o,^�߮��������?���O?��s��ӻ��o�0������[��m�O�*RRd�I����t��x��1�o'>�sݟ���[��ݚ'����V�8��������g�V�6`��n����-��;o��pa�2P������Vp�|��%T]��'���28��n׮�ݐN�U_��b�Ӹr��v1�o��|�-�k��Я�>T>��tP���� p�}�.*&�&�g�1��{�Z͖��v���e�}Z��-�P�إxz�z��<��;]b^�$'�^����l�AN��a\yx����߃�2;��{���A�Y�/.�2����cc��t�R˨��\�6��]�+�cnn��ś�`8T�l�|]wA(oԧM�6�����Y>���	P�(��#9��rVH.�5�a)+�u_������J�]-��]��Nŉ-�
��{��?�)ͦ����	W ���rC�E�Ы�x8�η���{��c�������m�]�֝���K�}�_\Т��{w�X���]@ለ�X'Eka��JVJ��#n����M݆��ޜ�*_􏀳#\�=�����7��,g���(����%�ٶv!�qOd��H��R5f�ϙ��Ǆu�0�z�)~T_@a�b�/�o����Y-3P,�u0g�΃ؔ�o��U���p�]�*ځ+�^��W�돤%'w�Zu�*��9�ϖ�%�m�=Au�y?ڐt������'W��Y��y��mQ�0�It\`GxǪCԄ5i��K�� ��G^��.�o"�n�Q�?9[UU;RkLYj��/�sK#[DmՂϖ���3s�;Kq�o���E�R��=��^�b[ب`�DTq����ڪjk�<��FUr�!\��#
dܳ�m� ����;���?O�6-4�����Sf�]�����T�s�Vm��^m���߼�߄4�`�B�q���w'���V���9P��!� �`>��M

;�(2x��`�b�'�Q+��>�АPᩖUɕ7��Hg�����F�����dCh�]K$�~H��c#�K�w4ݥF��7����'q�+��ii!����.P��}���;-xi���>}�t�i�x��8u�t��ԙE+Y�Z��EK�A�{��Q�gA����0{J�;���e��j�(h1�&�P��}�^�LcC�.�����	��G�v�F�Z�V;�Z�.�*��ҷ��-��Q�]�ioP���E^�cLvgSq�F��H�@���?��3��Ө���6��c�t���T�G�G��s�[�&�G8�zb	Lܠj�8��ꔀ��#%ȸ�6���º�11y����QN(x��ݼ�,P���2�5�b^�!��QG���\Ȳۉs�8+�y��O��m�7;oN���N>څ�?l��d^lb��\�GΉ�6�fbj:�B0^�t���Zr�)��z��X!Wp�nÕ+V��w�T�p	WUF����_�h�pP�㓑g������H~N]'�xT__�R�Ȼ����c�������Zń�ꪠ�"��8���`͖��k.��.�S�U���4�����75�<XJ0��ڂ��U���M��Q����u�{��$��$��q���*`hv]!@�&��'�}J�I6����!R�=��t��>>}+�=5D��6.�јӧO��u*T?�l��+����G��dge�>����T_�2�,H��ī�;��=��X�8@��@��n7h�M�f�vJTQhɯ�(����(5�)�N�x�g�N���]��8Mfˡ"z�k�|�pa6�G���ݶ5Q۬VZ��7)S#��ͳ��%�!�9���~��r���^�?�ª�F%�,Q��� ����HZ{���]�*�l�`�-��J4�f��y��0�j�L��˓D�hY��/�A��M����2��I�|߆Ϙ�B0�@�@eʡ�*�`32�T�uÖ_��9�#z@V��+��c��f�N*��fk�h�7rE^�yiMY���%{����vd׭����.�����/���5��>��!����27���ťK�"���è��S��ۘ=GP4���������WH��R�{2L����]��՘�gP�́c�ȕ��e�
�Tg�֨��7t63�(��{�����"by�W�7Ko1=L�hBcE8�B���WdT��6��f���Bmbх @	���|<۰�ɢ�`}��d yGҍ�+di�/��x������66A~��BL"�C9Q]�Eݾ���[�k�/Š�0�X�^�'�S5[��W06 �4�h�i�M�/��4�E
�F0W۲X"�j��"0+����q\�Q��"5��N�s�&��s��7�̝��r!��J6�6����:f9�.�T(�+�]�G�Q$�<0�kkk7e�]ܑ)w���I���eCǉ����S�t��%VU��վ[�]�o;��~MM�ac�@h���O�~?�$Q�*3Y��� T��/�If�ަ��Sk��& ?Nx[
UF�kJ1�t[Y�b4�ڏlɴ�����ɗ*��_II�g��k�Y�98.�`T���y�d�.Z�W��]!�y1=��{�<Nx�����eBN7 �|p���9/fϞmp�+d':�o�ْyQg�, d#L_ɼ�-�ȶ�F�_����WZ�b���M��w��6|��!��s�ہJ�Q7g ��Ǆ�����'OYʭ�L�	�Q�<a"�-I ��)[b������}�)zO�$���-�h�T�_�N{n(n*ޅq���@���Ċ�s	���"�;1�Gۚ&�p�Q{ ��:놀��LAM�~8 ���+���mJ��D>�\!_�?2\�Y�,�����:�0ݐ�q��1k�GƒH�����A�~�/���g�Y^����m1	U��T|1��r�d�y1{��h[�Y�P���ʷb���Ԣ&~�%���"��)�v�u%m�B�kC��ac3�S�e�3�g����t5�,'�r�$e����[�x�����4)�S���ԏ��dԈL�kz���HB�9fT�)[�lY}���=ᠼb9���k<u[{^^Z�62�5��ko��Ŭxf;�q�3���1F����TJ� =V�-�<�%M'���׽�=}\�_�H�n��������M9��g,JA��=I�⢒c�9ׯ��"�}N+��k�(s���E�ˆ.u���>����:n�q��ER�gk�+�'�@����8�c����Y�ui�� @������NTTT���VJ-p!��{�B7c��*�OeK�D8�o�fއH�P»>i��U$��N]$2��)�ϴwδ6\�@��/S�9���XY�����n��@!�ϻw?3�2����]뷳	g��%'��t�	�l���e�F�����6��b�����������:v�P���*$���455.p�YAH��YJ܋v�O/�^F��  *�D��W$&o�Ci�>W������G��� g��+�b�g�sR�q�+�;��d?rK8�#̑�6>�s��Դ?  ����)
͒z���
B���
���ԥ��b�$�}�����8����:�rEe����+o�@K��w�<e�1��w��F�H�[K]'���iklū�A�w�?�3��J�4�n��8�ɖ����V��mx�`�/uo�뱿<n`f{{{y����S��366�$�,c>%d����<�y�o:�I��̺N�e�چEdV���|u1K�{�33(�5\c^�%���S�\�[�;�nζ݆���U��b�^�� e*���V|vw����l1g}���E���v�eD�/(�f<�t����,��(�����g�����4�HkM(=�>Ė�^`���MU�dE)M�M�d'�)�Dlʮs�Ri?�*�o�<e��O��xrMnG��n���A���ӡ��ָ�M*`]w����u<o,�?e2#(H�ڿ��G�w"v%U>���ƶ�:O��5��΃�$Pt�1���q���$<lg2=ȆnRe������G+�C�
�%�d�B������6�`w��6+�$�5@�,!%�	��|�����dTw����<�L�P�������K���ҒK� �>�P%C�P�N���x���
K��7� 99��M�T�"�@�d�㤚�������,�ʎD�.u�UP��pߒ�zѬ2�ۙ��^�oN�3�r 磷nݚ��t�.��ؘ=vGTq|,d�<�_u�;cd[?�� YJ���7N����з�o�N��dk�ק��8l(9�S�Ʉb���n�0v%''����X�W��ُSy �Ѿ�ϋTZ��܇���q���6��u�,-����D��A�tU�o~�K���1a(\L:���*��n��Q��Aʫ:�3�����ġ���M��=�_+��B
�C6��X��V��J}��X�D�1����m�.��hZ&B�T��O����STY�d���G(o�� Ld}@{��n/�g��Qv����[˄]x'�{=�������Z��å��/����^�UdJҸ�����J���M�LQ����؍��ח������ �l(/�q|=�F0J���Nu�޽��j�$ֳLj%D�M��Q���c]{��h|/�'���Y�`!�����)�<����.��+1�ʰ�,�sf�@@a���g+r�Y��p����;�2�0����ƊɨĆ���	h`����D7r����B]}V5F��܂���x��̻p3j3����=
���Ҋ�)��S�>_���x�� ������7S�.]:@rA�*��^����ƴ���Tuuu�Ν;s����)Uk��l�A����0̀(5}h84���^��bɻj�d��u���DEiʧF��"��#�u�B�p0����,��p�c)p9��N~�zuvH��U^�iܭ�_��2(��<y�V��*u��{s.[�N�k����۷�$>/Po��m��
nE��G
��ћ�R5<�!��yͿN��1߼�;�sY��z$�o{F9X�up��J��^P����[,q�9�Q/}C��F$��U�.ģ"(�V�)oޣ����: ��ǅ�$��Bܷ煬���Z
3��U4�®\��x�&�]�jYG$|}��R�d<� CO�z�+�KP�BTyUT1͌�*��}�63�N�t�[(耱��s^I'5�=Æ��E���;�G�U!r���}�Cy| 	�Rj뷷Aq��o+jKp7�n����#G�MO��W�rr���yw>��g7��!G]��.hJkŶ_��e"NTu�KV302v��K7�8L`�M�r#���}�U�����Dj��[���p}��n�%[���Ե����tf�嘨� �u�T�d��T�
:���Kz�ަ�%)@=IH�e֥��m�+$����C��� fF&�\U��]���D��������^�wQ8MNWҏ
�����
�#�j����US�a�5����5�+���7�"Bh��>,!�@Ԥ �x�=��F����Y-|l�I����l�|^y�eQI"-�п_�Zm굛찗z,�A}}���ׯ�y!�ø�/�)yi��"�Z��ϰOJN�������R�,Wp�nWM�B+�'�`�߻E�i�/_�����7S�}���������?���L䋠l.��xN�P���&L�*�i�kթ�jX>�� ��?��|����q�0sQ���)��="[�[&?v12�]>{���6e㮹�ڰ�-ܰ,N����]��5���{{��΁��(�3�ȑN!{�����n�oaT!����Rp�l��ۦ��wf5�S!�NK�-��Z�|����m�ի��ғ���k��Ny��p������h��
^��l��Ч��8����*O�����-����:o<�L������W����v9ٔ��qz]�[��k?�	��+���P�� an(F�|�M��ꗓ����@L��Bסg5�Џ�Q����U��q��CNQgΘ6AY�h�Jw}no�f�|��#P����h�Mr��9���---�X-5|�K�����,0�Q�IgC&�}CI:��^O�����������x`�*��w,����kQ���+����o���;R��tr�=�$0}�
8�?��4���"�PKWB�{�T��$���� ���t�Jcb�V�C7����Z��ͨ�ZNkO8�	�ޘb�_�)ڽ�Ly�Q
vQ{��բ�&���C�4�[��ǅߣ��zq]����(8�Tqϕo�0Νp�t��������7�%Ӭ�|��:���IϦ����z�yP��yGv]�ɻQ��V�,�5������z���~���_�����}��m��H�%����:C8��z/_8\��t
(l<��)͡pR�RB�Ƽb�k^���6a;�g"�1�SL�]���X��L{��~�e%L6�T�o�E!_�G�I6���@�.P!oF��%<���i�7�CX�A���e����=T����
�j1�Ğ��W���������_p��Ř�;44T>�ب$�.�z�C���N����N�t���%ʽ��XQ��F�/ch���F���bz�U��yp���#����?����m�Z�Z^#V8߽Y]Scx��a[(^�ٓ��u���M*�tom+++5�F��S�5��o�S�^A�bh4�[��}�a����I߯k�>������Ǐ�ƻ�&d[��m9������%�	����d7�&'�Ȝ��E5O\�K�?c�w�xDl�'����o��k��%����.��9];>=��z�jӓ�x;|<���>n��Q���w�6;�KᗟL_�D���������Տ?���b����MI�V��}��g�4prCo���~zqq\y�]�>^�q�~���P&u��yς��֮'W��Hk=�S�c��Q�hr"/-ʂߠ�v��`(�5=%5:�{o���?d�ip����+:��а]�
=��]M9۹�d�(�� ^6��׮]�~:��o;���1&�b^!��W�A�Z6��kM2\�G�5[ʄ�{�V���5u�c�i�'�ne5��'^�� ��"�8Ա\p	uwC��V���Nߑo�=��b�X������	�B�&������q{ł��:j���*�3U-���7�ݖҗ�lM�[�r��8jkR����$.y����)�-�5 ��E͠.>07��dw5O|��%�Kq^!cP�<ǒ@����h�J��������*b���\�꾑�;HS���K��0��K6F��Bq� ��{��������P5>�r�A�]U2���?bl�.�b������%�J2H��=8&�Fo�����#��o~q����PwZ$�����v�q�B��o��+2��{,�IULy'˵a��)-w?!ݗ�&(��b]g�r�h���COf7��u�B9whSr�K��&
�āG�|��s8���'$�W�M���6�� ~^1�Q<f]i�w�P\x=V���#Vb�W��wdKf-���vttXI4��젶���U?4�<�p���B�Ԡ5�2UHiQX,��U^;eHw?)
)I���ZDf�]�6]�L�3=amL"X��n��Sb�L�W(�f6ct�R[V?	��	�:ګъl*J�toNx�F���]��鳐�b~���"�C���1:��הK��-^Ê��9�lb�.`63 ޙh�fwZ>����Q��2����|�&r ���fw]z���PC7��e��%�*�aR�����K0��PR�l������c��S�4��+$t�i��{�����ii�XܻE���\�;��V:��w��8ө&-�e3{Ɖ>�E���&𡜥���P�JĽO�=�q�˵�'U&G9���lw���óٮX۫���ϗ��
F��1�!�h˃H�Ȓ��\ID\	��/c�V�^�L�6[.є	V�!>anT[`����
[�*�sTvi��^د8��Q��q�#��g�T�=<���ᙟ�J��i�s�=��.fff���`B�Q��h�	��-̞��l�᫾�Ř�Ը̀	O!Z.QѢbg��Rg�,N�K��eq	��ϱ��U��~������v.��=���B��#�"E�̳����z�~'��$�1���K��JDi��W_�Ut��!KXխ���s���N_U��t�ҹ�ր�Y6��w�
.���mO��ɸ�!��kI�R�M{��P#�G
�H?�	��~�#a�&�W[�,lk�]3�Z��8�Dcj���BDQ�� MA��g�G�!��r��!u.ٝN1�ɥ�EQ�H�ݻ�������e5ڣ����g�N.�5�(����\�5���Ib34Jڵ���Sؕ�5}�P���م�d����Q'/h�s.+/O�ыS}!��R��j�����Mv;���m>q苢�y�a�ڏR�;����*�P��Z�w@*H�e��`�u���� ��Ѱ�7R���z�I��t��o$�.��r��C����v����Q��l��x���cǎ%��IJ`��1�CqS�u|��9uLv43?�w���x|��wX��D8���E���ܾm۶�h� 2�4D��S"��)�"�K����6�����x>)z�U��ʽt�1k�DԞ��ڳ�7}��sa䅸)ϯ�1�AP@=�
���Ak^=����Zo{*��G�leU�t8OQ�p����:��	���zf��N\�:��;���������ٓ^�A����r0T�n��T��C�^�0��Spir���%{5[\[�7<� o0�
ތ�5���R�־K��e��k��f����ɩ����+L�+Z����|����aެXc_���Ǵ�v�{�(�?���&'���kW���V�_��[���*���)��H�G�J�=/���	J���F�9,�1�[�nL��k�-�my!���ՖS;��	5~J�<ByP��L(̦8S�#�0���-����b��5����K�M�������Rw��5��Nÿŉ";���8h�3��*�+��fW꤀r��IPU\�r�{R��Rp-���ݚ�+��6*��<�%��7}�D*��G����X�0�KV�Ă ;�hCV܁�+��!,p�UU>�%op�^}u�� E�@z7a�Ժ��{\y$���>�ە����C�#G�*SRR"�Ʌ����n!�篢?���KC�_�]��ܨd�sNԻ��$:����+{�t%�{ʢN�3u�Ļ|���*N��\y�֘������K�y�fS;����`�~�w��З�x�ak���l	)|�=(�}x��yL�M��Y�I5
=���{孧�sv�ᆊQ� �����(>�����(�_�jD�!���52��S�u|/=�U��v�}�Z;������\�:ȥcg�V��� �Δ�%_�\������� �i���Ww�ګ3�5��ț��	Р2�����{����:YT�(�_���J	o"2��íڑ]l)
W�za{� :�PHΠ���s�5/���5���0���đ˩�cf�:��&�٭��U,*G*> �r}���P��CV̠QP0o����T�r'7��2�N!c�N(��._^�P�B�{���T�����L+/cם�Y�L��������Q�;G���F�9�"���L}����u��?M��^�	p�����M���G�G�$xpE�4ژ��0p��o���M����,wq��
�����ׯ_�K/~����\��
�U�&��&�cؒ�5���G���YM*u�}�U_*��K�����,D�#����4�ݱT�>��e�O�am�3�E�6ox襔;a�os"7�;�7�%�;���i���?`K�l(�c����z�t-�!��a���	ԌQ��m}�@�����A[j���E�l�����a������d���w4��h�_-�F/��]0[RC�U>E�{�߉���wL	/j��rK�޳�|r�Co���"�=o{�j�ʙ.��+��(\��݁6��.��%�R5G�($��;4��=_nrr#�f1���c��ΧJ:]L��cTMA^�p�p���9K�=.����S��4�J�l�]�v����+��wSݸ����Z��r_�9��<\���ˬ:EvH،57/Ѻ ۬�~��	�"%�-]�rd;Ⳕ^t�m8�4��9���G�}ZK���N��ZY�=%ō�9l�g�����>��J��S�4E���Sܔ1��|l��=>����0�*>?`иL�FH���t����c��*Z����P�Ol�̥���K��չ����n��V\y�&������̣��]oo����K�0kr��?<e>��YxM���dx+�CX�$�`TԻ��Jrp=�� U���n�P�X�x�l�0��\`b��U�D�#���ό�A.�ߌe0\X�Zy1ќ)��0��Q$L���w�$����OY��y�T��+ߎ��L.�hgʹ1_ߵ�[O�U	{��I��2y�}¢��v5["W���
��"���_��aDp彚-K�x�m�S�x���J%ͮ@�����%�r�u�6�^�K�u���!w���dC�P~U�����Iz�H��<f�qa�l3���\�Rzѹ���}�����-5[V���g�I�<Z�����؄���y��L��B�HW9�F��ֈ�6�*+f�;eq��oUEE�L⚟ӳm���z9Ӄ��D�����5�~z��5΍�u��)U[�R��
�C|L/����{<���PK>ڈ��m����֣n�Ѻ �\\k�������X=���CU߷#����@�@F��#�4Bx�az9p0���,_����������)�E�e�R��!C�!t��Ԡb��v�7�i�@F��"22�JN��v��/
�_(�����w9ò�/����ɬ������Ya�W�i��K�Z<��5a.SJGf�w^%�3a�;v	����`P�.cK��q_���%�8�ig�+�u�R�+�(26Y�%N��O�c�>��lieG����$F%K�v�԰߹s'�(8Z�NLW��)�g�� ���Y� �W~u��*��w{ ���PP����Ӈ����3>���r�l�UX���f����/����|M��Wrr�v�x��w'-����q���?ƒ���b��C�?7�t�W�B?��Ç��>���X	�3��wym�{�ҟG�܋��r.P� 2��〢'��'zBQ^�[Cq��,V�����^,�3�cH��Y�~_�z	���#�H!��&�H�Z�|l3:}�����U��Qq�>�+R�%0��V�x�O�(�~��*i@,���zy��"���%�X8�������h��\ya�]`�y%�k�lP�-�͑��:���i1��\g@�|C[�ʣNߦ�2eǄ�Dz�F�]vv�7�K/�p������a�"lQ�,�c�l�_�}�ї߀ĉ���Q(���j��]��xs�7?�5�
��]8��)}-�кn��Z���q��T�H� ��vL5���T��ܣ%s�OԽ�،W�O�˹\�ސ\�~O����9���y���o��F�p�pG�<�'��~l�y�EQ|S,<�}LOV��>|�+�E�F|�/�އs}69 ��C(܍��.
�����O �he5��nJ�̵	C�D)ަ�I�/`f�t?��w�M3q���Fe�kh0G�'�/�{�:�xM�W�o�K���H���,ta�?>H��&�|beU���8�u��g�S�
�s2������*�	T�G�-��D�)�X�x���|�Vԃ��+J������I���$X��;�
P�W+M��~�0ѹ��%�i<��u�]��e�'v͜�ξ����6���hk���~ژ=�`є�W�4t�@����������Ŭq7���C+V� E����q]�S�vO��W��IT���(���`�M���a¿���1���Ht��>R\�B�&�jP%R�b#^=��m��)Ӷ��qG�裱����Y��j�j��%�;K��k.��
���+�%d�d2��U-�@���	��f��,���j�����c��}Fs�q���>3���1����9�1M�V�+[Ҵ����*��
��Ԡ��7�^�!p�XX�&ܣ��Ɇ�{HE�}�kX5~Ёf�R&�sX��Q$��U�UP�� ]N��1��''����r���]��j��jN��
�����\v
�~�����n�
��(}��p#�P9rs��zcQ�>�JgL����E� ^����ü����� ����}�~D����v�l�|�Ԯ�v�'���N�;�Bx��ǫ2�����4��ܦ��T��&��dac9�}m�K�{�F+�`w�g�"L��w-z9DD��� ��ki��þ`�#m0I`�I��|�q���*G��LKk� �;=�fl��ڞ�Y��E�/h?�q��$9��S��K����hqW�v���l�/�|2�ri��6~�$����5��IK�*K�e\�������璓#�J�ٜ��̘r�#N������G�?�m��w�C̙���8�-����#!�:�ad܃���ӧ���;�Q�K�洽mʿGl�.��y�-�!8e�Q�� �p�fZ�O��}����0�z�^��P�Dq�
���/4wM>���0*hK�������.�����.mN�� ��hm���ҟ��k�K�GA�?(��l<�-�pʴLRE�r���MÄP?i*&�q���E,�MҞ�������5�9HP��P<G�Æ�(D�Sl�wSff�1,N�VO�w='g���� ^^|'�V֞x��y�C���9�VU5y}��';�X���a�J��C7<#/��P]�����H_�������f3Vs`���bʡ�h��ct�����:�+O①������dD濫L���0����|���ޭ�?����h��}| 3^�,2�M�:0f��-͕JHuK�A��k�z~ۇ��=�l��_�x�lԘ؃
;�>q���$$+t�YZY5�1ˏN `�����!�愨"$���[-F�VNڪB��S6�2�g��Jh.~��E�lk����{���i�ţoG�n&��~���n�;*l�\�9�M�bH�ю���U�����B�~z����=�NE�ǰ�/���jO�����?#NY�.]��ܘm�Հ�y��!�NX��8��$�1h~o��m��	߮�;�����u���X�����/�?^�v��L���e�Vf�H-]V��.���3su�Vtj�����2���{~������?~{�����_|�KzV��V�>s�m�ee>	^v���c��n.��ߏ��T=�v�knk�P�(��� ~��^��fS��Uq立�w|��ӑ]���ں���͏�]>খD䄗mC|�28��a��CZ�������/�������U�Y�Ϫ,�֞(��fVk;�|j�mc!і����^)(�i*�9����t=�Ws��!Gio��LII�(��d_�������rp��Gh�ϙ>�~�d4���zUdQ�����נ���]wtOjߟ�������0�TƥDGK��e�e0(/U�v�c�F\IttMϴc2�@]əE�.uq���F{�V���[g0���k9�@�M���{B�쬛~��L�řk]������F7�ÄB5�#�i�E���g�J�n?6S]�Mx�
C�E�Л���י=���f�X�D&*Й���Ꚛ��U�o�b��0yu�ʲ�\��UTT�f��t�f�����<{����1�m�D����0p���=N����@j��n �m����7�Um],�����w�.u�Q+�tX6o9nta"�d��rI�Z4�����\���,����2"}|���2=B������q���awV�=>�	n����r���˓��O@�-��gV*�:�������c%�o߾O�@W��MN1/��R݄�M�ԉ���������1����ze �g�����N���R ����0�"���<b:���������w_������cD�g�����}���$h��ߙv�/%>ř�%�%0h͂�a9F[f��Q+���5(�rZZZ��X�ƒP����C�
ʥ���wy�:��/e�,3��Fe���~��̣å��C7�S��V�Z~�d��vZ[x��(uM"Z�j������ $��9E�8W��qa�8�j�K]�݈}����������#��,�R�i��Fmt�HϨ7r;*@��4��-�k�]�,�Μ�7*�s�2u�S���r�ϛ����|��k/bE���s{U��+@���02$۶o�o�0{����L�2�=�ퟔg���X�u;��1��s����H�AT@a#@%���n���}��w��\V�M7��tC��2qɖa��ŉ����wE�2VH��i�'���ݘ��Բ��V�dե�,j��ӎ
��eb��ᗕZq�z�O 
L��0/�n�����'խ�hZ}�D��5��Q(�dPn�|i�TR�Ǌ؇����/���з�?��{�`�S�� :wxl�֓����87�D��T�_"����f�};�x�\�F)�hխcN�QeZ�ʼ��� U+����4�8T.C����;`��&������:t�`���!��[i����8O�R	>L�4���ΝC?���
�q�$��Nh $q2��tl<�ZDC�%��^��Npsr��HVK0n�1_W�_�	��4B��p�f��U�3]�=~��핽w"lg3��=��t�G4�J�`�?�c#��#�Ba7�Aҋ��u����n�r/�����`�6n�Xr	�
����g�W!#�.�.S��:s�<ح� s�3\v�d4{pՔϣ�NNN5��6��M�͏�Q�'������X��p�����S���+vM����3�%��(�^�m"'���*uC[~��y�9����E�dj�q�4�ٍ���r֜�0+�N.�h��兗��g��R2�����x�B�����W�O�N@���6��
Nt�����95��c��-��JF���9ȃ�K���P�y���:�>ʑ&z[P皟��߹��.ch5��R��酯l�v@��˟\g�<!t� o�`�G�.�%oRg�u�ԾlVK#Dw�W�ð������@�˺���K���#����s�D���U31SLe<4�TExE�u�ԫ��Zt�<<z�V���q$�<�R9bQ��@�@���Fm��BZ��n@iAJ��jp�Wto���6���VE�I�,�؈�cޓX�OW=D�����+���$x)���fy�y�b�a�
�;���IU�Cϣ�d�Ӻ8QPȍ1=�y�pa������zGN
�3�a���}~�L�ޘ�8�6)�u�N����R�\�v�֟y'P�e)��!ޟp &c]����� ���Zv@|���z�J����V��,Ѱ�z;([��:�4�7�~�ŉ���#@<v���	D�ƣ����|��Am��cr�A&~�ώg���yV���ͤ�P��d�P�oV(�Qv�7~�	p`�j����~�nH�����#>y�|�	��F�K]�;ɭ���"U&��h+�(������N�&��O�c.x&3��������7�t�BV�Z^���K�*X��'_)M���5��S����\ �b��+�l��&����E��[2�	�D����	��{č����������F|��0�?R9��~�`g���2�����x��) ��2P�h��$���1r�PX�f����?__�u��`��>�Њ�Oޛ�K���ֶ���Yih�9�}�o�хGG4[�P��2��~�/'�\|����Ka�R�������]��UUU��~���3�X�8;�1�^�(f�q���K����ւ��fc�}����t�A%�����p>����i�S�Oz�MR-~�٘ġ;B�h�������P��K4竇n��ރ9[�3>�t�X���vk���. ���� /}��
PoB�D�0�9���^=�e�`��9X�,�;6��mx��v�����%3׼�Z^��� �ܢ�u?|�|?�i��RSS�/�i��Q'e\ڿk�����)�{4!#�]�i_���.��:���a���{?���=�"�#KN� ,K�0�^�'w���P��;�-�[���)�C8����yv����vu�����n9��-�v6O	� 7�M�*O:��*7f�Ƃ��#�z�G��?㧏�p+'$����L�_�9n4 �h<�?��xAg�0�<ί�0g
�����5�r]V�� ī����� b'�L�
u�>��B���G��Ї\t�z�|����y,���UgMf#Ĭ�-�𽑁��t�릂�J�'������YL{��0|��s���9���'+��v�CQ}�Y����|�rPr��\�7��R�k@%Ow`��^h�� ���]��{�M�$�"��&_���'W>T]]���$
#5J������.u�$�vD�|d��
�qƑ�揭'�}gY��2�ָ��Y�;(�|��0��ɬ�*#ѱ�I�b��ə�����K��u��o�M��u{�ۨ+�@��-I@�ː0vFQQH��-zO���Z��0��Щ{S�)4�_��Ϳ�<���i�/����PK   ��!Y����<  �  /   images/bdd7c0cc-86d6-4eb9-abef-3fcf444ec41a.png�YeP^�'X��YX�C�$�������;X�ӥCJ�E�nI%�P����o��wg�93�g���͍��Q#1����H4ԕ���v����NI%��g=�M����z��~'C�Nzcw{��K,~'7o[��K~w/���2���4�
	��bz.k��wx;xq������[�����H�S�^��jz,��D���K��
9��+O��,T�"K��B��l�&�|?�u���YTT��1�2������3�a�!t��ư:��4��ޖ�[�\È��9�s(&�k��������]7]�ǃ�A�})$�%y�4�?u^d+�O�����k�Q�b��쫛�'�k0��b?�����ckJ�,�}��+�Kd5��Ҁ`͜�FJ h֊�d�OU�Yz$��D.��Ff�I�g+��\
1��{F�rV�7b��R����	��b~���&()�Rz�(����,��0��K�JQLD�9�R*H2��D��x�щR��㷸6ΞF>��U��a�q�Z�$Y~2�By�'6��ZQ2��`k$�bI�������p{]����1 v��X��f��2��7m�AKQt���L�;�{�Ե��h����czBSiH�D��!Ź��[La�����;˅x~\�%�f��T�ϖt��ߞ��ǩ��o���m��2l�f�:������>bE3^
�{�V��(a�r��^�.�L��)C�5{ǌ��!�?�W���ѝ>cl�4'�p���؊�g3+��G+`t��n����^V�L��4�}�DV����f�Pj ��޲dq�"m��BP^���[7�B7�\����7�:C6�=���\IIvZ�\����]�������
v��vG�,l���=?L
�0R=ƣ�S��8U���
�d� �?��>�[Nƻ�1���sLP@k����<�oD��ZY�U�\Q��q�\h�]� ���jnB�uk�I�ōre���<�ǀՉ(��^��/���3HԞ�b�M�-I��%+o�.���׍"K����hFt����}�a�����iiC�����7}O�6}�`���^st���Ƚ\�aB���TC 5a8Ԉ�,J�s#
������#�H�cS5G�|}�2����6�B9Z�I�&*֖_:��-i`�U=�1L����ӎW�o���p��<D0Va��qC���"X�_�/���7��dB�.���U"ST��u�(�;RQm�<4�E��c]��?Xfa 2��>�זY!����]��\d��d���9!ɐ�*�ѯ��o�9)�b��w�iF?a�
� ?������wY[X�߶:^OL8�-"+k�Fp?�f��M��]���v.Lع�O ����pL��g�,��&�L�릆�Qk#�C�]�g���*�_������N�F�G���i!U.�JlT��r��MDX	��J�L��p%����ƻa��k�>_� @��$��i�G-���_e|!o�Ш.�x�I{�XS�[5V�<0��`�X
�	,��RԝD`��6r"��Ya�[Ǌ&�+�����g��������^k��qBT~GG���Cޫ	�7T.�%=�Q�k�~z���_ǣ�u�*2�z��p(z������L�zkļ�Ŝ�#�����
e.6�$��O����ެ��	ZQ|��"Yz�	Qj�h�S������.�}3�����E�i�-��䲵��0MR;���<]Rd�d>Ɩ�c
�P�w�����ЂD}���{���zΒ��2�R7����;3��������w����9s���1����g���glS�87�*]�y�C�|6�Gg�4Ϊ�i�j?�3��i�9JuxT��f��� w7k)��YLY)�l�#1Y�D��u�-���*��>��!�@C��)�h��#��V"��?��Σ�d�?�r~R�S:��%�{m�F	};��Ě�c�c3z�}7ܽSa}��g5C���f�\Fr5�
�B?���(\v�7�/vI�⧥	3bb�^���������"&��,u���(�~���QD ���PJ�L�^� |䵖>L*� �'��Ԟ�URң�Gїv�Z����C�|2&.���ܮ:ۋ@�UX+�fG��Dn�m;,�oC�ݗ�{��/�p"��I��b��`�Ӯ�[�nXK�7a���!�WIې��j�*����eЦ����V�7��|i�ܴ�����фRO��/ţL��B� M(S���~��GVa>#u�����ӕ:DD��=�r�y� ���zi�D�� �Ò<� �J��it�e��т���+-L�:(�I"bZ8/�{�F`�i����1�j+�+!��qJO�B�ZM��ww/��-5¸��D�Ulv��z�2��!��P��G8��ZT���G��4����x2�#=�k4֍����O���V� ���pбe�ˎb�ǧW\�0s��<���{���Xa���:T�i����_�N5N�(��w�?=fd�w�Ƒ�ֿ]�|8�j�4F\'G߮�xً����a]0j�*�By�����@��1�L�����
?C~r�?���n����j�{�?��5�P�.G(]�8I�i�*2F5{�#��]�����l�X"ȓ�>So�&U��Jg7�^��GMd�`�@hhw�6�;[��1��YZ1)͍y���ǫ�q�l���S��-tMM����Ry�_�hf��Lf2�����4L����I2]�2�c6%�٤լ��s�ha�Iq�y�)%qP������ڿ)x��%�Զ11�x^��Da�t���`���x��H���;��c��20q?hv�4R��|�A��TK��4�"�����[������h|��hyg�߮P �J�ߞ�=,
낊$�\x����k�����W+Ԇ����(]�b@ER�J����������/�X,ү��b�	x���Mp�E��L��q �)TTlٿ�+�RC���a����"�v����.��66��϶b#���X��yNı��U�j4���ԥ�9���{I/S��Ola�A���}��Hԣ��Yg��5��p=8�)w�%�c�B�xyRLu��\5S�I=���BU��wْ�d���>�JC��_[s1�p�ˮ�(�Mkd�*k(x`0y���ϼce��"�JrU�_�6����X<��?"����ۄUD�Y��k� 	|a�A/�zЛ"����&��45p{�wo�7���˗�-�Y�63�n&�\�G)Ekq�#��b��S}i(`�\椨k�o��:/�'xL��.{���ǂ?���(i��p���R�$*�S�e��ͬ<���Е&9����d�*+Z�\���5�6)+��@�O�>���#�a�5(�}��?&���F����t�C4��p��Y�ݽ�0Dwdz۹��)KNؿ�&D����Y.����ʊⱢ���=J/�
��S����U[7���-p�AR��@�r,���t$MS�����XrZO�?(`)�֭R�H�i����]y20�EU"����=�Y�Xܭa�q&i",N�ɵ���j����]���������`YG��3��ڲ��*�ػ�y��~{M��@� ��:j?Ď,�3��7�頤~��1L��"���M��!�|'2�2����ʩT�۞meIR�xH����J�۶�E�Ĥe�Sj|j�݅������ �M�frP������n�U����<�C����]��@3z��Z=8Olֹn(�Z��Z����/i��C� �dݍ�N�>$��4�yp��o�rO^Yۈ�ԻB��Е�ސ�jFɉ��Ö�VYw�K���6����wYg<6���ɹ�d;~d���j�e�a��Ld`y8w�/��W/��Bl(h����ū�&�ATA(}�W܈��MIpT�>���m�uq� �l�^����R(]|��ݮ���i��Z��x�j6�j�L*�~��
�d�ꀯ�H��nq�G_2=_�螄�� ѕ7x.C��nyq$�R� �Uv�=eHF��cE�9)Q���m�M��&^^G���"�W#-5��x}=c��5X:7v$ԥ�>�,~Q4-#n�i۞�l��+X:TV<�ѣ8�xI��ε� ��Hr�3F�S��5���B������uQU6��Q����9"H�Zzk���l] ����4�K*n$��fg]:�%��ɹ�]X�Y�e�l^7}������hU�f�{�=�
M�r��^k,�^��5yn징k�Y������^���9�v�x7�~T�g����ʫ��n���p_�ʐyZ�� =��P{uz�6L�)�E8�����+� �^�h������j�UOs�R��t	�Y�\�J
����a� Gˊy��Q�xqq`I�~ 4&´���#�k>�M#6�Wb"w�����ڟ�VP�f+��h�1ֆ��������'Wy�6P�ei��Y0���w��L��@��ѱ0O��(z�p@U���`
��G~�Ӧ����pI�R
�f��F-��T�<�a:2%�^����4��
j�BP<�����=�&�W�������tn���y���1Ƌ�QF��_��.�8�s*_�՛�r��w�JG��Պ|g���+9ho�����9�ۙ��V@�fz��ȯ��u�}����Xq/k-���:q6M�H�欨�0R�T��q	�M�xf"���t��
.�B������/�*Q3����cẋ�dN���K�ǽS�bkFT^���"˼�����!kY]sQ�O����?s�r�U�G�a��2�^��ߥٹ���D�����f�p�ƌ7z^��$s$U���s�sfW�Y�+�X٫����?�SxN�;�� �%�L���yrny�e����`YNZ"�Ҁ�>�TEp��,��f�1N���DR�sD_~b�]�Q�|�`�6�+��bF���+kk���o�FV.��%9��7��}�G��n9q��@4.�}i�ܾ����z+l6E}��`_�,���V�q�o�up�e�� `�U<A��!?�P��tUe��u3?�q�"ʭJ®���@�TP2�s-p���,�O�VV�}�k�d��I;r�u���eOCơ���]�1��3rZ�l����q^$��Ǖ�r��D9�׭<EH��c�����'Mm�5^w��2�����}P#=l�1��I}�����꧵S����-M�d��͡�2�� øL:!�H!P���@ټ��ru}���:��S�s?��t�X��둧�bC=D|�5U��~��b����IH/��Ϋ>ݷ����Kc �J� �<�j⾔"�f~̑Iuҗ����C���"թL�C�_�LZ@�����זxf���(�В.�y;g&Д����P�2��H;�N��wQ].���t����J��XE܇���SRT�Z�j���ˮ�M!o!� cLS
U"~u�P�N�˻q��%o�~�"�a�����[�:�o��=�i=u��2�lHH'*�����͙��ï�w��H�3��c'Q7݉��������m��6���K��G{aK�(d��R�w�=��?�_�G���X��� ��Ǐ�&�' �5)����ߠ�œ�	�Q1u-\�5���x������������F���/hʤö��~ʉY��k��D�~� ��,F#N���Eĵ�����|X�=ԁ��'%ѝA�A��m�Ч��[�l^� ⷱ�����/��/K[��_I(��/���U)�Q���2w�y��mr�z�Jc��i�W�o����o��Z��fO�oi�6* ̳3Z�|��Ɩ��I�/���������4gt�S���~�aɒxn�6A����V��5S�5�=ZeC�1�W�S��ly�(���Z��K�r�N�C��2$��"}�g�F���N�u�hI��UZT�Ǘ���QJdgl�3���Z�l̐���&��U��?x��|���@��L+�U[�	P�i�U���Y�ݧKG��̡c��K���"��
�q�m'�T+���}����{��TY�3���/�z�Ș�>�E�"i.�z��w�����cW�1�o���ݴ�r�9�6�.?8���Me��*���?{A�E��c�bL
n��y��w�Jp���Խ�O��̷���X�����������#�T�5FP��b�����N�gO=3��+.�5��;�>��rɿ����=���'����H@��}N��U��3vտ�,�M�oTK�cX��VU�i����X�?0z@U!S+X���Зm���i k���O�Əzy6�x�",�XJWuU(�/S�����fM��F�������܌6�m�/(�n�Ѽ�ĉׂ�	�1��cf4D�#�6�lͫ���L���l�|E�
\R|�=珿_�Æ?1X�V(V�%7n�zح�*F�6@-�'�o��������*�����R�bϸ�j�Y/!ojݵgl�[�*E�
 ��Х0/��A���'Kd�+���^�,�_��0v����w�_�˝���~!�`�u~餍�s��x[�v{�Y�۟�8� �z�����MY�k��#Z�Wr�������N�vS�4���drI������Wh�,��ԋ�X�E�U3�8@������%2+�j���%������n��[)���+�Kǁ��3q �?��^֟u��N�S�N�Y�Ð�\�"��RQ׋�['��#�1��^�r���(�z�I�]i���4;2��ʙB��1p��[�Qno
 Q�+��u7Q|}g��lG� l�=������Ce?��޳@"_�L��X�l~~���Y5����?h�D���bD���U�a	��3��-��ۥld�gH��r�ޤč}�F���.�Q��E�i+$?��'r>��i�}�_׹b��Y�V�v�s����_�nk�J"#�N{h�{7}u!�����n��R3�s=|����/��s�˩@^7M����=��=x�級̢��a�{�.R'ٝ[ً!�!�L1�(�z��$z�����]����*�&��ŉ�T���1��N�3n���c����$�@��;�-��=�q�x�#�:^1�� �T�_�%`o}��?�����&2�}��:�5=����:4?�&���Z�&����:S�,2-d ��퓼Ɋ��р�JU���[!���{�'�gM��2��Z�}Kr���9��]�P�9��Ac���P�S��#�u�n^��sN*���à^���7�	ߕ�p>�l}�ӂ���Z'R�y��E�e�/'b�%@��3��Z���
��.����V�A�H�K-O����Õ�n]�it����6 ʆ�7Bo�'� �5H�vl�K�F��=Ԍn �F�c�i���̎~\���3�/"Z-���8��3p�z�}(�L�"|tYz~����?Kj`g�ע�		�
�x{��;s�$u9�+�Ĝ��|���}�]�
���׵X14�9�KO�E��=��?w���p�9�{i�ks���oip���Ww\�\��{�"XA=-c�b>����ǈi�����f�ǜ0:���sh�;����QC|+�U ���B��	��O���H\a'�N9%�[��c`n�c�N�rn�����۞��:�f�h�n�[vZ�_�)r�ۚ/1����S�í*	���W���hp͕�?�z­�����8ڸlx��d�i�:��/���zE���PK   ��!Y��g)�
  �
  /   images/c1fb8ae3-abb7-4800-a199-c8a1e0562abd.png�
!��PNG

   IHDR   d   B   �s   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  
kIDATx��\�k���߻��d�dK�jA4F�H\BK��N?p[���/�C�P(n�R�?Ч�ҧ��o�@����UR�QS0�cl�.�lY�W���jwgz~�=������������;s�~��9�s�LBD�O�<�D�B�0#�R)�L&E�\��j�*����$bϞ=b�޽?��o�YLNNv���#dvvV,..�l6{ƶ���,�;*��!L
�{t|�ɓ'o���v���#d߾}��ݻ �;��n��������W�92H��I�z��h7"G�Ç�����HR^V�h���e?Iȫt~���Gt�#�l� �aQ�>�����C��m6�����F?�jK�Eİ�~�O�^����/؏���m��\.W&���������!���bbb�P>�o�V�#D���������
gΜ333�T*}�:��'��h�u��3���=I���b��	D��X,b���v!�o�p��
>pR���={&8Б�G�8u����ܿ��D��d)�N���3�������;�������"GM[1�] ��1��$ #.;�|�����z����N�:ձ�G��+W�xvg�1�T�P�����uk꣏���?�޸q�#m�!Q�sB��	�2D�uP�7a����;�B���MY��۷E�!�<��!��aw^y�uw��!��:>�!�t���'�����ѥ�·��"�Dx��dv����y�cc��4.=�����vD�t(��[YY���L:$ ����d��w���&����(��P[4g~��='d���.ҹW��&�v >YU�&�رc"N����0��r�:�P��ᡡ��r�cI"J�&vtx=ச���?9��[u��r�DMOOSL� cy �H�S͝0
�F����ˁ�V'����>H�#�0Hm�I$(��. �	��ras j��J�!���_��x0�u%5�OJ�*"0!���h���������d�C'.-/c��*O�m�ȧN�C$�.��:�UҖlo���˷b��ϋ�J�a�	�H�(��!��m^�0����͂���P�\I��!0!��8#T��`��ُ�2�F@����יt��,����BH�������>̕4��k�@�jnb����ٞ�(��5���`�7
�)!L4�
��2�'�G���SL 0!<;	�Ӹ�L�I���	�t�2Sf�~eɝ�a��`uez󃖄@l��4��4! :�7��,��U�&�B����4��.B�d�I�m����u����*�ج�;o��@�����J��.�v@�=��>h��@+�v�����κ�iG�:.!~e��< ��?M�t��ۅB[��݃��&o��|>��:jbB]uBM����9��J��!rX�"š��;�{����G��6U144$����V1�׮]���T�g	Q��TWu���ctl__�$!��q�������c/^������!6�����t��9}	�"��t��gGVΓ�;$%����~R}������{cjjꗃ��� �7M�����oY��3�.�:nCԭ��N�w��Mˉ������$=��e�))�f�I��`��X�G��g"�W�.]�300�aGgY~����_Y��� ǹ��s���]�X^��xNrT�K��xK�V�U���1~�lB�y~�h��Ż���;`�k\7�Ћ�Pw���z;�M���8-T�JKH3R��dB�`9-Bt��mZiK�XH���u��#=he����K~�/�-�D�W./���4�W$;>�m�����x�r@R5�|n���!����!��U����9�V�??�mC�H��u��W��Z�F˄�$��i���v��V;�����*�<���cx��6&��sq���"F�P��':�`?��OB�#BxB 8��<[Ӳ!��� OL�#�-�	���dI�+�I��ȟ��6ꬲ�V+��2	Yu�/Gk���5�!�kE�C�:�WiYe�yΕ6��D6��m�0G����=�>��C(���5ǳ�Q	Q��F]U���!->Hû�ePG㍫?Y��5;��S	e��T櫵r��)�#B��$�S�����E+���)���-is��CTP�Z��~�����6|ޟI�*"	��B_��7)��ׯN�<�/����9�8j�!�mB�0��Fj�-L�Q��8z�lI!vw�w�f`qH����fg��ŭr�r�5 �~��Y1���������+u \k����u�a2!��N�:�\�{�m�N)�D<�X®�˗/�x���m%>�QZ*�ga"{�&�JHPpI

+�Lf�}�K����و ]!!rX�$���Q3ݽ���9����SHR�I��%�7Kk��d�jB�3!�&��u��&�p�~�\i��E;�ʌL��l�I������#5C��l�oT
��m\;�]�����׌j1M��BB,� �
��8n��{���!�n&��Hㄔ�ٯݲ7^v�Tn�qJJf��,�?	��{6M�]��u3NȾ�����<!j5���%���p�-�M��m�	+�z�R�,��	I���<dD ĉ���P�\+���:�nW���t	1�.�T�R9�n�B}	q���|������۵bص*�
���7K�X=v}��P	�?l��v�l��k0xO�n�����Wㆰ�v    IEND�B`�PK   ��!Y���]  [  /   images/cbec1558-c992-4de5-91c3-4ac90e5ffec0.png���S��i���S��>�����TJA� )��:��8I)�����Ox?�������~gؙ�$���@ �����#_>z' �1���<��K������������1I�n�g����q�~�����r��q�?�g�����VS1*8($Me�^]9�{ؐ���D7-;��ݣp����ԸT%�Q���%�B�ބqT��|>Z::o��x�A�4�3:߸�(ep�t����� ô�r���7�][7��G�ч���e��Ӭ��P����?�����dޏ�+3� ��O�W���U�����{���R0��Y��,��.����/ES�X��㺐��7���ZO���qlll_I�
XZY�ɩ�������/�?�?Dof 1�͏��>5U6w8��&(�l(�K��*�iyH��MU29��=�,���N�z|��;"��sQ�\BJ�<P�����kt�S"�*��ǘN�F,#�O}�T
kO��0?��s\�#������k(��u�д�F���]:���	׹b�w�)�5��b�r���D6x���NT�n�O��r�f��a���������JR�1m����СUPJ��1�6_��]���~Z���.����B2��Ŗ�
�S���Pp$q��%�O�k��[�ph%T�v<=9M#*����[2��}qA����h�!�0TT@���IC}o����	��� \Wv��v�霾�n��G����H���ե�ہ,2�D̍�Mhq�p�A�c�.P�~�ϛ�S	��E�F�,��J�:��@�EA�=��u@&�I�5���o�sg���J	���q`\y�#t+K��7��&8&�s8��$��ag�bY����L�:)p������m��9QG n>wU��	1cYNoqc�������'9����H�o�����(�:��_y��YS'��K��($H�XJ���Ox��\0Kr�DF�>J����z�?�7E�:�0������If��'S�6����Z��j�)��qZ(�>Tѻbz�_�J�K��sX��7vF�T��:P1������vf�C�a��+��,dK)�#���@�dy�\�ͫ2��zKB���\�,����2r�<�_u��^�U*�!��6ut-w5����e	L��)i�KG��I�L�r�S���`8?E� xaaV]����0���k�\&W������s�ؽ�*�-Y��U�=Z�����[��}�xOy����:/�P���r��s��+�w��׸�b�bm�F°�(�hj�l>b�S5��)���3��Oo��/?�?]e��F�_4T�R�0�}�u���{���iѱ�2=��CS���rLm�w��TA W��5^3�>����w���bܪ����%y"Mj\�2Zim������_�$�p������~�����~�:�������׉����w3(M;�ᬣ�L�GBҗVp�i�>�V�\.���e�êJ�/-{g�>8Z�w��E��O����ȴ��N$
��b��~���z����>P��לq�И*��L���ka��BƷ�'���̰1�W�)�у��#�|~B5w�5lX� �2�߬Bo8�s���h�I���ٳ�Dՙ#��?���:�Қ��+&�6y���hk�[�f�m�b��=f�� {�q� &�
ⱊ%�Ɋ��s���3���ט#�HA,��Ӛ���"�~�8�����#���q͞2Oz�Jg��`�"��*|\R���|dÙX�z���Q�Q6|��6��𱹻�����=�baf������������w�� Ip�8WB8���9��Th��ې�<*Z��/��' ɶ��7����d��� S�//Q��O��e�O���ā>y9+UJ!E�qg��:u�����5��{�������=Ҭ�Sd�l}*V���݄����aQ\���P��jO�+���3BѰ��:Y@����a�4c���ys�x���e���{ⲳ��n�mg�n#H�c��A��`�^X+����7KTVV���(O���熇�;�6^EB�1Gtaq�0J��m/�74+���%qF�6
�>Y,���ϟS���b P��O��D���H�;/ܗ766�m�p�L�a:�u/:*,$�%#���De����L9�a�M�ۓ������DTr���������z~>�s��͘.�[L�����͏�#�	nb�,i�3���7j����j.��v���5���WB�@��f�,��,rc!�?��αuZ�w]^9F5hC�444Έ���5���32��8Y�����S�l��[Q�d�ǽ������%� ��N������s��	�����21��33��#gg�CD^|�y&ʛ��E�:�e�����T��8;�K�;I3�IF�d�-gE�ao����z
a;}{rrrXUU�ܦ(��XFN��<=\ٙ�+�\��q���pR�{#&&��������&�M��� U�lv��όD"�!� �z@A�N��Y�j���_��^yz�>I:5�3�'[1b	�3fiJ��Wb1|�J=���gs|���"VK��II�p����w`[�ۍ"n�a�'�^s6����+�-rF��H��{���u:��d?�`6�l���$��`�O-5ޣ�w�LyÚ�t�e���ί_�����0?d� �n?ɦM�;~�}�T���-.����2'�z�Z��zS����%I#Z4[)���AR��-�j���z�/x^P�|�IR�Zg�5�ҏ��S�w�����Ӻ1@�V���D�JulM�z���>2Oo%LX+�IkЏ.��,��v[��0]vv�z�{$���P��_
�j�Z ��e��D���#�ͥj�oj�z/����6�$��n��܍p��4�D:g��'/�Ϙ��h�����f��[�We�\������N�+a�^�PӸBbXE ,D��*UPV�D} ���L2e���|�L�5:�Zjim��S��F�,F�E��w�B���0�ߨ����6�K���MS��:� �5�A�__�U!H�d��q�����1�M:��b]I�svVs����2}��a�7
;��y?�7�����n���Z/�Ifz��݁��/�*,5L��@n՛�"rT�[%��Q��}MpRG�����Qj�=1�=����'!��Zm��5���������!��U�>�#�5ߥ�(3}O��[�t80� a��P������-��Pd�����Q/��>O�\V�~��v���奦�W-u��5b��Z����1�i2�s�/_�P�����1	G��ks�"r��7�%s�jYL����_K�C��ɟk:l�����Ù��sP{����B��	xkJ{E�Vn�ί�_�4Q�/���/�uY���c�����cZa,ǅY�-��W&��]����*�n��Q})뵠�-+	���ڠ� �"SS���	+�"o�o��{G�ɛ���2*+�d릑�4�Y�ɍj����?KO`�Y�
���p�I���@��߄�gb����9|��wSp�?<��=�}�:��d��S9Փh±�Y�f�2S��ͧ��0�2�ܚN~�|W�I�2��b�PU�5�~��bm�F?�	-�V�zY��.\��U�S��veZ>��L�k�����������is��^��.���yz��t圕\�H0�3A,z�:~�Z�4�5*��Z��¥�������(;c�9�V&��"�Aq�TΠ�?��,e	��i���c�-��¹��*�x!F��Y\K��1�N�!���<�ۨ፩�6��4��'����K]Q>�<熉w��V=}��O<5��.ˈ}�}���y����b���Љꉌ�rdZ��.K�4�w[񧾿vf���pq�]@�e�me���3��޲G�zCBc��6�J=�|a3Ύ��$-��`9�w	��uT�0�����QaNMm0�H�5�[��DD'��s�!�����j0�6�ͫW;��YՋ��ͳ�ɂ
���a�7r���n~:Qفs�YU@�]�������#�o�$��/�Z3by.��R*��w־s����&QU���p8<
�S]GW��7j�Miˏ�-�/�:��?��Y&���*�R�̤�v?=;��В��	�JHHX�*ڍ5*�,j-��� n7������1��l&ۿD����Y�M����F�a�L�_��=$�K�b��Չ�}�n�z���O��E�@][��)�>�J����<;;$e���3.#���Al��ǿ�0���J�;$���:j%��'5h-�v ����<0	�4z>��e�r�A)]m�k4���[p�~{}Z |'>���#L�jll���W���%73�3����L�ޫ{YJ6~u��0�L�yq�(�,���r~�|4������Pͧ!�/��#�$XC�j
����o��(A��n`�ʳ��*
���&�?���Gs4]o�t9�	��zyOH�ˋ=��×j=��Bv���&��5�߭?�:	�� �� ���k���i�L�E}Vn�Y����ϗ?��'�Vo����{X"���BM�c4��(��L鐳�@����u1#>ǧ�Lm(�a)�RXۆ4�/�~S)�
Q��	@ӱK�ISe0�pj�?��;���fS}(�p�?����O��Nl꺲�ɟ�U���֮��6C���3�p�v�i��8�����p��)k˾�Iqc���O�	R�-�dy��k���!���T�tI1�LG�*�w��)z�]y
v�\s2<*��bA�IC�.Đ�����	n�!�wd{=����ϰt�E?�<R�w�_����pE�Oa�T� ��6]$r���^������)�~e:Y�&_� ϏH�,U:��`��@-�
���Fӭ�M*m�Z�X�Ž�I�4�C���b�P�AR����.�=����5��I� zÏ�=�"�	WNt�5�z�L$��Wn@�Ḽ��K�+]�_�"Ti�_-h2�
?��(�K��0�JG׮`�H�r����bGu�#�J�TJ|Ww��8\Wj9ͨ�~,I�b
c���M�Ƒýaxh$(�6ģ�|?"�l#ļ^�w�\CڞGpV^��X�~ۯ�	��.�);v��ZZ��(��ZH}O�y��[K��>S�垎%U�!t�,�PRjg�����#�pn3����\זM�H�"w�?��&nqt8��p��)��W���L�p���up-������t��	�ęշ���$�gP;i��C��u��w�OKn�S�W:k���~�4?#S-8<2 �֟\����Ӭ��=�D�>L�W��h�����@1�PK   ��!Y/yR�c  ^  /   images/d2af519c-c065-45b5-bffd-6bf239de2b90.png^��PNG

   IHDR   d   P   �	��   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  �IDATx��]	l��gw��c};��ΈU��ф#H�4�� �U�R����HU�V�z� �rD4��F��\���І�p8�Rb0�41���X������lf{vv����>�g��f�����������*�8ˏY&�d�xY���/�m\�BQ�6��#���a< )���������������~��f���rݟ���M�s���Ȳ���x= �IaB�� Zl�ۗ��������p�I���zV��ˊ������۷��v��/����,���$1�#L[ 	����t�ҥK���_����Y@NN�;wn�RRR�_s�â�Ͳ�e�[,>�7�AI�5DĐ�ˢ����I�&��2�M��	b���j����͇��cg��3,����r�x@c�0!W�\�[vG�p8���/���#�)��Qr��>��3L�9�e�OX6�FN�^(�1G����:joooHKK���"����.ܻ�e1�wYv��(�S/��t����P�������;D\I�Y��;,+YvRT���h�p�Ȼ�������Ғ3x�`b����M	��*�?�4�@�!�R�?x;��������/4A>��E�Yǲ�4W�{��(�ۉ	2n�8:~��~XŁ�Q��UWW�C��������Y^e��
&c�MFyy9�]��� e޼yqՏ�#)S��kg%���㏗s�=m���Ɋ+����
?o.?g3s��qLA��À�"V�k_�n]\�8�OI	���a��ڵk�9+2d9�N�&�|ʔ)t���)��@��<�zۇd)R�)���d�x���F�O��dgg��W2�T[[K���b�-�b�O�>B`�[�{������p�}RC&�6�gXo{�!��
b6o�L'N�S�N�p�]�}���Ni1w-�u ��ѣ�\�������h�ر4|�p��ʢ�S�Ү]���=�R��`8�)1���㡊�
�Ng�QSSC^�W([|���)4!H�"�T��u��bK�)wYY� %�� ���w������1		qdCo�B�p��R���L�'O�dXq;x�~��i6l�p�S���t����DEU#�)���y�2��SK��י �`\o���bU��1���@q� �Sc�����̌���A�Pt�K���7n�nJ�S ��Յb��[dS��o��f�q�V�Q��2(���]l}�4Q_?F�~l��=�������F���u8�)ܛ����R�2-�W�^d���is�uD�NXCC��5e6�u�LG+=9t�;؅����j������)/�y}����D�?蠃��G��M�L{��P�/�f�Iv[����-���p��N+�n A�&��y+')A�ج]J_�p�-�c\	N
̘1��/_N�������e��	VBA.�qd�̙��~I)h�v% [�Jo_�25ys�R���ug;=��h�����=[(1\���TO-���������tQ/+��2���Y�q,��!���l�U�������dy��V�WLt9����'��IA�0`�Ha�]�d	m߾�������`�cdn/��M�0!|��W�
f$�G�|���B�����a�r��.QN���E��S�e�l�t�(��9?�f�n$���,��4�jNO��"t$-�����A
Z<�pa�c�ܹsE9b\Z=������D2n��Ѱ���RЪ�����\A{/L�*�B߻<>l!�*զ)��qd�����.�a�7wO��n�f�=�<����nR'F���@�$��R��"�����/:yP<�-V�.�0ta �3���j-]����nѢ�lXHt�bq�C5����
�B�c�X݋Z|Y�V�T�����3�x� @]){��$�]`�� ��E"CF�v���`�޹�yp[pu�`�)�6�:�.�f����.�d@y(3[Ay�禋Q'��]U_	i�aAqA��ߣ�=�v~83"�{�V�,��1	]�p9P0������"�Bl!dVp] ���*�!��9���6_F�֔��Q�^�}(<�Z(�X'\n8}M��(
�Ҭ�4��2a!p;��mA�1z��gg �
��X#�fʰZ�Y�xϛ���1	ٸq#Z��髊1&��D�(n1&V�n��L�����Q���ƾUg�I��Ç�Q0��p�BJ��;!2�����X �C�Dn��ʕ+A�ZZZ�$J���28�T�y�f�}�>~ժUaRt%n0��TX�c<^!�,�IQ�u�����%�@�#�MT� ˈ�E'����6�=��z��B0�٤�H�L�w����!��	h����A���'�ǃ�	��SIH$�	뉢����!	��A�9�SS̰x�bw�@�u�������8����.��$���Y�9s����e˖)2�Jʃ>�zNN�M��֬"yܬHH�oD�F(�E�`�A[˒��e@�1;(1	n�[E�#�$����4���0xXPP�̟?_]�z���z%)2�?�p�\J�\��G��`���eI��X ����;��Z�;�x!ř� eŊ����ۡ[�СC�"p��c�xԨQʢE��M�6��d�HpV*^�q�UB?7�|������*���4�u$?PLՑ����<v��1hXb�q�̙1�����o�6��i)=�f�4к�:����yx?oڂ�0�����{����z<�=�-2#\�F�H�{���z	�~l����gY���O��h�uf0c�����>eVl}>�d��K�,ccU��P?z��k�Neǉ'�<�	E2vt����Ԏ��[�n5�V��$!�!:
����$B�/	I!��=ѧJY�"m9^,�!	Ijk{y��?��Kښa/��.*bJ�$$EX�tӫ���XxlK�dXb����t30��fڲs�ӣ�ZX�f	o�MZ/^ZH�C���늟���w�ÂD��&��$����38�MXXC��XK{5bU��O�諟It'0�T�vMu0Ȫ X����/�~¿"��t;LQ��'+}ݠ|>5�4��e?�v�߰%���?|饗���nX��,"-��;8��,{YvKBR��_+��wi.��1b�|IH
�ي��������_=�3�A��,��|��Q�\IH7C�)��+W�~��XO�e&��4ik�1�=����nF�UX�h�ol#�k��W�he�g����-$`��0���RFZF��F�e-���PW�`�ΨQ�^����>Â5��(�|6*<,	I�m�ǌ�>��e�|������,��V����ǉ�H�B���z�����_��V�B�0�.�|�4��$|��9IH
�q!n|���k�}bj�UB���9�X��]g�0�����V	��=�Y��D"��Κ�7�,dYb�|����$)�d@wm�����0)O��)B��fA���u�u��l��"��`���N���x�]?�~���&�e�_w:�x�$$�|��#G�|�ԩSq������A8c    IEND�B`�PK   ��!Y�GDU7� �� /   images/d628d844-ce42-4e82-be63-f5fdfa438334.png�wTTٷ.Z6ݢ�@w+���6�d$g[D$�䌒s��
[��,Qr�PD%I���"�Ud(
��Cy��w����1�p��[ٵ֚�ߜ+P��T�~��+�����1q����u�,��oT���g�����{��%���Ώ�����3-6������k8Y�#��Z �H$������gn'W�D��5�O����5���?�9t	��T�;N���h?ڏ���h?ڏ���h?ڏ���h?���-`�9����t졚֏���h?ڏ���h?ڏ���h?ڏ���h�W�����w�>�d��c̯��nq�������\<W�^�)�����WvK��[���<���N��s����vK`_���jv�z�n�����[�o��p3�=E;G�oZU�y#3�{��4�.�����o$��0�5"���x���ȏ���h?ڏ���h?���Vh^���a=)n�$�pX޿���g�\�+S�(�6��](Ӏ	�N㱒�w�'ӪJ�����K!�:Z#�|��fXN�Ĳ�_���F�cv�n�|�؝v��T��m�"���2��/�r�f
y���f��XH����S�V����z��y!�R/󘭮3���g��o �3����Z]fk�>�)IN���;���n>����9�}M_iX�X
$��D���������+��\����4�ͩ<Ƨ4Ƨ���)?�Բ��W�`T�SY�V��o�j���$������eObՕ\���Ն'�k���_��_*K���5�\��ubK$��G�0 ƓT�g �\���	��i5O<�yfMQ
%��ޛȻ�T�����ښDq���F�{L�ڈVav��>Z�f���Ԑ���dC��^��?���~����~Z=Ͽ��%.�
�d��m�%����_�)��$��e�9��LM��#����s>s����4Ҩ�S�n{��)���i)���;�z�ֈv(�]sh!:�v��|7����e?�o��O{�'�T$!Ћ3b�V@^n;^Z��K^~_jҤO{j�/kM���u�<+F�K��)��{yY�T�������^0��,Sy�/x1j�N`!�X��6'C�c!sB�]����E=	��CMf��]:퍹����jؤ�gq��c<�����Q��.V�Ϣ�e�C�J�TʌquoA���Gs�������3�9-C�퍽.��>�ٞc�}���E�'���q���~gJ��^,�)G�M�O=&KyA,�$k5�呕�������.���5�9�Ӹ�?��6 �jf�����5��� ���˔��l�2[���	x���r����!-y�79'�f(K��Ȉ�cl�� ������]�R�?�g��EW�󝲯�l�]��B���(�	Q[�%h�yM^X����/{�kF���Xy�ZӤ|*p�W=~�
k����N��s�?*�K�.?.�KGi���>4��w��r
�C�'�8ܖb��W���Ȝ"iIS������)�3���/�c�^ֿ�����?�;�,XF
��ߋ�T�:e�b2`ȴÏE�n�m����.	��Y�Cj-S}�22���k��ͬp��@8A�(^Z߼-�H����$u�l�rg�a��,�:2#�'6���ϭ|��j��^�>��=�G�O)�*Yf��mڎ���FT���)CM��4Ly�'���>G�=:Iqc�0N����M��9{��I~Sf'�߅�=�WV=�,�9��Bed�H��Hbל���KN�%{_/����bo<��K�X��0n��U�����}��8f��
h{�춡+1#�f����Q��!Y� �!�~9/{
V2�����qK
n���X8<�#(c�!(O��m�G
� x<׎���������W���Q��T;4�����3���~6HB���ۄo�.��BF8�l�0��ܹ��G�d]y,��Q�Gx��8�oVSR(>'��q}�%�"�L	�5�#8���R��z�����`K���t��AygP�����A��yB�#'M�S�=q<�5�t�N#=�� ��|t�t����tS��r�w,�h"��J��\��.��mW48,:r����[C�":�ڠw��ˤ����Z?�������DIx�j�s�Fk)ec)��!#�矂f�e����ؐ :�7�&��l3� ����	D՜����~��x��`������BM��	�A��]���&�R��l�Q�ZD��G̅�,V�
�5Ͷ�"�&�����F�-�4���Țm�&����6�\z�Y��8������WF�y�×�����٤3J@��g5��ne��ʧZ@B'=֙��(��QÆ=���u"��ƫe��0����t�pt�����(�wL2Z�B@#��}�ݯ���HЫQ���Y�k�g%��Ǹ_l,�p<~�q���s�U��	�����<��k��9�J�7a��%�ԉo���y,��v�*&�?d���\͗�o�~�b?g�}d�џ�S���X����M��p"���������4�d��<k�z*q�A[���R1]��h��Ē��F.afG�ec/@Q=�mt�|&�caK��q;������_;�?#m�u��I���*_�U�+�ىPo�<�?��9�
�:Z%Y�G���6��^Kt�) +���/Ol��S"N[ɤ�~h�d=�n���;#ЮB��C���I�����	�|�`/Na�z=�w�s}�#q:F�����d-�F�\�b�����r;�kM���d�� b�B�q�
�hd���ȡ��k��5��]�Z|�F(>� x��+獩���"��꽡ͲZ�Y��:�m �w���-��|J���:xH����rC�p�b�@#���+�2sy����Ȧ2�וAu�"[�y�Hm'��};���� 7����z6-�L�ג�E�V�5Z��,S�-���9���JEF/,�hx�4��6�T�cޜ���z~��j���I�oGNoS���{h�͛q�v�~BW�O���	N5��≡p���Qdw@�?��	��¡�9Ц�PL�u���9{�F�v��k�z����iw8��_�P���5�@Pkհ�����_���(j�����Ԙ��5e�5�np�`�':2{���`�/���fج�NwbĂ�Ưz�����drQzDʆ�����u�B�N�z�d�{�T��9݄jy/��v��F�	��G	`cS�����-Czk�<38jOM!n����RKg8�wZH�J8{>�a�r=��^���ί�i��g�}���k1��Ff(�D�=�kQ����>�;�m�x��k����|\q_���
�*fy��ZDK����R���*i睬��I-n{+�y*� �X5�Z�Ū�����|��Q��34ఠ��0���T��[��P���Y(��Rr&�6�!��m�J��kV�])�f��t���?��n?/���`��I �f�����X.U��_�蹤�O/���ʻ�����X��¢ʚ܊��E���*�ApZ���<&�
��9����ƻ_:��6��P=�"���OD|�}�8&3���VT�x}�>a�}�ԑW_�7� }��]�kP��T�,�_�$��J��)���>��Ĕ�����f �r�:N�������gf�m,�&�h$�y���AM�% [!t��b�hz���$�9U\S�Hַ��7�©�����!���m��fs�%���}�n��:�ǖ𲃃߾���Yd�X��݃�A����I5�c��Қ� ���`�y-�vG_�F�^m����q`���U#&#�>0�λkK�����tGP��_�@�'"`�w�	2�d`�NBv���e�����,%�q��+A]��X8��tҗ�a0�r�	FU'����� ���K��%N�A���B;��w8Y\��u���ZB	CBl�Bi�T}��4����!n��!GF> $J�v9�v
����?Ɨ��qF��j���_��CwW�zl6���ԛr�@ 'L'gY���?3��O ��`��*��r�� ��W6%;�VzO��~�+/oP���1z$�}B��'ȵ��%Xc���@τZ��;Y�Di���ݮ[^�cQ�SYv�/ݰu��.�V"P�V�!�Vˆ��h����]�MM?�%uN(e�.�,��l���[�4q�+�oON/�] 0�޹�f�
�x�V������i�ow�Tp�Y�#@N��Ax)���.6�!Њ�;X󶁷�}i6��XeH��#�D)�}��V��k�Sⅅ�D���v�U)��$�����P�c��_A��d�,FQ��E�5����&�K:��s�g�&Q�}�da�aay& a/� YO���F@�$�I�&�#c�Cy��&�Z�u�x�Ƹh��~����/�1+2���%�Gx�%_z
ՉJ���`*
}���G��n3�,��$}�~�n�n�Y��ӵƷ�G<&M[XU�S`�:)c��H��#�_����fd��|ڝڷ�'2�;�\,�jP��� ����0����:�
/�dGGZ�!�q!׋�&)G[q�9)R;<��SNb�ኇ�1����o��>E�&!�֡��ޱTc��F�I������s6�s��R�<9Ҽ�Gc���	����bU4�/F���1��V�.��~m]p?��������� ��"�,sٗ��F;�QBF�=a^Z ����P!S�T-'�f�8����A1݇�$*�Vf06C��M�ƒ�do�A��R��W���fc�3�> �m�wq&�\��e�N<p |n Ӏ ��3�:�f����r�"ڽH�0n�;�$
@�
v;�Ku�H���j=���-��_�ç���F%˞�7\�PQ5-���!�n�"��?�?*�ҷ�-������P����_����Tu�,��?E*}�5��V�.�p�#v9"���3�%��	�R
���'@�Dޙ�����M7�T�o�X)�Z`�����ܞ) ��HX���)�/� ���i��jʨTt����f��e�?@���~�هIo'�)l�(��..y�1�yǔb���_�]w��{{�[]�t��4����N���K&bȓ���� ��]_!n�u@7��s��eW
 �V�E�ǆ��_�;�ӏ�����HR�H�c��/u%���!�b�)����=������:�F���YO��9~:��� !{L�$��O����Wڨ�F��v5��'p�a��;�m�!�
z^�"PH�G}������k5�U�FU��[�%�8�H����o�2��8�uиa-��f�.*	u����X��j�]q��7С�!�,���η�!�=}�����2����qK5���6���;�;���d�: ǝ����:��/s�en��u]���S1�F�Ě�b0p�Y�R�e
�/H)! 6�L�%L#�ч[d81p�[��~i��@��h��)�x�M�~��}t��V/J��eS���lޔ�p�����DT��"�Y��$��2dٗ�l��׎��LT�e�g�H�_�����a큏��I��$�?Y�� �Q"����HȍJ�F���QɅ������,$��򇕑��Ɇ�Z��kl�>��HUyW�Ң/�:4��&L<�������6&:���<&�<B�;����P���Ϩ�B_li��E�K:*t6��e��n����8�f8�b��Í=��j���4�^$]�����	;�=oL� rp?��L]q��L�<
��;k�j�=�p6dk��{�2�gS1�����>Nr��7�#��ןBR&��Rm��tc`<���Ȕ/4C�U��"���X&J�O������o�U��;���]��%�;�r�!�YC�/�U�H#n�'�+W�k�j	�'lO���1)(㽸���<cFZ#�!���lϔ:�F���cJ�PqE�:✯@B�man��R�+�"�E���9�/�0؆��� [��l��w��R×����:������ ف�s���m� ؑ�����0�H Y�h�!k	���*w|Qу���K҉��f�t�﮿�@)8��q��+�r��j	���Ie��)�ۡ�LX>up�ك�xC���q����k:��bZ'��p�Ƌ�A �D_������y��k;�|�f�h.�9��6.�s���zl�p{�1�GR-���v��h�H4����ґ&��o� �����2��0u��6�rHI�Q[og�*6,N�Q 4�$K�x�&���;(_@-T��ӎ�Oy�{9��h
� �)s'�NR}M�jiCxC���G�R$�pe7�G�e`ŉ��B	{z:�q@T?,�58�;�U K�R�$fd��Ԯ&4�ǉ����p��#�f���(ӷthA���[���-W��p����j�� ���0b���+��B<9�D e�;MMdL|Z�໽(��-h�x�H��^�j��2���>#4/��u>�����R�/����=N''%D<A��pM^���z �`n����o���ete��4����DRX_�v6�é�IJ�����ƳnC�_�#Ƞ��M�7
Oړ�Z�f%�3����5��nӰ��rk����,Ɩ<+4�? s_�C����%����+�y��P� �޿~�V��S�N}�̩
Y��S�RQBNÅQ�>�����h���g�d���D�Z�� ��X��U�D9 E�j���r���	��!fA	)�������Zqwh�n3�ސe�jû����G�ztp�CLA���r;�ѳ���6��<P$�9h�L��[��/��o���fj�� ��ɻ��#q$j���2Dv�Ԕ�
�O��<]��}�s����օ��T�����mD+�lha
���n�S-iUuzOjK:$��B�B����>��8��%���PZUI��绛i7����i��\+|����1���^����q�<����������x�͛J��
�������+u���p�� �V�T�SBCu�x4U�/U���|��5aF�xw_��;��=Q���f!T<����%o@fU�+��~ ,�2������w�L|����{��0����/Y͚pjܫ6�+��c�&���=2<&Z� ��� >8Х�sa��3~��7}�pV��&��m�g�^�-KG鐱������,(W�d�f����n�������$!�SF!��hNڽb��t�72М��p<��[L�����ca;O'�S]�Z��$Zi���:ӇϽmv�M�}�,/`�|̠.�@�n�U~�����h���[.�}���>��M;!��ܪ�sQ�i�����P�?u���Ӿ�̴��������:vE���z���͌UU5���GN���l���;`"���Hٟ6���űY8:�wA���]'�Z�����o*S�i@�vv�ȎԬ�_��G����D-��)���R.�3���e�����X���l�Ӗ4�\QWʁKK�Gv��)sR����Г�)�{Y�K�~ӊaշ��=�n�σajJ]���k-��&Q��H6ĩ�ݴ���5<N�lA��OH�6��kJ�]c�W�@��x����H�f�'R�ǖ�9�!:�0�o�MN���$���``�@�D�ξ
���T�y�ogϝ,x�q�d�$Md��w[M� cL�NO�g�(:�唛���L��13��,_	���Z�-l�����@2\��p�&�+�&�2u�J_��u6��9\۽�u�|]Ľ'6�H-�E��&�mf��y�:� ���z�,g�se� {��
�.f\؎MD&{��߇٬	�M�X�Q=U�Ho���.Ąͻ�
	���s;�nB�?a�L��5�����4����/>�K�7��}�������a]T�_�+���5�)qB#�w=��?�-~3�k������5iz�*Бj��fVc~�bI�X\����2��&a_�Eq�er�d�Gͮ����=j��r{+�'��<��{�n�з:��7�6T��i�9��L��Y(GTw��8���E�i�q��i�'2kKLV����������+sP=5�M����.�M�Oږ�yKQxJ�P*b��(��qR�׈�2�Oe��pe�CM�r��fx�֨��N���@������2�7u�%o������=`���$6���"��}� JHFҲ0}j��6L��(�n��S�`u���8���
�M���@�(�4.G u�
��)�+b���b��j^���I��)�X���.��i�FD7]Fڝ�X'n�2�!�d��/���	�N��d��XD�3��l!׾�ۻ�m��Ś � "^�9�5N«���C�xVט�y� ��o¤##�b��Ò��8|�À�!��m��rq�vW��g�{�
j��=Ӱ��uk�@o����[k v�r����5���9h��>�4�����z�#>�S�8�3|��G2Q���A)y
&�!Α���T~���o�aC�\MH,�]��Oߡ88y�������`uL��bAw���sY�����9���ԝ�2���od��^~�"j˖��9`m�(7c���t�/��:��tbl�/eU\,��N��Z}��y�R$z���ג��Pi^��U�禤I)w#�˽�!�[�Vh	�Z%=^i;�D6�d����e�Wr��VQ�R=?���]�M^kr�='�	�<븡�Jcm�r;P?ry@�	/bB�vo)����"!�0�t8�=l��gaS���Y`���NLT6�n9�j��Cb5��@VU���zA�� �){�J��u� �Մ�'�
�%��p��@I���1{�*x�J��6�Jɟ��>�c�o*w���S 	Ӥ���B�K�Y<�|�fN�D�����0��Ǉ����۫w`sXFy�tӈ��)��5ښ�
XJ��*zۖ�%}%���{��UB#��m�[�s�O����)��keDڴ���B����ה{E%g`h�oڀ?x� Q�^C��ȿ4&���0�k3�ةxB��&+mN���DCs�+!��G�մT|X����.�ڞL>8*F��|�?#���q��G!2m�����,_T���b��SjtaP`������^�ʛ��R
7����h�
�%~��0:�g�Z���ӷ�l� �/�W���&�i�d�;��Z�֣��V'�G�7��_Ϟy	�L����\��w�ӱK}#�)��5@C�#�3;ycT�o�����_�:ё71��#F���+
���B>�tON�������M-m8�Jk�=7f�g�`?���TX�Og�d:O�ߥ
\3��\�6V�+�z��{irn��"��ʞc��R��v�y����`r����K�4p��yQ��Z���Qȳ�C����HXL���t­�~��T��J�~�i�l�t�h�N�r�jo�����`z���
�k�Ȧ�B�QN���-5��*N���7��Ve���*&k�	iᰲ�2�Rg�`�M�U5yr&�����j��a<\վ��o���p��z_�������s䶻�@Q�]��x��c2r�~+Z*��k�Hl�2�]0ji�4S���{v4+b��Ն�W_QF*v�Eބ�� �����Ya�O�%���w�7���u�cW����:�������j��]J>�,?�D�j�2]�5��l�J��qx�qz�@���C��=���H�>��x�~��Po �:��Vf�4Y���gz�ܦ^�kK�Jy�!l�d:� ���A �x`gUMRYPhp������t���A�nTN�~1�lb���n����I��� ���h"�â1�n-� ƽ��d�-ݡg{�N/+�JV��)���U�kgz��a	k=ˣ���gV��!�M��	G��݃�D���� '�/��$Jx�b�T!�gL��mz�qÑ;�u{���h�����  ��	CgH��_�5V�O��-H�U���0ғ��TDU��8� m;�L�U)#�|��rimRî�S��)gn~��81�t
'm�XV(6VV�OF9H�n��=�M���v�����;'�i�oV�Y{�2�rx������`c�pG�����^��K��+�e:[;n�T@����n�T��	���I�&3��9�QeGQ�j+7�Y��<�u�fR�Ǧ����d�	�J+�W��j��S��	���z4T:�3����ۇ3 19t=�쫩X��Q�@�f,���2�f�7�KB�"|7
�H0���@��w%z�w+ZԷ'��]=Aw��Y�0+�m}n������JK&Hi3(hEd�Hp�>��#���Ѧ��"-�F��5��!��
g�y&��A�:;���|��������UE��g~�g^l{����9�����Y�b6��f-��c-K��=?:��Z(ͦ`�kLs��/���1�q�/p�6�;��8��=��ڃ�!4����Y�_,2ȵ�a��`��]�A��>e���lj{S��a��CG�����@uv�������@ɷ�D�e".�Hp!���K����NI�;~�pg�A�jA8�a�28Y@�ޅ[�"����rF/C�:��nPg�)*'���ΛVY�+ʄ2L9M�����<�9a�3���Ϊ�uʧ�
Jѧ>}�g)�:i���v9j�F�'�w�^��;��q�(N3��Uk���
����-Җv^�f�0`Mw�
W�#�jBY8}U0.�΅�p�9�#�xJG2R{gx�i^o�Mp�s�Ag�Уw�cq0h�{�f��5Nn��A�,�:2�C�&v��n*H�I�o�����qU�,O Sc�d��6��&O�#@�.��䨝�~�������Jܛ
��k31f�!��%B�y�����TVQ�8Dǝ����y'3ݪ�OP���1��ĬQ�ݼ8&��Ғo�蠂����}-.�_}����yk�؍b�bI5l�bG�̙p����t��?��%,a��6Jo���yN�8��t����� E��1:�Y1�'��������L*�J����δ͝��>&y�.��mF��o%�����O��)�]�I��G��?�3��iuI�Rk�(���+ez�W�AN��\U9e���0]V��e�ɚhS��W ��̊�S�|����3�{�\�����L�r�Ɍ��i��>l�qwY��Z��u��S�A�%i� 4r�9h��|Qnn�I!��v4�2��q�����Jp}-�0��K����%�}�y�Y6�+�p�6��@�3�3�K�n([V�`��)�
�t$L�U�+��#��sܧ\���fm���7�e+?{O��&~�Rö?�E��?��8��3�?���5���|4Um���/�6��o����fR}e�[_lc+��f�C|�����Q�>���]��+�'��Χ��DH��� i�h�@�����#$�I��o �j�����Fm�4�)��x��f$���h��=�;e��z��Y�U������ �v�B�-Y"/���b�a`�{=��8���"���_K�=�,W�`�AKq�Zez���\�t��r�>2w&����XT�S�~��^%\��CWC:�u�Pj��3؎*�O�c҉Li�"����PY�h�hق��zF)x?s덷,qʳc���A^p���2P/e��{�C{���"!{@�a��H	���6�-8b�Hx���u�#��yՍ>K��՚%�?�_y�;Ej���W��7�������e�]�8S�0���
&{�Q���[�4͚��L�*N鎘��]?/�\�)��|(�%��$H[�U�ꀷ��~�u�NE����X7 �h�w�+>1*����DE�	�#*��p�WU��U�*i�#g}�"Ȃ��ދ&+���l��\چ�g�~��'Xg���7�{��j��K<;I >|�KR�n��K�6�M���t;㙘������>�1�@{�-a��r����Zc3����!�+lT{�N�$RǤmѢ�ddD��y�'�'������Dl?2�e�H�s��'0{< W���8��d���[��.˪���;t�zˤ8�s����t*K��]v�d���&dbd*��4��坠?^%�U��Ԉ��M�'j�Aoܫ���
R�Do�sA�!�&*�?Q�ؙ	ތb���b�t!c.��jx{:w�<)�k�uj�k�&�����R2S���7�i*�N6K�ٙ�Mn�����X��s� $��%z��}�D�S�Y0j3�%.��8o������Y�
��R�zn�@��:�J�"��'˴�!����"���D��
��ӽјyv�G�z���i7J��	�A��)(|���X�Avw������b� ��n������+h�P����J�L�J�N:Y�c$*�)W����0Y��I.;]�&��k_��p��5:=�>��1�tv!�:���T���C�s�����=��@��"y�����x}�
r�� 0@�[�_�1����$x���b
��SKF��*!-�G'�: B ���9|m�L�f��'��6���S@e��Хjƾv��|��A�/�L�n@�M������
�#IYC����11Xs�ob�=#�}̫��PJb#|��m0�g8�m�����&�¥�:�T��`���T����̀AiGB�?φ�O��D� ���۸�7cS���F�\J�}��*�"`ę�;��K����������x��������� ?5��-��$�;�O�Ƴ9y`��'��cv�17�)�Z�ջ��8'���F��2Ż\�\�q����:"�z_�������&��/������J�M�'�o�ċ �ԡi������(��������L<NFa���{M�j��X1��<�1;�Y%.9���=U���j��`ڮ���} !�j��v$��p���:h�%l�nY�]@���C������cx^ӏ܂��W%U��)�6��䭦���e��2�$[�K�s�Q�����c����A3�{��l�C��%=9ЬV�@�>YW���a<�-!��� 
�He1��犹��&j=M�:�=�P����Yo^� #{"��q����~�o���Ō�~V_����X�j���tl�/�&)Î��&{q��Ϋ�fo�E�a���t�t,tJ�ae���v`��\"�X4�N�w1��C���cR1-�.24�^��ȕ�kr�������˂փ�Z���?�d����
�����-��}����L��.�i��5n�X����`�{��CU\vW0f%)E͛�e �z�=�̙���=M�[;OF*>q�<���a�2��3
�g{^8Ѱ�v�6�� �d+�~��a�	�����8�!J�����W ���v�Z����NJ��-�h���o��z0[�n�A����Y�hYYh�. ϵ�>����2N�̯�1���zoj!B��3�2^\?2�%��ש����.�r���6f]>�~[�+�XBh`��t*��X�W���O�J�A��-���\!1Y�!aM/�'��ύ���V6�����H��`CO�v�)N��]�9úڙF������<�� pz��p�&����Ƃ����%�/Z�:B�5�W�Ғ,Y2�cg&1��9f���=�O�`��5�I��W˒Wy�_`���s��w�(�F[�~)��8(��;:a��������G�Q*R�t@IlY�8�n(���Ơ����6E����ʑ��]����n�����W0�
h�H�P던ٮ/�+t����]D��;%�.�Z��D�������jt�6^��;T�[���2�׶[����5k�kUŨ>*�b'�)t���چ����ai��n��(�k	��q 	�X��!����W7_�ܜa��<6"3"���3��F7��T�Tn�Ak��;�	�'Vv��/pXs�w�ȫr��p�:m��k�A	+��9���.,L�ݲ������\�[��v2Lq�ם2�>cG[z��)�mo�p�2�Oz�������k��exr�aW���)�*`�/�<�{��HLL��i�V� x75���3u������0P�4+U�L�-��<��o�?3�L`��������S����%`��	����.����	�ap���r:�u��8n22��LĢ����� �3���
6�"z����7������:'=ԟ,�ήDȽ=�N�@5=��s�>�Y��'�I{�,�f6+t�+[o�<�)��Ѣ��ݥj��@v��d��W�~O!�ݧʖvb��V_�Zo�<D��� ��V	��z�\���
J�lS
=�?Q3��Ь!�B&G���)oGv#M��ahhz�]5b��l�֋Y�2W\r���|�����"�/c0㣟��I-�����5���O�݆��?#�!�I4Cqdx�}f�j�z�O%L�j]���"	Sǝ���!��'��U�&�J���4���pqU<w��2�{�2
k 6\	��[��̪��BKॹ�;��,�s��r�]n���T�����`{����j����b�*�ʡ=�l��&I��5�%���Á����-i��|��^H�`(�=:v���]�`'Tw�$?�@�oL?[3��49����D�C�dU��yō?�Xn����l�9I�u�6�Җ.O8�$���e)	�\�@�o� \w{���f�I
>�����X��OA��gm�X�͍9Ζ�3��:\f�.fgҿ�����`B=C1\�&��ݏV�$���"E��"�o� 8�"�����tA��#if�>[# ���׆��}_�:��NM��8c�'��L��I���u�:��?�cu��)��T?�� ����Nd{��t��;e�������	1�t�s��+�-��������������78�,⼕�Jzb"���6ۏ�۪�
������k���=-\۴]����B䏷ѭ����l#+��@�P`&�䴇X�z�?x�4�_���V��h�&�s���}�X@ʚ/SKTw�{���Z��D�L�Jh���է-ȃ[&��:L�Nˑ�O|���-���4
4�&#��n��Z\}N�Z@�y�u�3S�����'�;=CQ�(˻��ҥZ�/���m�[�b��k��������8b�G����;r�Wj�x�ᗝ�͡_̢pxR8����̤2j[9�dC1�vۡ�mt��sj�4����O��3��&ӱbko��y<�H0x7x�K6=首B�\{˶��d�q+����V
�`(�o��~�
l�U3���l`[�O�;�������>L�,�7n����{���%�{6�C���VJHD��?��W�v��R���3�N�:ĭ1W��y脏'\9��t��y]�ZR��h6T���]�z��dqg{`0CX�_��X�eĤ�Fh|yU�T,{+��`��ٿ���F�^��f�����{��A��C�q��;P@{	��SMF6��m�jD.�r,Q��O��}��4S�b	bXHhx�?�aB��9�N�:C�/|��/��4��d0�{_�'��K���fO�r�V����gF�s0{�'��Yl.^��ؚ�,; q�~%74Y��F�*�����:5.-Ѥ�s����s|��?ް��
0�z��\�~��bJ��G��ՠ{���*��v�j�/����o�~'-��]�1�/�����1���N����5�9`ִ�Q���~R�ڃbؖ�%/�o��� ���h�0B#ɇ֞F�ݎe�ޒ˿8�<�*u�8(�/;!li(@�����4�s��w�R�1�*AϰgNE�}��	<��
es�y��=�q�_�8�ݗ901�.$i�7"}V��0��2�x��BKY��g�_������Ƃ�n�{7v<���?!Ď�f��D�B��7ό�S�@2�/�Y=��m�C�G�7_��3f�|�şu|��~�s��<sW\v�&��(�$�����7�ߥm��)���%%F��)�쵌{)�-�~'�{���=��r{�=]��"�G�D�c=������3!�cv���ps�*���93?-�'o��a)��r����{����p�86[˵��[b�6�q����#��t���Ӽ����2�Y��'�i����Ҿ1�t6
HM]����5O��en�Sld��b+k18B5YA7�k!���,:*��W�ĥ��ڽ垈D���!6��>�)�|��}U�B7�k�=v�.A�A��lC��p��� ��&���N͘��%�^������-�A����[�3�_��+�h��D}�ʽ
����w�ఊ��]�F�Q��"��Ho�j�8M���wv9۰�ٝ" �ꂢq�aҡ�~�RN�ߥ��*F���O��P���`|�y4
�����E9)��[i��A2$���ۗ[�Uyp���Qb�̬[`c�/�d��YOƑts{�l�7��y���nH4>�Ҽs��%�+.F�R��x���nJ!���܆���&XSB����Z���vO�M5@�rkȦc�f)��ft+D���������aŮ��x��C�Ql��ˬ���l��M���,��"z�~*r�@
S-�(�Xt$.O�������_T
v�
�E]0ʪ��b�sN��ދ�p��`4)�r������Rv�y'N������HVzV�؆�C�o�C���9�{��=?$����` �����ۅiξ���F��l��J�jn3@��o��4���G]Ɨ��D�:J���J��9�Wߒ�?�p�&Ӭ���w��HT�Qi%W]��8���$ߦxY��S`��$��k@�8:����ހZm�i�t�+F0�eD�!���+�ަbBXj?n��.vrՎtF/��u<t�6��0�Ap�%����sզ�����]G�oU[���������%h]F�]1���~��I7鲺eOR1d�ψqP*�٥�4���w"����aV�Y���n6�~�{ĥ��_$oQ$�o��,f
g�jX��3#+м���p���>P��#Dv�[ᕈ�7/�$dً�OR(�/T�	���=�:h��Y�\�d�\�1"G����G�������.�#$5G���e��ܕ��A38�䵙����Z�5��xQ�k��1S�
�I��xf{0m��M�bW���
�����5�̽�w�����BUn��%��ԭ�����uߠ�;��	���U�o1�^��+O,"���QW���6���~5��}Y�������2������D�{L㾃IS�����?O?�9>.����_}������OJ�=��u?^��i�3��Hl�q���ɻ�L�
��qו�O��FR_q���Xt{�Z�\�?���<DL5�u�3�YP���s�x�o��L}���ʽ�<D@���S�r����ؿ�f`�;J�e�i�
�?e/n�.$t�Vbq5Y^�g�C�շ��O:X&���з��}����"6I�=��T6�w�C�KD@�ҷ�RYN�(%&[.�>L�����uB4KD#1H��?�*x2h�5��7�5KH"�g�ʅ���*l�|�\�
��)L}�"����%[Z��I��`���ց�����o�;Ța�_d��h�x�6��N�o��1g��:;���of��'�`! l/R�ĒA���9y�ĒK������Bĉ�s���hd��Ա��B@(R�s���T�N	�
.t �c@'2���;�fd�oE ��Dc���'L�D)p�X��]�����O�N��Ab Ckyo<h�,C�ݦ#�
ñ$���
'�T��X�&}aCOQQ�I����6��~~{8�T�[i��D>'9Y�J��[���wgμ�j�����v�,V�t�f��5O��]�L�hA�������tZ��j%�����-�U�Ċ�O?�X���q�/�����{�]j9X�p!+zg�Ej&��2���d���u����-[��m��z<%,�6݋[ԬY�W�*F��I�z������Csu,J�ɑ��yW���^�gBz�n�� �D���{��!������ATT	�R:��Hw7H7C�
R�Jw]J���!9t�{����>�~Թ��}�^{�}�=7~�	�j�oC3f�i81 �H���W�#��cV���7��?�!v�ŧ�=J4N�VOh{���	��DjT�N���Rd���b$���J�J=�XC��I��=�G�X�d�r�:EL�& ��$)����,�*A�k��6�����/M��]4� �yuǀ��#�5Rt�CiE�Ѓ�U�6��i>-?o�m:�!tU_���A�=N�5��(�ME��!Uh�A6�]�[���J���ƹC�X����^5��Ĳ��-� z�3�z?��T��8�c-w��E�����ط*�&S��R�������S:��_ ���ƴ��+���؂'pU�`D��p@��hקּ[!{�p��"tu��f�MT�-��D�9������t顸�o�����Nge�飯�e���zrݡq��A4/�1ʣ0���p5��t���G�8��Dȶ���L��u���X�8�ẽ���%j{q� :���l&�.l,�<5ta{���$˟�{����5@l�ʪ����{��hX���Jo#"XA}kh6l�L��q5�tn���s����*%���{0�u �����k^+2����M�R"w�*/M�$��:����ޓ������[���*���=��!��� �"�Nʴ;AJ�2cǋ�LG���웗�xth�AOmΙ�o�K@�e�k��IZ9�-	��|�)t���H�I���.�����θ�\�{I�8�J_��5J�����ا�g��G�w���I|�5:M���)��Aj�ġX�z�3�c�[��+nƲ�ܩ�k��R�N��a�r�HrS ś-%t����.c�
w]�`�G���Ӡ�b�i����&��0��a��\�U��� �V��K5�3 Oj<���=���Ņ��tm�g�܀�ȣz�����s�_�,����*"����d�/X3!#�<-׼&���m��� 88����VMJ5,վ�`�����em�����;���z�~;�z�$k݉��;/!�����]T��TI��%����&�\�ڢ�����SCbp�(v@�l����:o�͟�V�I�u����]л�����!����?�a�<�'��p����ޱv{g�⵵2dM!f��� ks��6�t^��^U�)�����4bg���>���&���w�ݣ-(�q�m�:`C'�<�t1t�9�-O���M�I�AX!VS-,��r^q��RzwO��x����1
Թ
�ߕ��%�T���/�<R�?|�H����o�q!2������9P��T:YQ^;s���/�Ї^���Hrx�ݿ��.� 9$P�
gp���T�]�P��H
�,6f�����i�UH��he:͂tBhe�3NCZ�I3(-�:24���!:�QD��M"�xԥ�^/.�6�LT�&8)Q�+6y����J��o/ �'��>g�jd*d;���y��*[�h�(�z`n6�{[�P�J�'�ښ�V�|��!��������(e��eҶ(���r����o�Az��q�+�]w�Gu/��x@���T��B��5(�g4����ᦦt�׼������s�4( ��U�W�P���(���F��f(���?Z����b�"y�\ƨ��E���Q���Jd�V����k��]��� �?��>bX����le;fM���̥�G:�O��.��rH`b�s���%t����5W���r#�_N6?2U�`G=*�8���,����B�H}�Lb�.�Π��~i�O,7h�`)��o�o���^��8$H{�q��a�4.���;,QҾY�vl��ŻJj��J>M���^��2+R��c�>�B�E�0SA�2V�~�΄q[�@�l�TJ�k�����*o΂w��4i��
w��9�.�!Ζ���ܵ�	?Giv��o�&��F��Z@7�	��&8�l�c\T�+�?��������L�"�X������23:����m3J^���6��\�s�%X�Q��޸/v����ib�;n� RHu'uµ�r~�r���Ͼ�-�}�L⌲K�{Wm��0�/�ڃ�V�j�(�o��w�=}��=�o���e�Vn){�Jx� H�=�8"J]��՚'�v-�����l��r7%ݎ��5���P���W�����6�����2Z<��	��w���L�?�+�	��_=r��L=���@[-m�Ŗ���Mo���_�S��Oᕭ�A�Qu�t����K���z�>�ѵ��y_o�bR62�������%�xj.��Q���a���eB�민�]�����^�kMoן�/���-�9��:�侮=7<�J&��OY�0��-���/���-�@(��m�B�ᣝj1�fk�=������s^LT�o�`�H�A!���)��	����Wo�+����)����jI_���tR�7�Y:=h �`���U�=���'�6/]�-�Sd_���r�#���H��<5b��W��R����C�^&�~-�p1f�o��������?�`0g��?�<�����$�Q���6��؞X9I�������2_��	��0�dD֘�]���7�D�%X�/5�5ܧ
��ރ�;��D,�K�w]d��c�-0��9Gm��H���݋�ͭ3D�-z��f�����xy���_�*��E��80Z�V�e�ܑ��1�-�6C��'�����J��?��\3�f/:���%D�^\>ޏ��#���)�����?��`�e�Ѹge~�ypt�3�6G�1k��

ñ}9�o��4ǰ�hP����`��p�$	K�S���*���ڛ����b�~>��(\u�!²�QMB%��<L���:H�>��h�~�(:��N��-���M�x� I��|�g����.�j�,,�w��;��ɾ@��]�=�#ԥ\�y�v4+�b7ER�˲jaڲ�Z>�y[�Y�n������]Mu�U;H��$��P�#T+�O�˱Y��}ek�(��%R�O~��k6vڛ\�z���Q� ��>�f0�Mݟֿ��ٔ���M+��d��W�~>�����~s��'q�'��V� ]��;�9y6��7Θ��6�9�.	~Lr���Atu�_����P_����� v�.<�E�Ǵ��������ƕ5��4�]4�y�����+�ɖv�QUɣb�g����H�qh�!mãp�;8�|捔W�RK�#�^����; ,��<����n1���-�����6&�z���۬X!�Ş6�>��A�r,���x��7h߾�{��{;QKA~��}R�Ӣ�}}�7d�~B��� }���ϣg��:A7�{p�������������w�y����M��
�ʎG�꺣��!�Ş6$��6�5:�DV�	���5����^��O��R4�_r���m �x���]� �����y�������:n��	U��j͒ʖn�'�͖�)0}Fq�U�I��\jBf���#]B�G?�t�63���{ϼMg$Ĳ?"�ر�&V�# S">-`GX9�\���f+M��9�+�_� ��4p�PňPw�@�K��b�|�Z)�ƅ����a:��	rbӯY��ո����4(K��:�z&��u���ݟ�Y�J�iy�ۯ�Qc��;��#�XaH3��ł%��zu�(�{f�l���ˑ`�׍֚�`tٍ2 ��>Xߵ�_��@��׺�j����肥�<@� �t�&ߙ֒I���Uͤ@�]�μ�p����L�yy�D��f���I�e���c��R:e���4j�Wia��S��ԵV^o:�۳u5H�|�[�,��,���-s���Ȭ~���~�E	���
Td�MLcj����S�|���i�o�C��7����V���}���}��p�X����E"f��O��~��������e6xA(}�¶@Y������XI�/-?Շ�.?�f"~)(׿�V���8}\��PU�(E��eǠ5>�38<��I����
���[�5m�Oט�g]n�<6o8�oq����]t����%y��D�(J8�%�{],�X�u-%s�I��A�����2Y'�/74���C���(?��t��I&>���2-�ĩj��{E�{L���<o��菙WMx��{��e��S������=9ՂX̏X!K���Z�1��Fqa��ه%}�h�� )�=�7��d疏�*)�T�]\�GQ+j��cQ2l�>x9d��T/%܁��lձ�����o䷘�E������s���Y�(�ò��l��X|ak/^�)��B͍����an����!�Z�>h@��dw��F^#�+�~�����\�n����o��g�Gٺ�$'9��K0A��t�� ��ujVhPns��py[ӌv�9�p�<�W�:�3~�����C=^�ogk�"�� ��I�C�H��U�n�QA��j!t�H�Ǣ0=G��x�O��'<`����d��'"5(T�6���Kn�5�J4��t��^�7[������.���
P0�E�ﯤY�?.^����7O1��t�*���a/�1@�j�f�hԚx'�Fg����a �A�&�,�7�r��"9����?����I�tH���H�TX��d�w�M���G+���҇^n�ALbȶl�V=m!�;�AƢ������>{k�H��<(�e�߳��G���f�j���k�\�aU�xaؑ�j�$!��n�a�oĩ�|ޙ��7(/1P`�#�	^p䏄<��'�͉���ﴔ:�Y�>(Λ}�VXUc�JȎ���g5��m���>	u�;3�/������I�jf�xؐ�l�L�)��F+��O�x���y�|J+��%)�(���G��7��)�K4G�*��lͳ�p��g߆�ɛ	��w�x-76轷BTr4n[#��M����PF=�b�������@_����@}������iH�M6�d��U�P5cɓ1+# �J�:T��o����v�k�����oWwj��!TǊ%R�1K�m�{�񝻒~3e�]���Gc�~�k^)]70�~�d�Ԝ"\Q��u�3 P�+��k�o�/|p}�:ݝ�l8����ک7��a4�Ԑ#��_����`rOfN�;p;�A�R�觔	w�qt��ʽw���� ���ͣ�/M����	K�����V?{D���&	Pa�����W�஀l��`^��E��G՛]�Mp�!_v_E�Z�����_$Y�e�L,X���D�RT������Ь���2���O?��Q���^�:hɣ�RAGq�gq���[ET��Z*�a���O�g���� ��Ǫe�~��Meu#8�~�����f+Y\iH��m�,��d8H��:�D>b���X���UHQ���޻vX��QV� C���w}�xD�b�%�n<��DJ�PYd��0<�g�J��K�C�oA�����D�3n�C8�����x �|f�qE��SUr�% �N�{�1`V�W�]~�%@^�F7l8�IR;bV���l�v��~����wv�����6'�Jߎ��>�{��^܅�$E�7H��ͣ4L�C����1�&&/Z�������/�`^֭mC��;�t<~kH=B�۝���;�{k{ё��@{��*L0��'�uw�k��{����º}*<���4���p@ZhR[M�U	���L��	
e��j�����$����4ɜ���;��������*5f�煫b��ªx�G/MƊ?ho���0� w�;�_�&��Y��7�jP��Zm��e�D��,��G�Ga]���в��b,��y	�U���ü����%}l�I}MA���~0�=�	S[)L(�z9�wjc�6 ��}��'�*f��P5�.Rظ�dvM<~V�PiP~%!M_m�w�X1���|���W_��	��D�<{~hG\�#��m%�Pnm�!rl6���dƊ�ؓ�֞ow�zVYa�A���ث���D�V"���d�H�OGq�G�a-����F�Lڠǫ����r���]�����7H�*��f�w�F���+���"������n�W)Qm?�a�{Ǽ�B�֜�[w���),\��+��"vO��c#�Q�{�b��"����jl����;����������iI�9_G�X��K�Bgtt�ݡ�yYUGe,��|.,n��֢��
g����r�ܜr��r�^+eԓ���;�c��T=�.�dR.����zK箕���v���竄U	S�N��4������2m��S��N��׃��-x�=X���_ ��h��s��� Ds=�7E\k�d�9߭\���# u�le>�͕�ſv�*w̋Ö"V2�$l5��^�^�Sgl�[�s��N�h�R��tn3��h&?�����>��o=a�.�^��\�f��ż��ݨ���q����D�9��;c�F'�t��Fv�qa?.�+����j�D=���is�����UZw��n~�i�PxE��gz`��;nU3|y��$�����E����=����jʄ��t�k�|$X�e8�c%#�X�����Ht�G�ol�@դL�Q�
%*)C������Q����+�`�pKT/r�b�������bP����3�-���/ZO	�@-P�->i�Ns�Z(}
�?���zb��Ј����0rP�.V�ro���*��z(������+I�xJ^������>���0�[Y�^��=�����_3x�Di����������T��q!�|�J;�]dY~eg����)�i��QO������r%��?�N}��5�GJ!k�FƂ?�Mf8n�`H�j.>XB�����f;Q�� (K}s�YP���]�M�	`/����������w�>��O��'�����mz$�J6�G���k�C�Ϙ��cP����g ���N�^$W��QA�,u�f�����O(}G��&}����v���=?�|��Z�N�W�%�����{��2b O���bc���'Р74DN\4gk0��>����O�Z̭C �� �sd�jP�[�q�CAM�2-�S�9�k��������)�ּ	Z��Y��_�bg؆l������Щ��Ic�%����"�@I,�  ���.m�Ͻ�q�rlAG:M�N`�?#�R4G���CY7�৘���l����:n�0K� BW�^}��'�D���t��spR�0|l=tDXz��Ǳ.��c�>��.�Nl����=f;��v.|0����O��?,�=GM��z�x ����������[^�^f��Bd�)��巉�ER���#�w�.�m_�#sj�a�x����Ve�U��x�x]Ȟ�7�^eװoH��KC{�^�q��v�~��Br���5/���R��%��� �ǹ����W��������cn��}&F�2К�-lʴ�
LN�H,���g>�q��_�
.��oS��
�Ᾱ�ϙ�p��&d��I�^�Soh��Ɵh^LU%��by�:������*��`���j*IS��#-ٴ ��P�h�ʂ7�u�����ok r�i��σG�n?ol��nj���l�γ�/��H;?�U�G���?V.��g��|�j�_:��CҠ aњ#�#��9�
k\�eC_D{��d����,��ok�-��GG�zG^f�����w�1mPe,1L�tK��u��|764�MF���@��OGIe�Wj���3!�0�;�g���}å(m��A�7%���s-*���6~7���%~R�< =T�s�`F�sEgo��_�n����'�ִ�o>%�0�Y��tj,��A�~`зn�TFY\קQW1l�pz�l�4r�"]�/��a�\P�'c�A�fr�OPڂu�'H��.�5{oH�B7���������>���4���C%ƪ�a��@��=�����s�"!J��i*�D����3/�("��)��o`9EF%�m.�m!]`��H��웲[��VO�/P�,���~s��Q[��\��ocߴ������eHO��.|8dA��M���Mu5TG-�]�bmf��>8_Tr�C4c�
Y6.�4yz\�I�Z>~�g&��&�0�k�	�x��M������&'��ٙ(���_���� ;���L�;C�$��������aj荪K�	��m� �N{���O����7�ǣ����/�=���L�FP�J�����.A����R���]�B��j�g�+�#N�����O�fOp���xO�Y������OU�E3Y�!^^���k@���٬�5��}�Rme�\��{z�k�j�$7\��;D���Y~<Ll��{}k�X�p�U�DB�Pwh�ta�u���O�����²�����B3k�$���kȂ[3��`�m�� \`�-Q7HgA�diw{:�GMf`�W��GF�.���
�u%.�R�m	&��T�͠�������� <���[W]l��=8�s	�5<8qt@4U��Y���D���J�����������(��'�&�!BҍM��{��v���f�tb����e
� $}�NL���� �\�����Ypۜ�7�N��r��W@D�+�t$\�OI��;���E���
���	M���lA]�]�\�W����J��}B�p�L�П�>12�c�A���E�8�MT�2$�7(��o
��E��U=���J�$��Z����Q��t��}@���4�ɻ�+�_���6��I�����I��ųDa֒����<q���'�����{c�K��}2���ᡡx�t�M7d?��Y>��%��F�%G	h��kh�(�����T~�4�z��b��)h�_�ߒ�h�Я�q%�=���{���i{�FA�7�"������V�X�s�r/����$;�]��L���}��9�K����Sߋ�qr<�6�mB���ښ,����	��B��NA�������ѣ�|j�s12�]����v��Q�v�{��p�����A��O����������<��,
|720���X*Г�W����ݭ�%�)�����p���f�q/��}��~����9��I�2�е;�)n0)F0U�a�6�)�Ǿ��&�M�.z�lP��Ļ���e�gS O�!`���N\%c�i�+�������;խ_��b;�Z� �L.��\:�����:����ܰx�ӻ�����,#�V�gZ���l���6����c#)��	���`i>;�-\��Y]:%�Z���W9;�ڲAK`��먳Q�#t��9�&<����-�|G8���r��F��o�3bf-��Da�5B�E�K/<>��!���.�������
YG;��F�9Lo���U��X#\n7:"d�����N ���vOs;ȳn�)�w ��]�p��HԢ�p7H.YK���i�83�������H��[��a���5,G [�G�b���y�6[�3y�2�D9��\mU���3i�߮�&����(��w:����,}Vȇ��R��$�O���=̐&��8�NF�����em�-aչ�؅�
�(�*��������P)�+J<�;c#gb��3ЀZ\�G����:�4i���3)�vd��$ �]��'t9pC�X��8{f����~�hR��o~�zǪ'Dѥx��C򌧾�<�I	�0av9eӏ�M)�|ڦ	���޿Ia�����2B�Ρ�C�w�XW�b�����/���=8a�Z�zd�k]�|�_�^��>�|��/
;���F���"c{���^/0@��o����Y�1�1,
M��]�؁Ң�*��+/Ei��8e֬�%�P����ۓ�+���W��GQ���
�{,1���la�k�1K�,LrU�t0�8�����f�~\�Xb9��0���!��$��tM������3�T�Kj���f�o�,&Nm�=�Y;���5I�we~`��1�X�=�ڣ��B�MVK[Y��f�&��U�K��<�<[�ǜ���zK�"1u�s|�͏��,)��o�mt�/����C5��zU6��D]����Ok&��N�_�Ҟ�&�n�i6�71^y�σu{�X�Qh�_�	(6����l����=a�I�Ez=:�����%l�Iͨb)���,v)Ġ?�.ye��,�d�Ɠ��
��-��QoC6cr���(�,)2~t�7s�m�@��0�TڗO��$�z�0�Ӹ=a�˛ȧC0v�^C��	{�2�+.��*?`��+�m��.�E��歚C�����ֲrA\{#��7t�fLct�2�b�җa6d��{_	��ڛT��K3��?S7{�u7o�e�J�~��-��ß����B�\A^��;�E���R����m?�K:�Z�]YT�C�Q�vz��R�x�XjGœM ���n�O�$��u�oW����ĭrl.���/#�����Vo
��x�)�b�V���^���Д5�gN՗�p{pΈ^�F�%����s��Y���|]�建�0�k�+U��eEn�	&��˻.�HjfH]5U��~����^��+���8#�qq`�1v�Ҏ���C[�h�k��q��<q�����Z��,/�K���g~����5ɢ�c���-���bh��3�ԭ��XгK�=�G֞
�1��Z���h��yyy�L��O9����?�פ'$4�5���q|�i<J�亽+pL�9WCm�F)v-^)���`�`��?�^�ag�n���j&E���vvFEQ����M" ���=u,���x�4�ſ:W�ẘV
S�+����U>Z�-���cy<x0λv�y���9�k����xz�V�j'�VV���R�]��}X�à\
��n�a<�=_j��ܞNU��kˣ��Z6�*b����\�{D�p�\'��!��V���*�ESZG1�LP�c�y,��fh�R�AtB�j�t�ʃ.mo�{��Pc.���J��۞>'ӈ(�QV7���;��F�QU��y��-j���m�~PG�|�>n�kn*�e�#fz�4��LE-�(� ���V�/~��?R�(�Ms�K%����e�L��d`w��Z����/���ݗC���G�O�G��d	���j9դ*"�"~S�.���gv�p>��P%��r{Z=��"���l1��e��ֽ�;+�[��}u�ׇ�x̥�*�0lN}<Y�,�t��Lw�[Uəu�K�>�si۷Ծ�^�̻��#�UC
��9y>V�v���)W���B���e
A�q��H�6����?�Lds��"ڐ�v;Y?*��й�=�|y��U��(��Q����o󋨶�a���\6�IP&`R���5/���_�d���oyA�:^ʆn��Y������^�P����|Qji*+�ɟ���L ��L�Hy/K{?@�{��b��s�~E��f��lJ#�7��\��\
�t24�./����qR������m�E�F���-ѫ^��SOMwI�X�-�`щ��<�pW����LA����?��6 05;�1GU��P����
-L�ܾ����14{N��Sk]7,��s�=�;�1S�Of��WW12�˩�P��o���ƆEmJ�G�|�Aڃ�4T�X05���5�C	4k[p����C5�Ч�r��$8J8�~���H�����L����^���j�YܒO���(�]P6�H��=ef~�������"� ���/�^�����pU�'S��|�C��_X��ܷ�_�æά�$9x]�%���vv~.�y;f�f+<�zy�]xP��)�A��l�R�39�%�	:R��<��&-��alGQ���	��ߞ�W">Աh;L��`S�>Ĉ�w$0���j�#�Bѽo 7���Rr�q#�u�V4���ON��[#�PowS��5�������!}c���ӎ�C���iU��Y��HĆ�C}R��P�	7���7�ӕfɈ�l'P�L4��G�l�o���f��J����Q����K�����U��]g~������ψ���y^K���B�w�w)�s��q�k��M�ĩ�L|���{����κ{S?����ԥb�`����|�و	��Z��|t���;0�X󽱝5�?��P��m������4"�^M^�cc`.���=KN��r��W����O��3$e�i���L{��S�}�;����"���ꃮT~m��	uy%@�b�@��KG�'��#���N��m�'�/�b�$���E��5���y��^��i1\�8�)�$y���� ��IZ��/�Co�Y<���`�����6h���������;��q`����'�|����WH���itF�A}�2���F�M�}�Zhz�@H���v�Q#�\��T����ud��\�k&���*V+���.�<�G�n�x�Cb�;��t�6�P�kXW x=�e?V�@ނ�ꍪ���/H>m	���A�#�ݎذ'_����#��~@v�,0r)�}`w�ķ���S���ݼ�P`��f["��d@e>1R�P��h`��emeM�����,�}om�����T��%mE1�Gߔ�9Ʊ�v��ؚܑ�#pߔ '��V��m�l9?�Pk?Z�.D�R�_]���;�$o���h�4��-p��ޒ�V�m��΋�>�۾n�dgU����x��Sh�$�_��șZf3�R�:��C�5�x�	�k:���L1��kv�4���&���ֹ~k��HVz��\S�(���d���idY�e3e�1x�o�iʒ��վ�_H卌�͸�W�1�y�M��9k�$>m����i� �\��5Y��w�]d�e�I6���;0P�?c(�����zR�kӇ����"�r��FҶ��ʿ��a7�9V'�L�;a���?t���(������j����gPVف�W��q�$92�A�	� ��^8]Y=8&E�k�E0��I�p�}��!����RU`����7�����;G�5�L�U�P�k�.g��K�wK�o��8�, ͑�m������ ��Յ��J�#�X:��p� qVS�����s���2����h�H�O�N��ȯ��U�X�*�������>?��D�(҇����ǅ�1��D���pr�>��ŗ��*���mOA2��.Z�К�Cy�ޟEcB49X��(�Z�HZ�fZ�Ju��f���_6�6H�8��dǠ��ɮ�*�x��8�Ã�eo5Y��M�հ T����r,���8��J��AV���ʜ�H�.#m?$�%�~�4��)'�;H]�t'qCMF��a��*�L?�@���o���T�dʅX��a��S�Ĩ�8�}�����!���5��}�!%B��[D1Ι71���N^My�<��U�V����\�qTL�Ov��Z2��7�g��ݍ-��B~���%���R3���+Y�9??��fe<Es3mZ��'
�������6���C��������V�&��gf����Gm�Zd���4!�b�B�]i_�N8���\��$6���� �1�j&���v���Rr+ܠt%�X�W���ͥ�x�zꕱ�,���T[,����d��9�����¸��w���ކ?�y@1N�7��B��J?$L�Nu��F�H*���LA0��a�j(Q+Q��o��� �}���0ƹ�����)���1����Q���k�2l��	KҮ�̄�Ȼ������u�n�����H��z�0�'�f}@�
rA&��"��*�.b=��./�Ŷ*�V��k˵WPa�l�C
�]�KU')U*A��x�+�6�Y�mI���w�]�L�2B�Deި\#�3ɔn��j��~��ӕ����{v~��҆&}`��ּQ)O�������#T1��C
arn���E���}CP�m=�3)>�h��+��{2bZ�R��C����a��Ո:o�m1[�f����M&*%JT�TRn�~t�쾢��be�Wjf�0��.��y;�'n�w��O�E�F|��ld&�Zʘ��m��R6Z	Ǯv0_���Ft׆g	�u�O�%��3*�|�u�B��<P3F/`��;�'��ƾc����e��8e�F�Íd��~e��T���r�Ԙ����{MN%�T��Q�O���F��v��U�D�>��76�8�����$俯Ҁ����Ŀߣu*�I�R���2V�����aa$�l�_W�?Y~�kޤ<�tW�6K&��yHo��;uv�SQ,Ϫ�Ang�X��3�RC��R�G˰�� �ogK,fm���^L��3�J�E�\��0,�w�'
[(�?؛�*3�Zd~ �l\��r�Rvŋ�Rb��×w�w2��P� ,�!�
c�X��/���D�zc��b���ؙ/��YH�47�
Oɘƨt��^�W!\`����hG��x�Y@"w�M6W��k����e_G8��)-��1L/��c���@Pf�<��V�.E���>�p1?��u��gzr�c"HR3ܬ���`\G�IcX`�X�I�Ӱ Tef���<<́%����cc��I���07�p�>�W=d���\����o;
MO��	��^�m+����Ll�������A1 ��B'�9��.K��6����3[�*�%��`��~,L�������K�vVh�IO����hF���W��0BX�f�f��gM�p�R!�e|������`"�n�Fж�wZB5»o}�u{]v��I�Q�7�����2���S���D�s��Gv����ɠB��
��f��H���1Q����WܩN;ʁ�(�\���t]��#�Up0��դ�dp��R��5h_\/S1L#H�{�e�)`�ݣ����#Vu��%R:��F5�>!۾��˩��A]@���Ͱٝ]f��tFｈ�5 �ZI�S�`��>�`�E��U���$�jbK��[����Z;�Dd궷��� 1�P�A��pW6�~o�>�W����XzNd�O���H�r'4���������e��+�FH��@���RDNC����Y�Y�i;���5�*�O�d���9ޕ�g
�Y���e<11&4.��7v�7�j�7��*=�5TAkR�[�8E5���'Lob�����n��v�!��� ��c�lyE�@�l���K	��@���G])7E��>|�e9��4t�n�b�=�=a���U�d=R����Q��qR�U�n'jo�R��C��V��^��*�X3��u�Fu��Ah����#t���T�J>�Q,5{�!�½�*8�%?t��)jlG�J�#K{Gь�]f'�{�����x�I����ޤN.˟��UJ�BĢ��h�~v�Э�a��d3&"
�tP���h�L�u&@xn_tW�>���ȅ�d�;�����K�\�f���Je��ߟ.��)FP�X����'L��4_��Dy@�q�C-��w@]�r�r��2�A��Y" k�;�Xز5���;�⤟�5v�?bQֺN�V���Fz5;/�~���γ0�Y$$����s����׷=����o	$���KZA��5+��p�0MZ��N�;_M�\~w����V㋨K���3��,�vț���9�X �V+yOҬE:�e&?���Σ3ϡ⭹+9U2�U����"| �~t���y(Vl9}��W��b�W�;�\�c�ò��U,�ml�B��"ݺ�AD�j+��1�9������g��+��3�c���l����w�2�/%g��^nG"��!N|{[1om�������A9w+ʒ�T��]���ȯr�9I��~��Xh�{$rtjE5�	�? ��J�H���ņz�$w�g���v�*���L"D�V��;����L��(�M�8�l%�&��W]�A�W�Ki��wK�4e��L�ȿok�V���o�Û�eǙq�q�ȝ�ޕE���N}2�` 5Y�M������}kw��gj�a/��,n"����{����2Kl�͝9��fړ�e�$ᆽ�`;.���iIe)�Y��8��գ ��8X�SK���d�!�@���������~�m�0�@��/���d��y?�8iFF��S\/��}�I��^�ު�"&�OA�&�7�O�*	ZdV��eA��p�6l�^��B��I]��O���O�.}�\O)ܭ�t:��Ô<�-or��K�t�A�Ǌ!��Sj�,�G蔓�����KF=f�顈�oy|?��qx�*[�i&+��(*z�T�u�u�T��O��9hF,�T��g>�۟���]:���V�b�h����_����&��떁3�zPᏍG�	��r�wV�1��Օw�4�:Zs�s�v��H�F�B���?{I�,�����m��]:�O=�����l�����r �񘓧#��'ϝ�cz^��f8�P8^]%*\�~U�Z��]	/���ʯ�cPΆB�U~<���"��\�2���<���+��+�K�bm���=��\x,�3���3-�V�V0��6��A�����n�D����j~;x`%gс�?�HA�d�M�/�o��$��*rEW������c��:C]�5=T����3���3��C�Å#�!��f��]�ۆ��rgu8��}ߌ���~NJp�P�����^��Ma�]�W`M�?���Ҟ~�Rb�^�z��X���/�w����T����l�{X|:�<�����(�Ry�;M����h7�.9+F����>�]�歱|��'*�v��I�����I}����94�3��i�d.v�2
��q���	T4�XUĚ�`�f�����2NL���t>�Qk�t0�B�c[���+-I��W�aP�#K󸕭\_��z�@��-7��D�Ǚ��ȞXv����B���y�[\�eZM՛��H�Y�;㫁k����X��t5�:���i�%�]Tӫ̈́<��rߴ�{�~�
7��Q�7�r�т�w��_�B�JĐ�8w���u��x˩J�s���j�q����+�BM���C�?��*�G����oʛ:"se���\��@��r	�f=���e�ۻ����v�V`DeH�ExK��2@[���K���d���Y.��ڥt��ԲVʝ&�ј���������ڜ�/OƠ c`]nd�x��fޑ�����y�q���]�o���b'"����B��ގ��ld�$�f�$xS��V�zh1W����(aߵ���Rh�F�Z��ZrGWG���)���#�K0��8
�$�6��wEy)��o�k�(y&x�EU����9���uʻv҃�;���տa؇m��n>�T��a D�i�\��(� ��@iW�u����WD�oƼ?;�+6�N��S�F]�nUW����@s�����O]��'� L2ً���ߦ]�g,�8�o5A���$P�T��Ȑ)z9I�8�l����	���|W�Z
쓧=V�1N�bdF�~��	�����79]Y��T���� $6Ɖ>�LE���g�դ/(W���?Vz�,��P~�=�M~�_�;�9*D n��U��#M���PR:u�≥IO]rV���o�<�z[-�\��&Y/45�,��7�/�(�m�k[{y������Y^�SI�׳��	�]"=�C%�M���s�'ٚ�v R�M�Gu�Vrvƃ���2N,h�E��P|F�\A�t�A��E�}���7j_*P�j��z���9lÛ�Q[Y�Q)�މ�����3�Nj�h*_�/�<�K=�l5l�Z$��z��HL����?�ӂ��S���3^
�*w���7Ģ��z���^����.9,�_�j�C����� ��P;�٨�)���Fׄ�r��Lz���O��2�ݗ�I߹3��fU���r�$陫���z�(��{xXVp�`3*QA@W����3��$IR�HN�$I����4��<���a��}���s]��s�=�������nK����f��'a��pF�{ּ�&f���03rx<�u ��`�oԳ�p���O��z�+)*Δ�>x���Ѵ��W�I �X�g1R}=��9zF=Oi��۷|0�f���|@�iD}�u8� g^0�^OS��`8�HJ�	�������pe�?e�P=��ĺ�����o�h%e�2V��7�$�=꬧�ؙ�>�Y�)��y��H|�*ς�Q����#n�s�hjOE�8�s>[���7�8-_VSX�_�u����65U�16��M�6��f�k݋�j�����"Y�ћ2��_r���Z��5��6�h������,��T~���%�n��(a]U�Tja��f�.�η}f�����T?3æ}�'J�t�� �=<ò*O�Ct�u�Ps:���?8Ѿ��^�ޛv��c�c�	���3e/�>�M/̅����ŉ{�rZ�Z=�Q6sm$vc�5�(`m�2P����1�ٱ� �T{+?�rPm�6}i���)�ĥ_�'\�&�rB��#���o�T9����Ci�����ZފcE�dg�W��sU]qL����a�Ms��@�p* ����k�MWUD�$u���<;7;�ժe�;;�g�vДq�)S������1���E�y�|ѥW�,?��x(�Y���[����|�9��d뛞L�u,�4����tʬ[��ð<N�p�(.��
���I��J�Ȩh��_vM{����3=I��sX��T`P	7��Iˎ�͇<�I�E�����}�S�� X�m���ӉN��]ݿ&����_�5ӡ{4:k�����z�x�5�|8M���:�7v�@�d0��V�ڞ6ۭi%b��G$.�-�Y�Э	�v.9����u�vO���*I�\���,mǪ�1�����(��2���&��G���j�~�	�F��|J�M�9�����l��A	��9�'�����w��,RY4��n�{߶-<���G��z���1���nc$r�Tt�	�9��F�V�5㢰5���_����4m���'H�qŠX�^�.�1�z���gK�I�ǡf 8���׮#����<��ư���P���uQ�Ӳ���'sOm�æ��18�e;	����1(����;k쭛1P�m�دmoi�6�E������8�8�(@��6�V*.q��T#�J����Ǹ�6�_����(7�W����))��q/�%��l��B�������|�s�#�ؚj��蟸ab�$�"�)�������t�*�ܣ���6[[^����o*'%o�k/oׯx������#ʞ�$0ks�Ӡ�IB��66�i̥5���?k��T�����sG�vO����N�����(z}A�R��v{C��O�뱾NУ��^V� ����ņ�t�C�(1�(�4WY�<��cW*
�����6�rQ��qZiz��c;�4��
�מ��� ���ԃ�J�ě�K�@�l|��G0
_�,E�������W��0��
���pm�����`܏C�%�u�镠X����Rps�����t��hVn}l�@��Dg��Ci2[�ffP�~���fl�W��ofҴ�]wRP�r=���|��M�b`���2:��X����_�jr5<���閼���;ZcƊN,|�*L��@~�X�0u2>-��$���ϮF%�i�+�T fm��P�Y�=c��]E�ȷuN0��1|I���f��g�����8�"���μ��</)��ួ�>�[�*�A�Ot<����8���MnFj*D���P3�Bo�������s�X��� r�0��}5�ߢ�xՈW�w��#��j����^�(�]a 6��������e�L��]�FB���E�|��oŜ��	����A�Lo���~��o#3|�QN�i���t�)�+�)�3o��xM\�9��[H�ǉ雂h�E�H��+�=��f�8r�N7$�D�E�(�U��S#�Ds��S�Ⱥ�Քva:��d�S^3���we�V��jC�y�T�n�KWPES�H[*Hې�����68Խ*m�un,�\�SZ� �J��}��pIn�P$⪂rN����C�'Q�Ɏj"�s��Ď,���J�<�b�Z?Vn��5qnU�L�Ꮮ}B�l�]Ĵ������q^pĞ�z>Ɂ�3+2N=�D`.\`$���H��Pp6�9�����Rمe�Q�� �v������?L07��J?�o�Z�������:]�-le�~�Ĕ������yw�R��O�X�{V̯��zy�P�!h�Ʌ�K�� o 7�eڳ�Q��Ƭ��>J�O�4�A�����)��S��9X�f�/ F�H�m�
B��c�l�k�[j�j,�?����oZ�}`����,�H�H�T�u�.J=�J����z���8ORc/s-IN�uUKPCG��ȣ,K����l���4sg�,�TÔH6|���a�|�$��?&A�����O0���t���ӯ�d�K�ڠ��B�*%�8Rp8��IW��+���'��c�e��>�����83eB�G��t�'jϫ�C�L�fZA��;�
�f 
m��}�4|��Q�Lz���;Ysց��Nf�y�sTU�b�w�����㒢B�����#���ܭ��;]f~��6a�:�'���F��TT+%�ޭ.�?EGH�{�K"&>��ªs�k�cRk{�ua��i}/ gk?(Q�e�՗��
x"�_(=̟��~3�41;A���@4&��sz!�+��Y�4Ղ9 ]�5�J��<�R0h5��vJݚ�_ϥO��B�b5<�i��sC�ߛ�r���b�=�a��&_�)8�����+���^ �;�Sb�7~(�_ �\
>Q���i� D��Ȓ<�i���X��r`��&P��TR��.�kɛF�^�2'�w�I��	���~�� ��5 KyM>���V=^�j��!��o�.��#��>"w�f����S'ݝ��J��q�ف�^�/�F�n*k����#|��ə�^{���+���~���!�O�˴������fÌ���iBX�vW�
k�W���;d͸���dV�����:ɕ2*;T,�͟Ng��t��G�B.�w	_�:�13-Z�4~�J۷�1��`&w�����(�A\jXsH��!{�(���}�j�A=���0����O{=�~(�{ZN9��{qn��B;�Ij�
K����	Lp� �o!��D��>��� ��N!M���C��ߨ�+�Q��]�p<��yB"�>��ϊ�(����5��Q�aNET�
p�Ǩ�(��>F�ܼ=7��3V&)���.$c�����R�.<CB��@e�Fkܼ���-`k C��1�T�e�q�M ��Ǿ��`��@���bTqތK���&b�>�:���nz�0�
���cx�����̌�(%M0�M*���\��7�~YWB�F[(Gu�K>v|>�S��T�񣅫�	�e�> uG5{�3zޤ�����䤅�H���b���+���g'��7���^>�'��Kb�k�OP��p�1bpb�l�h�ut�A� ���W���&l��=u-�ٙT.+����3���H�6��A�?����7j��a��O��)wH�����v���wH_�s�e�OP�!�=!1�|�T�+��R횒�y.o0�u�#<��9:
H�7�jހ+Z���e/���ũ]bd�����y��t�3�ވqR�y�5�/�)��gD���o �o��o;hy �K�=� /\��4*��<ؚ��=L�Y��=(7� O;@�\[;���@�����Y罭�r$����J�`@�0̺�K� ��9���>(�U?�!1kd8�[AJ�7WL*%X�X��hFp�~~08��}�oY��]y�u,�w�,�P�%��>��ޱW �ǸҬNI�ŠQZY@Smem6�aͦ��>��AӾB�N�8<	��ʂ�V��3��)6��׶�?#R�u�h5-h}O h�_���<^��/�����Nѓ �����=9����_*����i�Ǡ[�����k���^�q�B�z��IH�N�һ.����<��b.{0��Ye����%6;����i��6��'0m{P��L~��V��-'���߂�������I�J--|��9!qb�|`�� 7��6ٵIܽ��Ӥ_3�PB�E��cr};���B��{�w$}�M���rY�o�a#3�UE[)���䀗�t�΄R�ϱ�8'o'iě;��*v�_����+MwR��E��_(��+g�����-X�0� yr���\����{.��x*wt�����}�Ɠ��p~((�xi���ko���[�����S��4)��!�R���|������A���v���c��d�WXb#	P1�� �ԯ��vE���{fv����|K��DQgOh����y�_؁�y�R�E�VK�(�ԧ�J�1���9�w<��CEw�����D
܀V�߹���G�	��7�R�T�W��1����`"%;��2������8f����)�Wl�,V�,Z�ՇOS\���\����;1�
�����z�H֒�al� 򭐲_���H$%�ڮ�T�\���;����bK��`�� B暈��}��`�i�'e֩9#�f�с'���P�q�is�w�y{T�q��TDy�U�|MmajJ��Ѷg?�l�,��}{�w����B�}�:�j�Ԍ��!ץ6T*tʷ�Q������͝�Z�xM�.ׅ�y�~��zsHAU?�o����.g\�Z�V!�֨�p��i� v�'ײ��)���SoCu���9:��Lm=~A�uw�u�d��{��-Z�~���A�y8��¨�O��6Ew��z|у��Xll���g��F~P�oz�۲����b-�x1B��
(eޥ�;oM$�uvv��N_�/��u�	�����.uG�@n=k�ށ�����#��Ϸ���|8Y���Lv@����bgx�ǈ��.�G�.J��gEG�,��#eLz֣��k��!�K�vne��M���z�=�+�G�
hϯ�w��*�Y��9�
q���M����CM����g�W�w����2Þ���)�
Z�@�>nWo=�&����W����	, �'6�γ�f����W�9u�k?��v*�����������/k:��G��K4�JRv	k��W�oAd޾�i1惰�T��:�W��pݔ���F�����;�k<�C=�����-�N��w�Ue����c^sj&+���'i�xQ[j�l� GWZ�A�!�t�`y��K�5�-\�o O���`���@����5��t S3��/�G�In�-��.4>����[tJc������`ס
>]����/����� ߩ���o���k��ϩD�����K�OQ���K��9h8G�|!
�ݹE!���A�ݼ�/�p_㫸��|���*��-ᕺ�/�?���l���<���7@4ε���ޮ������$8	�矙��?O�����y���$��.��9����mJ�jRF�X�<K��ug��V)�[�9@��mFBM�f1���T�Yҝ�s]�^�m�:��6��6�W�#�|��&?�m��d��T��N���fU��rIu�\'dW뾆�WGvZ�g[S+� �)�I�O7^W�};��\���ڭ"K�Y����=�9�I:`��mEv�3��VͻI=I{���6�+��=J�덫�EԎ�,{��'���� m�����?���0�2��{�sA�&��{��oB�P�(ݙ�"��Vŏ=�/�D�U��������� � �b�����cf��d�fc#'��i��F[Bq/�8�-��3��w�QØ�&CǱqF��c�fOO�K}�Ț��V��<����i/o����:���#�>��+���1�xHf� fWܦ^���B�(h�;I[= ��Ag:�*�v�`^j�٪I!f�o���C-s	���[k��|j�,nP8���u}���ǋ)݂Aݗ�m�|����rv�6�G]�(�*Stv�nl_R,/%o@#L�i����A~l6w��V�����}�w�Lx]�&�;�s�A#�MWz"節?W4|��<v}q�կ=��sР���<AY�Jx1g���	h��12��pP�n�u�>$��4��pjG0���K��{�,�w�����R`f�W��A����mom�"D�'0�h>B��A�H/����^�ꀗ���
��**^�5�⼘���DwC���_�ˈ�!��7h�<�(���їV��ѽ���8\�f��JK�޷����g!���y$�-0�O��w�zǇ}@�
b׌/%Ń��8G��x`�W)Il��ՄLG�/�[`��pŁk2t]0�U�*��v�!	�U�U�@8'M=^�(�}~t�]7��_w���`a��b�@�Wz�͞áu{ �Z���h.�� �?��]���oq}f�K&��I]�m�/[ �S;ሧ+WmU�.|���������7g�b͵zR/�MVs ~3:S2���{u�u�$�o�q�t~p� �ӷ"��D�˙/�I-mqʹr���%�Kr`VՔƕ��=��j�xϋ�!;K�;,��������z���F� g�|���T��>	7�ؚA�A�������|�o�'9P���͑��������h^{��D�<mna	R�8�I�I��v��.|4[Y�ѿ�W����Rq
�Ĉ�����{���=�V/��]Y&WAuK�O����k�H���5<�v��{^���@"Ѻ�i�)�(�<���WKC_W�!߻�|��Ǆ�!?�+�hp(��N��1L��b���'/w6F��.��z�nN>�c�DߐR�sn%�`f;��8s�w�c�A\e>�wE�T���J��jSa���͘�:
c�#i�=���݅ �JV�S�l�糘���ͅ7$�_(����Xj�Z�i����@�+
���%f��	�]LJ�X��B��8s��wH�ǝ�;E
�e����թ	f��Y��"��mN��*�,1�[�ت�5`u;�!���R���oqIe+F��ry�Y˞� Hq���������֤�݃hAu�����ހu�&]�Ke�*t�9vs����ā�ͦ���1\SD67�K��;��ѕJ0�53,�5��Z6���7MV2|��&��k�q.�7�f�DAٯ5 ������E�w�[qQ��^$�k�Pׄ�l��W�.m/
�����[M�z`a�������f��Øk��wLf��1��粐&��T���ou��_��7����z�� |�""�O� 
ڰS����v63�[�!�L���-���VQ�%p}H�_��B��i�ƘA?�:����&�?�;+E%e!c0�@2J��NÝ���Wa ��������|�L.���q�%����ދ!����s������ĖnZ���F妘[�͆���tg��V�z��Ns���0���n��n��[F5��?�k{��w`�c0VyP��.ֺ���fpՊ?%}`�Br0�L1|����ݟ���[�^�Nuk���.�Ʀ0@��
zh���m}'9r��c����@��!����ͼ�>MN�X.�������e�8�n8ǭ>Z����%�f��a)�Su��H���S�:-pr�*A�'&�6�r,ÞՖ36��@��%�:K��������I$�;��ZX狂��ފ���a�!�,���k��EH7���������k�W+b���BMf��Ϭ�Xdp��~t��f�`�X�]����4=M��ᗹ�ޏ<<Tv�����z�{�x�{x3 ڗ�8�P��O�~���z����E�\nn	%�YR"��5��"�.���e��F�ma�+�����������k[e��+�2��J�ꦘ���B��4D�(��m�xЇȄ�>c�V�)���ˤJ/Y��`_�e~���t����6��ÃC��.�8�($⩙��Ӟ-�E��;m{�MW�: Mx����a�A�����a��6=��RB�'��z�ft11�_�]Eb���
����Z3!��B�B�K�ކ$(n\"5���:��x�G.Ɵ�`9+�Yi���&fh�*U"�����VF��z� M:j'���%�`���3�B��i���w䶶&P
I�J���[w�Qt���T ��^%K�T?�)��_�%�Zu��Z��X��6�h���k�&�{��Ȥ���ėX�mO��Z s�Lx���Q��ݞ|I���|�����H:���\ϟ����PhO���v�C�\6l��ᶼ�����˶�����1-��: 8�!���th�{�p�������<;�0�:E@���gǩO�-(��("%�S�q�����425~�9Qr��O� `� �֓�k�գ�y��+������g/s�{�!�ۭ\K���G�i��C���U�X�5&���������Te��|6CC�ݵuO�}�׿�|#�we+@���	�e?� ��5ݖqD�%;Xڛow���2!G�(b��)����<d��t��퓐��`�8���Q���0X~Y�� ,�Z���%��T`�e�:�������B�#�z�����>���:
�H�y���+w�)�So��E)����
sTL��͒X���}K�T7�9����_Ր��V�����X��%�8i��/�E��ں=�!q2K���b=D�۴.��a�A"CI���h3���E`�s��%��ۄ�ض�m��>)�LO�H}E?g��1x�@�	G�X�� ?�iҡ�����g���_ ��v�0���&4�Q _�+�/=�2���aR���Ue�`.Bj0��_��`W1 �5��<Q�F���O��ټ�US�/�C�n� �w@�8���ڳX#���h���PT�PRԂ�E��z#���v�gu��;�`�x��L"3 ��,xw؀:MJ��-������G送�'�욹=������u/�9]�P� 
�6�}Fz�����4Bf+���a��Ǚ�~��㞟4��4b���(+@������K0̕x�c ��ծ9���Z��1is�[ܪFi$�I=y�hEv���^��1�+�B�K6�1�v�{��>��K������C4HIӱ�ZkBjd��B�	��<.J*z�֮ϗ��@!t��^�wB� !���Ӥ�����&����p���c.�3�g ��&G�JcNb� ���񌍺ѨT^ҧ�;%J%�-y����3���v�i68�öo܃IY+��8�W9	��Ic:�K�B+�R�{����þ���Cxz��a��I�m�#�#�U��0x��n��(J��QO�u'*��!PK�a,����rm�?7�|t*-'��!h���[RZ���M�%䚸�&������p���8mW��g��e���Ez@n.<�(��2�f�]�G��t�����퍐��9�"�?�?����`
==�A�T������6��3�tq���^a2 w^�`K��h�����[�����ִo�",Y���wj0�ʤ�1�S7k�@N�PB2����w��7��!.�
K���;셉H꣼�"H��K�;�st�Ğ]��K�g�GǾ�E�D����	�� 8P"W��ٙ����	�Ϫ��_���B�a^�nl1j��-beY��t���H�	D�|`�5�.h�b��@�����}�j�x����<��"-=���(�nL!��>�V�m����i�5�tN46*~�2��.;�x�l\�l`�k�+6�X�Du��"(Xbc91gJL�?MR�V{�
pK��O��ޢ|>�ó�5��'p�C����
�xt|�����J`�T
b&��(�?U�B���f@��;�h�#���$!٫�Tٹ��3���b� \}���ʞ�ZB���'opn!��SPt]�SڬH2Y`2?i��g����/��,_�M�ֽ�������*�������$�Z��!�LQ%��'���>/��D�T��|�����q��KݤoDߋSgv�xO��u�n-<�K/4�ѱ����䃟�����s{s��!e����`a��3�W�^{3to5g 
�W�4��g���-m��"}�Z�/�x�/�S>��UC�3*0��aV��5\ɞxS�IzZX����@�1a�z}���qU�Ge��"��U]��z�n��c�B4f��n�֥��,�DNt���]U��P��]u��y�P�t�L�aq�}���a�7�|���'4�g�j�\�d[I�uY����w�!Q-�z����6L��� �+�~B�����7�Vh�M�|��&�|TJ+�٣�e��O��6���Gy��h��[JZ銂t|��j��]&�#��*MSOᤢ:��F�͏?�V7�:Y�(Ѵp ���k�g����^�������\m��×8�l��������n׵M�
�|mM���n}�����ᚧ ꘴a?)��ў+�K�5Z�K�UA���u��W;]�i��e�2�L��m�Lrp�N�ܮ5�;F��D�
r_��6���m��L���ӛt�߅�_��1���K�a�-��`�	 �q��/35zk�%�S�IଧR+^l4 ��N�9 "|�/=��� �ܬY+�/�Y+u���'��D:�o �um=:��@|}��#ff�¡8�����Dq��d�{6{��
��U���gO�"��O���Q��/�N->�^�\��͆N٢�Y�i [��%�#�={'z���V-��K� 4>پ�)���g�PѥV���ͷ���;��i��Tu��O�QO�L�]��.$�;$=��i��xӶ�u^]:�U{7P�%���8�&���L�MM����f�e�$���܎�-Ӗ����І�^�;�2X_���_ȝ�����r�h����R��x�B0�4����:�ہ���7����J����ȱ��K�0/�]�{Ig�	~#��U[���O;j����!d�I�>,ޘX��$��ל�~��B&������U����w�.�;P�ﻺu�̒_9�`q^�!q��+�W�sxB�R��h�-�F��o�6)���Y~D�� �[-Q|%�z�Ԕ7uf��0��W��U���Gw���va^�'��byeC�����s��@����V�� �=Ȩ�C����_�Ƕ>xL7��2 ��o��k#w�|�(�t�5qD�旉�0�/LSf	e���;�l��jHC���v�5T�y��@�Z����X�V�=^��~?�����x�C���g�v�F>�d�����;r���œ�T_:]v��7ӑi�7'�&��*����K��*��D3��_S@��З��͸� wiGO�yϿ���1���/J<�b��/�Y'���<�t��K-t���Ao��?��&5�Sl��qhV�,k9����������+�F�Q/�� �+;P��!X��:�k��?�_��������N�K�+R���v�
[]4k5�]��G��_C������M
�$��Z����^%Y�1�\h$�D&v�"��u�8U�����_�o8�N��,�0--��F��ϋ���*'�ޏ�Y�Y���u ��Qgf���2.��N+������fP7��yYՎ�D1�#4T񱗠��뽯�%��:4A���[�;IE��L�olQ06ya�����*_1��h�q�[oWW�O5�U�X�7��X�_�M�W��Ҁ�*�BQo2Z��ī|�TS(o2<���t�~p ��\��V�l�X&��xPk{8�E9"�؈E�#3����;Q>�k����,֙�,f�W٣� ����i�3�������Lø\���R����w�ĭ�U��[������m�ѧ"OSJ��h21M��kUop�����'C-�=#��޲�����0sv�K��+�Ĭ��A��l�6ЛԜ��B(aJ�9էg�O*J��(�N<� �Ur B?O ȁ�����-]�9`�-�%���m�lwR��^Q��e0�]�SQ�P@Wg����Z����������x�8���a�_Ո=����o��>�_ā\�^rx�J~ruQ��ƕ�ja��9F`��b��崪�C�9����_
GIT�F�ʱL�E(^e%S�$꩝ͭ�@]���Z=�Ew�c�BBɓ��,��G��i̐���T��Fl��'=?G���ۙ�5{<C�n�oM| �S7Y�x����<�;z�C�Ŭ��$5-�4��*&���P܇|r�!�ԗ� �׈����]�^f���澇�p\T���=ضK^TR�Yk�XW	��̷Y6�j�S4hr�O B>�h K3?z���7\����7��/&�By����i�b@�K���=��WXA�|k=�'՗DzeFF���L��Yy��~R�|��_ -!{9�]��K���_�8*2��]�y��_���h	����9l� ��o�Ț��ݗ������L���~+);7Ru����4}���6tZ��sԙ���|��S;�K(�9o�'���4[7A�J�����S�O��+���j24���^V�hY��|�I���*��x�:���C���m]�֍9h������t��-T�}�3�ʃ���� ��:�m���G��m_�6�o���y�����Z�2��}9�i�I��x�)�1��'���/G7���Xl0��ǯ7��_��L'W�?d��ܒ�)3L���������ӭ�DT�#�|��Cs�4�[,q�4��ȳ#@k\n2愊��, ���D�h.�rK�:�B�T�^��㐿���ً��]@6�s�#d�zǨ�l2H�Ro�Cq�)����n�D0�Z�P�f�����U�����c@�X�9��@�*���'u���R
�3��-����M��:[R���4�!fN�+��M����_��H?���rݒ�U�ɢw^�`�A`HB,g���� �*Iᢔ-o�(w�/Z	�1�'�x�:�3��v��!��5o mI����i����4�^�/W7eE�4A:x��{_���+�n)��f�3��.uViR�r,�ꁤ�Y)������V���#f`��݋<Ĭ�Fr(;:h+ ejTB¤��u�d"�p�c:�w;���Ar��hF�� ���RY�<�V��l������tx� A�Q��#�T�y�/J�;zI7e�j�V�kC�/�OE� �oq��Aq���^N�,J��Q�,'y���4z ��"�;���ֱԉ/� ����o��%ɒ���0�}>���(����{�#z��h�h��]x���!U�{�]�	�T:S������Y�̻f�Z3X�;D�<(e}�r�����_��s��E� ��,��̃^����Ǘ	���xOB��-��!�9�B���ԑ�ר����iW� 4�Xªߪ��h~,i`h�;3M>8m�2d[Q�l��BO��w�&�.�N�N�Dm)ˤR��b��>o�=�[�����b@(:!��M]$�;xx�mv���z�Mw0�������:��I˶����}���JI�
��1��{��Q8����r?���J��HU�j����A:_�'���4w��ُX�uLBIB�T�\�Ş��ϡNz������#&�
�Hԡ�̲�)�s�v[+[++QZC �����B��"�:��[�N� ��ˑrR�cyk%�D����̝����"���X�׆�ɑ2S����8��������'0U~6l�[zgȄ��X���(�����(*[�i��*��M�1�>.2�g{[�~iі�� �53`��nU�^���6F��VJ�q:�7apOKUx��,e6d���PXL*��b�z+OX�%(�x:��"��[�	����M)����/�� �V�g�8�����q�p/�c �o8�J%h�j �����o9��j��e7�Z��w��l��4��-�ݧ���;9��a;(�@)�����yMCxC����'.H�Ev��Q�J�±鄸�R����@�CjLpő��c��[�~�(K���)�4�K�1E	K{wr}-��J���S��!���E���䱍^����������3��H0���VJ���_`c�a)d�T�R��콽��x�����&e���`"/�c��:|��, 8���b��w�;$A�������*Dд�g�ኀ�G),���0�t4Z,b�*��.I[� ���mFg(��j!c55�6}� 0w�exp���cp{��;�Ձ�S-y��������|��O�|��[v��ݗ�����ٽ�\����Խp�p��Ra�m�4��x�����uc�sX���o�Iģ[=S��n-��ʊ�h�8����.�|���0��[{$�`9|_���=���ׇ��,�b�a�
��'N��\��ֻ\��VX�U;����pi�5L̴���j�3����=5� s	��e/'Ε�%X��y��m� ��l�l鬨Hu�U�{W6���8�l��۟�w����q�D��mۡ�g�_{��}��l�c�c��`������*=ʝP���ъe����Oڰמ�z��V�r�?ͯEk�>j%���ܨo6?ܚ(O�"���b�!�_;�qP�=�K��.�{lMIS����B������`�hy���j�a
85�T���v�Ϊ�rt���簐����BCk�2wG�����e���{	�-�a�1�����e����G�?���;&� k��š���]�jڍ�3L%-.W�(<ǒ�|r��ܨW����;��d@�rѫ~�M���W3B��-�կo��=��	C��F��J�kk	tȚYW|�G!%�������]�ɟ�C�\9aʠ�l�s����JTm��G�[���"
d�[:?��C��B[XyOșjDJ�M��ؖU�2�*�!����ϙ�m�|�d"1����!Q�!k2�$$Y�owL'[ ����ŧ`XP������Q�?�d���_�g@B���=�X�lF��f׵w�q�W�(=G�� !�d�J2��
}��s��!��������rM�`[�_���r�έ�L��"���n�n� ,�z�X�%�$�F�58��N1+ ���o�Evq��Ӱ�X�@�U�w5��UǍ�z*�W�C'5�[�D����}S������]�=���XWN�I��2�>'fv�̇����W�כH��A�ߕw�9��⏞�Y�����/v�%��EnT������!���(�BP��S���HҍAZ-�����d�����J��u �w=���P�[���Xu��5e��&,/�[�O>�,�SO�! ��4�]�p`x��rp#F�}�y���L��4r�Ktj����)��U�I�y��$�d��w��E�+����e���~>@��x ������a��uǱԔ��~�l��w�0����F אI�����$&+�vN����w#p���{�v;���۹����}V�L�;~��-$]���BǮ�5%|v���Ξ���]_=��?dֿD�����0tʹ/.l�/&+���}[�q�`.�J0L�G�4_��k�l��k>����;���o�$���
:�$�ǧ���k'!sa�Q�V�>$zp���d����DeomA�8�'������F���N3����̐3R�c���7|���Ɯ��wv��#���9s���A����`��Gމ���&�+`)�27ko݉h���%=�Qp][}�<�z˼���濡D�y�qy�3 W��~w7��~q0m�Z�&��L宆vqtF_<q�M)�˴ܾ{VypOx�ҭe_*���Y�Pk*d�Ȼ�C�{�����"�4ծ�b��6��s� �gΏLf�Ē��������Y?��`��馿[������1>����C�%�C�x�ӽ.�a�t*"���t�����y�A���d��Q4r���l�)X'F^q�)�\�Ǭs�LTT���ԩ�Em�ڐ���z1�o	��f;Lqm�E�.���<1`֥76= �!8��s =�bY�ڴ����g�D�,;""�6��4�����C��z�F���k�9���\�`ܛY*y�,aw�[�K%��y���u���q|�m~L$Av��*�ܧ}G�ύ"�X�>!�����W4[��xL��ub�B-����%6᮷@�����Q��G��OO���!�ę�X�l�S��.(z�9�����q��Lp�%�V=J������B��-M2y�|�k�(�1�O�e�m�2��$���A�҉X�+���b}@�f>� EKz#7�v��| rh��M��"��0�g�'{���X����l�庫t���P�㟾�4Y�����|����@��w�)�ח��vݱĠ{��4�4�lNS.���Ԧ�a�;NCs/|9���������1�Y��|z��`/��2}�����	�m��H�$�!|{���	 �lÂ˺Yt�"�&��M��qP?�gr2C&jիA)L����2$�rn�A���j�3F�G��9U�� ?Wx��P)�F�+'�p5�����?�m��h�$�K����XS��shqXe�[5�6vcҬ�r����ږM��k��~�*�@���YYq�닾 �Q��G0�&�'9��m��J���)�k�l�m��g{;���@".��5N6-�}�Oi�@v�iE�-��!�<O�4������1ˡ�-*��c���|��c,��^��!�X{S��ior�6����e��l"5��w�� �b5���p�L�f��`�O^Y_x�g�jЙ������ۋ���"��wfn����HFV}��AapeJ�a:΁��6������A�ܴ���c':�a�#��������PakȤS)j4�Ю������҆3|� K�fju��T�\��2��N�����������f�����"�OW�G�W����a���zѨ��Q�4�^�3�	��a�n��A�mm�iD�u E�!��z�|ri�r`v
�?{Xy;^����/��b�eb�O��ȹ'�w�ז��$���_9}�U�#|:>���!��� w��|n�2\�E����1��7�n��#m@"<@"ȉ8�'�/'����U ��+��������;�P��#�R�}��-(��+�����*�H����I���ݞ
5 
n�e�붯}IL&XV,3�y2�㼫�4�Z��#���#_�f>��;6�z�.�,�^+m��z��7ٌ&���0��yk�=���(�����؁gC��d���U�_�E�O @q�DӲ]��X_�� ؠ-2����#��4Ķ�"?���\bl��/��"���s����Mg�'�|��{�����:� �7l?_%�O�!}d�n�!�!!�	��4߾�,�6�E�M\g	�D5�I�1�������-�e71*%�������8R�� ?%�3T��|�Y{f�bhG"��Iۤu&������o���s����1�Yl�4^."E��WQ 	]�@UI(��Zq��K��t(�]�?��[ ������8r�+��g/�9%"Z'�϶O�~��:dZ�!�Ds=��靆��\����y��<��(�(�����fd}�b�����d�sQ/�2�j֔w���=���kn�1yt�p��)��N�\u�ABU�c�0]�CVi��U	�����ݩE����B���!MS�^ [�$�u(]_n8�����x��+��1Y�?�m�ҕ����k�z�p�5�L�c���w�����uJS1T�����D ��q��L{������ТQt]��Q�2�ɗ����4��F����料3�:�%��Rg�n%}�(�#	�u#ߍ�������j��O`�.�'� �	��RX�4��-��d��I�##�[���VSv��n�J������`�ik ��hL)kJ^�����d��=i�84��b�O��ǀv��б�P~bG����dǙ��Sg��fD��mZ�jXz��h�S�7�T��� ��ͼ�QY��WL<���V�&�²�a��t	.�e9�DѺ4�:07�j��w�q�o��l
ߐ��=����7���g��K���nW@R4ͨ��7R�ͻ�����:s�^-.K'n %�!�]3�ɣ�ߊ�q�4�3���|�~?�����R%��o�����R�����?.�(}�ڢ����m�4w����zۏH��B������5~�c�߻y d�cK6Ba_L�7^�n-l�����`{��}���1G����-r�~���Oܚ���S

��cF�X�H�E]�v�3و���#ː#y�A����@�s�ډ�JpJ��B��L5t�q��w�MK$*&��Ҋ�`�rփ��V�d����*z
���> M��&��߼�A=y�I�>�ewuL�I�Q�16��D8����Cd��r���b4�J�5�h�Ͽ�_��e��a���x� �Z�J��,�D��0��A����&z��=�պ=�kށ���:�Z�C��~!{��Ao�}���kz�q6�ٳ��88Y)I$t�I�?=7�X� �U�tz��p�
5�1�=�x|��k�k ��㓽s�L��{��E��뮸�]�iE�`@@� .""�  ŀ Y`$�₂��U�̐$QP� HΒs򯪻q��u=o��?�:5]U���>�9�ӥi�Gk�"�?�[��ց����)�]�����a�;� r�����i���"�����޴�Xl���`��m�@}�(x�%6�2�����c�����F�¤M���M?�M�Bp�	���r���� ������V���;G��-�5��l�u�J+kPڵ'X�uGFIjߎp�XZ�T�TAlf�[����1�j�&'*s #����܊d9���m82e����b�س��*� r�8�1�),��FӾ6�e,��w���1;?�-a�:{,���e�C_�[���C�/��Ye�����i�O�;�og����p�t��(,gV7�!ԭJ��s6���.�0������y�M�h�!�}��|MOt�LGbï��c���j~��1�ĳX�����z�}��Т���x�aB5��
F�;�~���S�����/�R�BL�+Ua��^W�NlѼ"B&��Z {*/�\��M�M·;�9� �v�V��q$R �K-J�o1�� ��v�۶K	���z�����Ά!�G�+ف��y�_���8�����o�����*X�|&þ��جΥ��}+�h�ZJ~!�xڄ)�-�/��:
���)�!`1{�u9�٧z!zCX[��c��V�R��x�ڰd���U�P����&���ry�᎝�@�A�"��hf���9��.���Y/���`����$�Juگ�/a�d ٻ�w^t�	�|��&vH�S��A�޻AldE��_���q�0|��|߻n@���M�ⵯ�xJ��⁂���r�o�X�)H���F>���8hMt&�ӿ���ۡC�V*��m_�[�d�K�R���6�;/���Z���י�Cl�����FS)�ZB#'�\�ָ�f׏��1� �w<k�=��q�(�"e��|�X>�	����O���D�T���툴�.���D�������2�j#�@��o��!B��z��N�ހ�˥�,A�)@4����s�/�X��*ܹ£K�p�b�R�,����TJV0'�x�Hk�ol�w�qY��
`%�)�";��e��\�ǌaK�
�׼G��/Q{��L)g�.�u��~.��o���#������&�iTZ'=�=�x$��$�v�m�(ǰ� FM��s`|��q2�A��m�M����HM���bam�dk��|��[�%v[ß���Q����o%�컗�,M��c�;(�l�M�MG�d̪O�;�ZQ�G7m-�l���K�c��)�>k�Z�����)w@>�����=�	��{`ѭ�&è�Kzo]�k��|-�e%\g}��}̡Je�^R,�M��,R_�=&�r���ĝ�����/�"��Q�U�6c�4x�©�팿A�����C���A��M����+�x%��6ੲ�hn�F\��y�O��b?g��N�a>ݲ�{E���~|�������CL�&�4(-H�l��_�M[Y86p�����:�Jb�5�a�p�-}m�nL�{0�v9���_�jf���6���-R>9b���>w��O3�O���@#��,��3e#L����l���ZP 8ht��QȈ�I�7@����ҕ�A~�A��J����,���Kej���PJhilk�����Wt]~L�l@�1��e/����b@j�J�L�N��8���S�)�Xk ~�� 
�W����cX�tyG�������dR����)x�œ���V�<��&�E+�M�@������S��Д�m�ࠆ#f����\���C��7U ��2XJX2�1�]�섽�<�X��XJ�������H�ϥ�pཱྀ�O��уR^Kԁ*?�<������ �xi��!�q����������&���/5).�x�O9c��~�]&0]��J�o�#�����{Fd��J��Oc'�@D�j� �F��{<�.ƙ�X���E8QE��T^j����m[��,�ZQ L+�UK��A�X�>˒E�Ya�Z�ne��
aw��%��YI��2�CT���\�Or!s�����ۍ�@�{l+'��\����,zC:��z&q��?R�қ������(/���XTfZ�N|����%�xU	(u��-h?/;��� ��c2�!rM��~����Lx����3�=��������6���ͦP�� ��(�]��jbܙ�݆0̧(�E�&��[�*���y�����aK#'(h'z\�73�0cs��G`0t��Y:��S��~CL$,��RȔ�^����G&��z�Ԕ'nVZ2��niT��U�v��&��*� �#O=!�o����c������׎
� M�e/T�tI�n�N=��:�~�Y'�����}��c'���(O5Y�;��D"kk�����S9[q�
?3Z�H����7j�b��}�e�7��#S�R���K�7����և�g�C��r��
 ���������`W��9��Pҁ���bsk¹��-�lRx�cv��#��L�����OY��æ/����l:Qmz뚓��B�o]j��U�6+zq��|��W�<0<��m��$�3R����	��쐢��?���ڷB��j��9 ?� �!"]Ʌ�Cn��p��%��e�KBAs��cD����nc���� ̐�	;��ݝ�j�H�Ch��@%���J�l� &�H�ܴ����i�gj!r���J�
Z��2s�[�N-B)����|�e�N.�w_	�%�+Ͽ`q�I�Z�e��_`�J���D�^}���ȯ��nkPY�nV��m�d>V��n�n36�����N.�=@M�����ޘFl:�&�BX
p^�>"ŠN����	���L�^�R�Y��<@^��H���oT����6K|�=�xʹ��l	F:�1~���",�G�g+��ȝ�0��=�����k#�U�T'��^��s:Ժ���U�� �N�T#ʚ{9��&RC�������Î�Y ���[#z�Zb6���[�5�����co���w�6<�`���uE�i���`RL��	���}�%�ݺ���� ����ODB�;��[��ͪ�����Kh�h�ws!�t�ZK�_�p��4GՓ�b&�&$�L1�rB]��T��f�{a}R	Y��6�n��1��A��gw�y�A��?!Ƽ~Z?�c�Ύ$�Uկ�����(@E��YAE��,�j>�[���g��KQ�%#�Q��_�a�I|~R4�0#�M�~?�F�.w�.�?�F9yU�A�y�%Vxze�+oY8/�y* ��n��G��;v�܍A����X���L�漜:T(4"�k��o�\���$w�~��2�}��|�M=���| �u��Μ�Y&y��VD�&��W�����O*c=y����{��Q���$��:ӐM,��8��k�m��h/e|���n�K�*b8e����-:L_qAE�5�4,��j��K�7�N�Q���m���H{��P�M���?�v"}��f*�Hl�Mϥ)����P�P��3�7�pB��:�,�#�E^g+6[jϸ�}���]�|v������/؟�<�T�����uK�x:&>�٣��YLP��R���eS�Y�`���A�X��L�jn����4�r�!\B����A�Z�m��,G}�k#�4c�f�i>�E#��W,3O	�Su����I��o��@�i���z.�uO�r�C�QG���0c��9🭒.\�����5�UG���ɨ1Gޗ<u�g4�@K]��<Z,-�eW��/�-���ǫI$��c��J�<�6�O0�nzq��_����T�U��ѓ9�Մ�n�O{�e���}�A�����Zb����ǡ����H�n�p�v7�=�~�ȧ�ϴp�%ԭd�z8x�E<w���_CJ��Õ�W]|͞�}�l��������>!�n�Jw�L3��n�]C�gʍe�W�,$��C8q��x�`=��ĔB~��(lX�2�����}������>�߇�������}������߇w��&Rnh͔n�_��IV�{��Kg��b���O��U�wM�7fM��ow\�tڞN�(1��V�r��Jz<Z�����k��+��k0��a,�A4k]��&G�� Nk�>{t�C�V:�gyA3�#}ETv����f����ؽV�}o���^J�RS=4����[̽�7�3>veJp�S�TM�t�.8[����f�A�2I�q�н�IU�2�+7W��%�ɌoVʳ,��//t^I��6�6?�>#������4���6�ʧ���?�V����L���cr�-�}iO/]�L��ط�����<|=j���S��RB�=V�`�����9wbO)���a����o��������$��G�0�J��O���g�v��y������ �, ��\;$�C\"U���rj�	�,N�?`'�5f3,��.şX������R�7���^�;�Bh[�{�S�ŏ�p����y�^���zU���_��8[��~�m�m���Z.b��cǿjpGr'Iڼ��h���0X.7�Z}��fn����ޝ4�J\|j�"�#*az�+9�\Ò�y��vM�&�ZW�j�l_,p	�Noۦ��oyf;���t�Һ����N�^��0��_bʵ������il�>Z\t�'���h��ө.�tO�z%�H�
p�d.�B�z]K��#Yo�ɩr�h�ҎBKJd
�Q���e�,M��=�[�3,���F��ќ�g����"�x0��위_��^�O+�7oڌY;A�^��F%#wv��.�`�ǹ|�7��v� 1�Gu5͚�Ф�}��2K�J����"u�PO���#�Lv ;�"S0n<a�Ԗ���Xӹ{��P�d]���kp�MaW��,�Ľ�����u��[(��Mر�7D�I>K_�y&/���c�j�q+�OF���Iuqj^��A_��5�lXa�CZ�dh[݂n�	�`�5�$��L=���H��/-22�K����+Nݶx����8_�5�.r��=��nh�_1�6~�N���w�P3��*�?��p�2�8�a�#wMU���m�L��p*�mwﬠ0�0[��yib��a�j���4��8��L��v4�4�^���X��m5=�$t��13�^�~�o07��7�k�}���y��]���l�,Z�u&�o6�&ee����>ʒՊ��V����r.�Cm��_g�{%F�g���32l��u[���'������C���j\���%��X���3lZ/�n^�uIzhV#�\����*Bcm;�4ܸ��Z_|6���,�|�䎷�)��`"נoIQ�b��6ȿU�1�C�ں���~'��BЯ; ƙ���[��9�%�a���ř1�L���_���}i���18v�_�e�\-Y*_<�;���oj��a���r��ݕ^�e�M���I��n��q�:�#l�>,5�W Y8��挡Q�9�>��_����u�Ƹܻ����q���sM�$�2|�.����Q���w�bNR��7�Du�Ǽ��z?Z�l�(ꕵ2���lޔ!<���R�H@l�)WW{��	|m��y��FZA�dn�K��pi�<h
3>��v�������+ղ�}ߡ�T����c�ϑ�֐S(nmVHjN)ƫ����b��m��vJT2+� /��&�k�8��7)S��[�\�a���4�[�����lm]l��6�<�zr�X�x����x�m��Ya��Y���QMN7�V��s�t gmHM�@�xJz4��m��G#4�����HC��FG����ik_=z��������낦[<�uZ;WÉ�&�96��H�TZ�t2�j�m�)�� �����}�#�"�����^?�=�̍�ʍ��[�qi�8o�r�·�P��w9�	k���Ԍ �Ѹ4|]`k�lu��ۋ����%f��YSL�y��;ȑn�q9}=������1��}��� �Uk���q��-���)��<;�����/6�'�����h�gId�۝,�_����Tb}��&�]^uC&�4�����©Ǒ&7�c�����9��V1��חT�tN���c� >�й��&?ߨZ��)���G�nd�,�����'���/z��Rh~��R��M��������o���	�նj�qF�MRՑ���Z��vi2�Wejx�*������ :�{���=E��[�ήܚ��'}�D���Ԙ6;�L33̽��1Wh�څ�ݶ|���\�`^n����!e{h�Z@"�'!B��H�B�C�0����I�cT׌cъx�{l�k�
R�<��sP� pj�w|ݧo��$=�_TTy��c06�.k�%��G�Ͳ����\?�H��,:|���9[59��/�5�w7����)oSeL�פ޸fK�c�6wߟ l�a�j��V����?�a�p�9��Sd���R��׌R� �j3�0�ܙ�/i:�L�� /�l�X�:�h�ɇG��9������t�믿�Z�L��-��c�[U��}�<1�G�<����\-ێ= �-�s��QI�a2d](G����7����N���M�rJ�g��� J�ހ��4#n4d�H)�m�q�����A�D<�s! HB��L_�hӉ&!~z&�TԍE�lq^󣒓��΍74%;R�Ǡ�k6t��gMέ��k?��a�� �R��SMVX�ä�د��f�!��b��B�֑��Iʛ4�xf��)��������[᫦%��[���H�@5��S9x"���x�uk��7�D;ܼ�S�u�����$�&���������j!�.�@q�(�Mp	m1=� �A�m��W��^0�W�m��&�1m<�;�+��/��˄�] �;�������H��4ܑ���y`wN�/J��yyf~�[/(2U�Q���~��[j��ЉOx�l�ι�ݷgj���/�(�I~)tnq��w��y�Rf,���İ`���5���ݘ��uN�"�Ó�u�L��L��r�w;&G]��5}�Ѝ��Hl�0l�O���_,���H�T�r��S�7A���͏W��ރ�V˝�_fb�uhx�!���*,���D�Fɘ̤���X�9Ob�O�fY�y_��?/�h}3�*�r�=�8��J��^�_ev��͘���y�u��?���v�@O�|�p��Ə�\M������:�m�-�W7I�6��`l\T�n�:�4�rWx���P�Xl;*�Ĭ(�����=�����LlK+������� j��ݩ��7�-]}@��h����+gx�2JڍS�P��4��:o�ju�oB��d�aoF�N�n��V���ߦ�>�l�=�^�W���3'�>�40�����K�U<��m�ٱL�s� �wӲ�WI�r�/,��ıT�[TA��5g9!�)v˳i����R��N�6p_ �'N�դ��x����ϔ��M��
se�]�^d�y�	�	��e����m��c�yw�����A#k�7IJ`��/�����k��^U���9)սyST�Y7��.��J�s"�.N���� Z�ĭl��"��&�A�^��ç�9����盜wv���ݚt� P6-M�s9�������r3���_���������m&ҙV�w�.����B��m����٧WV+m���M��!ϭ2\q��@�v�1�Ⴎ
�43s�O=��|Y�[�������+�g{��\Y�����
�v�+� >�8r@V5'�a@*��.��s�ƚz�����dZ��j�Tz���/�4��L�����(6���x	��5���Y��2�=����r������±�'�w�W�� y�ܼϻP&{�Z���l�U����� ~�EB�˩����fh8�+a+(��Q.����VJ���C����_I#��4�}?	����,A��ͅ��,=��ձ�t��2��Ykt�zCɶ�P�:��6�Y�9��`�jz��/f��Y�nFX��J�	��Ǔy�λ@(��$ ��)�����m���"�?PrKٷ�;||��9��-.��^��&B��$����s%�����'��V�ra���� �R�$�q�M�:�,:��;�b9�\K��i1R�������Qg�	a�Rj�ə\�K8[��o���n �X��ej|NCQ^N]Oy�Rx�[����7%���P����+)!�?�0�{GWI���$������e�eZ#��#���9��^��ƴ.q�1'����^�h��m���]����z?n��ޝ��-Ե����>S���)�m{�ȝ1}����	�,b������-Ԗ���c��__�ʘg5���Lf8\a9��6N���k_q�CzI��8�I���""�`pj�\+D_o�����������E̸2?�[���D��fC
��b*��+�<X .�\�5P�:���O�S���oj�T�r=0U��>�+���0�nEi#݆��h�_й��=����;9�)�QS9gr-�|.���u�ѳ�j݋��tu5t�i|��ƮhI%�I*L�s�s��g�9yb)`ƣ�����GA���r�A�`Ͳ���{��Z't����p���/�	_�6֧Yav$1�@�:��-�V�8v�M�1Չ��(P qn�]�?݀^{����1K	*h��`�����$�
���yS{�^��u�T!�5�S��UK��:��[R���ή~ �dL_)j���{�Bi��[q���?�8����R���?ٕ�CKb斃?똈�,iđ����s�)������k�l�a��=��"nN,]�eZ~#��C�!��F��p�1@#�M�r�����I���������BRϮ�j{DBE����e_���e����h�u2�P���Q��
��=��G�d����{5��!ݲ#���YݒR�Қ_�/�b_���?��#��&���
��RSWcb���F�G�����L����.[e�n\�/Y7�Z�?���=w-�u��~��RB���R��G�5�z�HW׬�:�ʥ'1���Iᖫ ��Mɏ���g��=!�Bl���~��OӍ�H�Փ��>�=�q	��ܿޘl�'�C2�֢d?�N�p�Ǔ�����4m�οhu����~�
j0�,F�)����'gt]A�<�B6��\eU�6�1v @�~�����v�:	�ϝ{��!\";��'p�ΥQ:kA�[�{��ʈD��������x`Zݛ�Ni!�-��50�Gx���N�y���_+����%�o[$3���P�����0��h��8�c�����f� ݖ8�74���`{��g�Ǉ��Z����6��g��C��Ԕ�ICkPx)iȬ���y����axK�d�	��{�M}1 ��Ĕ�\M�#s�_?�~ez��s��C,q�j���K�2�prR\�k��̹"|9��NZ@�PO�����!�?��:��?���ӂ5
i�HZ�{���c<j�Fx�WA���1�]�9��D�ˠ��jo+�u�^�������O�v�aZ�����P&�zAZ��l%=	���x =�Q_m�ǔ]%��ߖߦ�c<��Ah)��-7��M�>^�#�?���+E�W+��Y.�R�5����s�T��UyDUI��T�t5n��0)T]��
E����Q
�o�p���/S����� 1:�Y�\_#A��2��[�%�;K��@�p�����r��#TV?��!��������@J�q���?2'�U��:�L�J
N���a}�b�Jcc"B^�Q�/ܐF���+cި����{x<�XL�V��#!�I\�������0s����=����a�٢P����Ǐ`[�CO���,���FY�(�y��ۛk	�1F�ɑO�N����#Jv����+�3��m%s��#R��<�⚋9K����������U��ofq���߉?LK*���K�ϑxQ���D�h��L���ui��]�#-"��d^�e�~�D��۾I��b%�G��.�+8�ߪ�Ƌ�3bq��<܁�\�0imw�!"I�ÄI�0�u��.A����u���C�� ��Q�?8Q����$Bw��:p=K?�iW]@��mq�B��A����F3s}et-G�ú`T�g�l5��j@�tw�M��
�J?�yh��Y�rGF�:�]@pGC��Zo�,��0�,��a@b|�p8RwR��aT�W~o�>>��@�ړ����uS��J~��M8&w��+~��?�p�;�t�h,lT���t Ը*BOR����;�C�AY�����ʘ�X�[�nX��p�@2Zm��W�S�3�ͷM�. �Ø���	�s.��)��CZ)i�9���5�f�D���F"��c����ŋ��~.�Hs��2b�b�!͑�����l8�`=��+����*`^�#��o�.tz�����m�Lm<{-a����J�iKL���%���'�/�g�=jP�"��1��(�Y�lm8�E�罀�ĳ `"��tR�٦�{�b�It�\B�]m��߿[�q?�ǲܲ��z�W.�� ��,�\ind�%"��W(zAC�B���܎m�����¢�;H����V�h�������Ѷ}��'���c���m�&Ps�����Z��Ыj$o��Jb.��N˖a��zp':������ˋٞD��7���3b斜�+1��Æ6�0q�V/Ag�L-]ꔇ��^Hc�}u��mi�v�u?� ɕ0�nȻ0�(
^��*�m4Y��BPY2��bDЎH,B���RJ�5&�X�Nb:!�{_�|@�'�@Q����B
��Lb���Y)=�;Ψ����@��y��b���Ao��f�{��ό��	�k� �k��g����)j�YCƇ�h�'t���ɫ��\P�䤅�Z�精	�'s��$�&TF�Y��R؅����`*=��Z7<	?�ڟX��N�����.����G��%�7"��ǐCV�X��M�ʠ��(o��F����[ �3�#��t�7%�b� ���zAm])�;�;p�"eK�9�E�| �� [������K��>����ɟj:��5�X< ���F��r���b�ϕ)�A��0�q��J�&�#��
?L��Ϯ�㳮gl�|[t��2�������ϦY�ƛ�L�Bn�dV8�0�X�'�	w���V��F��a?u����K��	&�?;���!T�� &�CD	�겆�Oi��0�۲�D�� +W!�ҋ��v�D^��}W9�FRl�!����W��[VLv`lII�2�,^�V=�yJ�k�g2V���L��woF� .��+�ͪ�a���}v>�H�^�����=��?ƛSeB��w���GMZx~| �{�����D/��{�h��v�\�_�2'�{Т��oXu��j0��a� �#k-x����7��Q*�����(o�C,&%���n^H���,˄���>7�=1�;��$�J� )!����O\�G�C�xo�ƱcJ$�<uC�����VB�k�����S;�@�@����In�v9訟�<)�9}�޲r�g)�kG$�şX�;�j\\�6K����d|��я�'�8�4�peO�S��ߢ&q���I��O�G\ѝ���}�l��_p/��H�O��/�Z4��(�x�tn��`�'{<�/7��W�e�t�*4t"�D�����<�01:!��G
R�z>��ȼ�\x�h!�a
��u�K}�d���ƚ.����ܡ�}aK$$��~���L!��L�?��=V��x`���D��:,�+1�+D�Ê����I�<;��caN������(��7�Ԛ*��F���.�R@����D��,J\��2N�^$b��e�s��ɚ��K�ͽ8�;�p>Կ�ၩ��( �f���sm�+2WB���WC��W�4��)J�&�� �ڋu��.�c7�����0R��:�|d�L2������ �wm��}��E
7ܙ�#������������!�O��e,��b����CK��yc�`*b2�!z{�����@�6���/��m0��A����՗�y��Z^��Ⲣ��ϝ�\n�<r�)2q��^��)�a�5�V T�ܜ6�)�C�(��Mb!lw!?U�r	8?k�#��	�=����>��r��kU����Q�Z�g{Բ��[�x�]v=:�bD��ҹU<�����7���c�rɕ`��{ȜY�B�ܰ`N�_pHCs��&a�X���ER�0��i�P��A�sH� :m砵M��$2��W{�1�j�nz�?������������P;��ϪJ$���;����W`��Ӣ���Q���0���RƩ�R�$�\k&�;dr� �%�=l\+����&X�.$�F"P�s�*D)��}1����&�r��˩�9������	�����b�D�b���4�c-5"H���_�M�q�&
��k��7	�����~��Ab ޏ|> �)j�0�����C@r|��D�^'�;P(b� ��?ݾpۂ.��t�zn�:�rd����R��dH��Ȯ8ul����������5�j��>�?m���N�_B�ٽ}���!ma��OE%
M7��j7!�]J�m�t0P�[�%��T� BG_��Z�M�+�I�D���F��&��ԼcZ䛸(�1J"_&F<��,��r�N�O�Kao��-Ý4���?��5|�<B���a��xS�g�����9��/M[���f��U�mڌXn��GY���׈���k����L�/�~k�(���w	r�Dδ�4P�U9���	����i��Uo��T�������#��b�����<��&�`�Fѯ�]����-|��q6��J�Ԍd*&Z���"�r
'����$���ɦ�σ0D���d�GM���"d�_�`�-��%�a�*7%�\n�iɔLW��� g��AL$a����294٫���%;?x�Ʉ^b��X�}��@��d;~WW#/	Ӱ�JV�;�r�3�J����Y�`n�
�$��
�DX�'~,��É��>�ҤK��%�e��A<_���.	X�@�q��
��#����k���`�qph^j1䦠������绸#5�x,a����)����{�[�qj��C�߫�d�����\ż0
���Ejv'���b�Ȍ�*�����x��L=|�[�8xD�=B���׍�c.sq��xG����e�]X˔��_�����2�@�sd��%���Ǽ� .�3O?�/��J�ﭪ�,�ݦ[�~��+5����8�b�U
�E=�$j'c�h@�B`-|+�r�kq�[l��#ۿ<�_������"���ͪ�ck�XӇ�6�G�^at�;���OT���,��KO�������Y�I{x�/B�R@~b�K82�W!gL�/I�ו:%�IO;�Ȯjg���/�70�^(�ͩ
{���z�7Ӽ/߫��m/�_�92�i���cý���m��V���q�k�&Վq��Z!�R�ڗ��[)o_g�����ez�ԛb�]��+��v�s)swv�5��q�d�ZY��P�ԭ��6,�
���z!;"��sl�⑌:������,V.h���s��->�V\�뭹�8͸	�����♅kӵ��)�Z{�##�&sii���p���X�n��X��5�pA��M��0>i��ʬ�d1�e�s,���\V��g��[��U�l-���/�4��FgLS4ѵ�QU���Kvd���EڬI��g(���.ɏ��J\���p��Y�tlؼ�џ���:������\]��CMuVj�[���g8D���bV�#0��o�#���v�Am߿��B��i�����J� ԬLp�%�!�955_� ��״��_���ްG��l�>�w���f?a�S�ݔ��䛌����ڂr����K6_�/�eC�������;\�'�FV4ί`X�.�&�H�	l|Р��}�R !rY��[������P�ȧPk���*�����S�Ғp7=�9�{���ˍ�yOf�zFSs�{�i�LFG�\眇���S�	[gQ���¤\w"����3�Tǎ�[�	/���H�G��|j��P�|��?KI'�z)f�5�(~4�����{f~[D+;�Q?���)���YD����&3e����y�C��%eU�9�q=2Y��O�iM�f�y�5���̠���nB��/0́�܋q�pR���t+7R�EAgO-v���}m�Bg�|7 �"���GRhe���C��lv]�90B#Pf�@��v�+3��`�ߐ��B���������!�C�\7Oa��Xz�{���O�+UУ9x�|N���	��V����l�os{�WŎ�}�
U�;R�lN�Tu6�ǛBw���$8�X�	�SL(�a��="}	ڽy�Be�E`G����4�ФɨT˥����-cm~���X~~qR�ͻmOqu�R�S�/�Ew2Tʉ����8{�Lt��i�w{X\֍�(�:Ư�/i�Մ�/�MlF�E.�5�F�0�h�/����;����*����MvRc�c�N�OU�� ����n���)�Z_j�q�2�jͪ��TKd]�e����tJs�i�_I9/:"a=]�M0�G`��{�'����^����O�>V���
��(c,1]-'b��s�W,�d���_���a2�q�>�^s������
7X+����&�5�:��eW�B��_�J{�˶9���4.8��-�g
G3��d�y��;�Uz�:~�n�]},�G?�<���H�f�����,M_s��U���>u[B&�������=���i;��k��6]u���)�ջ�l�X5�ݹ�pu誱�b�;l�y��gD��<t���?x<����꺧1���>A� �5�4#�V�ط,��.��xE��XFM[ް޽Ŧ��y��C�����k�u�eLs�һ��r
���x'���^��fq~p�f���Ma�X�:��:���KhNmb������=�}tsݡn�
����ߏK�7}���ԇ��?���A~��|e�����C7X�ikWl��������hW�������{�Aj�m��zx^7tnR,~��a����Z��N38j6)�;�56p�S�,+7��b�ji���wy8��9~9��n�w[��D��id����O�)�n��jޗh����4i\XO� �������&�
�Y�����x�Y��8Aw�u���a��NPW�L1�n���8�Vڧ����>�D
��3/�^0�
9q�x�\���]����9���`�)�29K\զ#q�>.ne٨Ñ�7���I�Vs!j��z�v]~����A�p�XU~��� b|�Aih�g�ӌ��{m64�s�5/���,�����]��b�{;�6��{5=q^rQ��K_�-�3#�^�/�Z��PM!�/U?�u��"Ͻ�'�n�2��r<�e�R?Ԝ9b'k
��ճ�м�m�Ӣ�G�[�H[��bw0z��n���)v�M֫EۧT�&�7\�ʞ:T0�v���rs��u�%��|�2=4��y���3[i���t��;ÉO�k^�N�9N��S��R�|��5&������͋4	��d�R!Sv���������g���mz�o�gʐ�MbӴdSD�?�_����A�:��ڝS��3�����8�<�A��Ow���D��*�����p����;�Yy��<U{�~�c�d�!��9��cҽ�d�)=F��!-c�{;/�ջ:���49��� T�[o���eSÅ�zǙ�a� �U�ѱF\��I �4ިZ(}�"Llz/�Ȓ"[��н��S�TvM�g���wS�:��B*�w�.=�d���$JK�~+!��� 0�+�m����7�/h�G��u�������e������N)΢��A5(�E��Ŋ�L^��h<��I;�x`םG��;��f�|R�	�pbo8ߝ}���l��m�URvq���gw��8zr���hR��}?q����{�e��p~��i��	p�eS*g��?o*�u(S�n*��Z�Ul�m��^Hi�񸑮Ա�[S����u�w�NW8�;��'��=r��W�a���;4�s-�t�ݸ磎�o�LÉ�� ��1ç�m�~��Ҹ���
Y*ˣ4�������_�����!���n�������ğ)߮>�+�5���OD����l���'��}p������N��I���)�����.��+�,�Ub�ZF��VW$��i.��X;�~�Szm�U����.�>]�i�o��ѡ�y����G��T���[+��i�'z��a�����<�!G(x��Ū�xG�k��*^X�&@_�$��Pt�0��8�{5�sR�ǟ$"ծC׸�(�53ڃ�B�^U�׸թ]~�r�G$i�)�'$A�z��e[��@��t�z��/Q�������v����h/�K�ߤm��ҀMX��瀾�?�N[9[K��/P�o�n�R�7��[��]� �-��K��cqzA�G}q"89�UG	�u�sTuu�wX�Ast'��h-0�o�Qs�5���4t/���-���r0zƖ/���ǲ��t׍��	c�FZ|�#;a+�Q���I�!p50��e���hX*ҡ�s�Xϛ�^��d����|=k��B̶I�;��ǥCِ�5C�����>ơ\�BԸˌY�:%�<_T�EF�h�x�&�94��J���Ɖw��u�<Z_�V�;��ķ�;�9�ʍ-Z���0�'���< 4�
��Ӝl~���_`�>M5�ۊΉD<�V}?��:~Ţ��i���J���(4F���a����5�VZ������V�i}h/���R(�yz������vd?��Y�����t��jRS�N��]DX��4��n�~����=O�*���C[��$�"����}R�d���) lK����(?waZ��4nͩ��K���������-���P2����:fC�(�\Q<d��~Ul�&܏x M��;o��A�AL��z�(ԱO;¨$�@d9��P>l�w��e�ａ:(���%v�'սD�OF���&���F�`�\:ۛZ������ۚAu٢W�����Z��b��n)�&�4q5:G>l�!1�e>>3�@L�M��q�@kq�@NU�9��q�
ݻ��T�΢�>Q� ,� D��	��k n�Ũ�àob# R?%-��[N�'��Ҥ���!�*�u��߃�Hz�1ʕ���r�2�{�|��l/���o,}�|�5ѪΙ�hz���g����ub1(��8v�#P�k�i�ʐ��{�xa� (�k���v�B��Jb.�����Ո*G�q幧C�x��n�&���=w:���kW�b��%�E��ɴ{Y�����K!�����cHg^�J<�yo�o���nY��+��
�$�'W�����£�� �?I�싶T�!AX=G�ۈ7mN������t�!9�6�"D6|�A˔��H "�(0܋�7~-Q�Vʿ&�����%�RV��J��5U���{�Q�m\��$�E�;��*����T�*��C�",����q����-w�Q�Q{2.[=��J�a�y$��v���)q�~�:S�T6u,�T���{�����+��2�W��D�`$�>ܹ��`�7?�����y�K.5��ࠔh���˵��,������_IW/Z���(��Me2��<�������Уڤ4E|A�eU*SQUi9�`��s��i�6qT����r}��̫�(�(B�~�܋�}��ԟxl$�8<o����}ښ��#7�73�n�/�ә%�H�}�МG��2T=� 26MQ63�[I8���ё4M�Q#-��D����L����*3��݄z�$m�v�W��v�mBS�FZ����>I����U\�j��Í�$}33CC\�1���H��������|��7���ER�m�y2�����Q2��� Eb�K(jE��hW�S�@�� >;~1����ĩJ��fd#��NG��� �x%��>D JF"�4���p��|��*�՟���A�p1m�I�J�r��pU��D�B�����?����m0ɹ���Ę!;��~G��k�v���8��1wFm :���f���!�����Q�T�I��U�H���{.��֦nk'��.0m��#�AO����y�0��С��}�gq�Y���vj�v����,��.!���+��E�r2�*�7y�F�ă�*{���G�����kZ��چ��7�9k��k`�>�]��K�
�s/���K��wA�/sX�6��>���(z�8�~]9g}�Q[#�$���oюNb���+�N9�0��Qf���������?�ӄtézu���-o3�Bn�3T�`̽�te�������=���\�&I�
G{����W�/��R״6�tV��O��O-�r#FU'4���*?O�5!�Ώ7�Y�(����pS��'z��̏�k1�p�ɑ�K�o���I3�������� 
gf��$<Wr��M�����49�$��	)�����~It�2��3�{�)�vB7@�7s��c��a}�j�}�ct}��4m�VgV4�C���_=M���qͿ0�L�=e�V�YN�ϫ¤%��`[F�A�0�g5}Vg�D�W�����,]���ųg�ߖ���}��gND����%}�3��"<�e�b80LUƮ��HsێȒ0A��B�0�@����Piᮻ�N�:zj���u� �� ��<f)��I���n�þa�r��0Q�6��%F+��o���ى���.��h:����?��e0��o�OjV�e��5��ǜ��)W��)~��LM�S�F>B`��������pj|���TE'�<I�%8�F����-.ŁrhtM�bD�k�Ku���2nV��u�� ''Ck'�j�z���,��"����EB�u���{t����,���,�5��cN;X���÷ӟ^6VU7���!���d��CX��c���?�����=���6	ak�x!.����-
����0M�9o8�#��"[c]�K
9�.C	[UV\��e��"x!W�:TF������l�9*/���D�$�4�*��BDmP��	ߠ#��S��N�;$��4nĨ��A7DIi���ش����G]'��-�B��a�m���K1� Lb�bB�xz�~�8R4K]��=�3ť�Y/*�0M�Q��'F�{c\o�zbِρ�qU�s\�Pw 6\6���ھEou���(�wbZ],ձ�SN��F�hY�f����sy��e#>E���y<���k��z^D�~]F��e4�Q���V���<�y
6�����k�V�l\(u<ޮ||�Ky|=FLڏ����1�GKk�q65П#�,?~G�Ԩ�#�Qb�P�)
ŹzJ�� C��Z��{�k���;��H�8�6�񾧉7w�  %� J�p(ŶV`��p|e(��8J�������y�X�k�������֛滜�܄�v]Bu�VEU���dЃ�	﾿I���@�i|� o��燲��5ӈ�J]Jי`��F�0���?�K�B��R�4E�� ��1��k҂���0R�b�2c�-��|:�.�g~*�Hs��S�N3F�V�|IF���%�D�F?�ix�4��ye>�X�8��&�(6�}l0��>mǂ��k��2��܌v���jdx�=F��������D�֯*�5��d�}<��8;���oG�����=z�
���6��?4&J|����a�!Xȿ�� )�6q�9�{S��u�Y/?3��E�/�q��ɭ�tt�����&��W�E����
�".�e�E�( I@T�����H�*A@�� 9JΌ�䠒��$�9����n���Ͻ�TW���SUӓq�+�0����@���Ը��o���෷-�|��-���vO���>�԰�T�%:��q
�q^AQ�=c�m�}�]s���7�#w_���	y~����
ާ^�q�B����x��]�@\�9L�03+�*��n�����Zh�uw��;��N5�f�J���'�9�]�|�Q���rT�ɦ5+���wY�^ �U�߿=J�k��rW����͝���K��v.��t_8�s&��u������P�.D�8�t����{�����OS�^���y��_���S��}��7����?�^9z5^�E���Dة�|׍�.Y˛�W
��++�.:��2��A�د�ةg��lվ�n2�H稍��&	Ҧ}�3�vg�u(m}�@�����Ř��N`���Fc������n�/�ݨ�A��,��z
STb�m~���ዛ��r�7k^�v'H]��ɂ7кn0ts�E���5�Ǖ�qu�Kۑ������,��l�Vwk򡬂6��4ӯ�o4B|�j��'�#��v�g�'�v�v�ۊ�)U�%"Dc%�d?���~�Fu�!Z'���Y�i��������}�+���%����ŝ��s�z���ʎ�����3fu�y3ЋjR�p��>�PM��mZ|�Ӓ~�G4��s��/}�XB\9��?�\�9��!�hy��gk��/p؇d_��]_��)�ZB�&���#Z�\�dZD�iKύ ���}0���T�E���Mk;D��D�_nw�������s��mY2�/<o<h��� �c0e<��h�M�FJ$�n}��h1�����(/x�i��!Fi�:�����l]%pcPDO�m�H���WH
��?X�.�����_�ig�����}kR�[�
�� /��y8��E��l��4+��w�M;�x#�f(wluaa�J�.�dbxn��4�����2z${%���������8q�����d�*����O�5���n�;�O_|�{|L(�X/��`(��b�ͪ��j{�T�L�'�1S��EE��Y�y���l7Jn�	��˭�k���OA�t(�>V�/SCS׈4�����q�7��,��B��6���I�Ш4�=���.+�T3��ZE�C��?Y6)t'FAL����uDf���W��R��=�S���M����tf �S�ЎsRV�SVR���C��A蒇M�%h�S�ZO|Q��í�e���'����@��p�ֱj���cb��ַ˭ϟl��2����h֗�;#-R��#���P���� H�e��1��ц����׭5�ow��	ʏ>w��u5�� �ho/9���ZJh35^�܏���+�)7]}���;��o����:��)h�M�c��d��h�Gtv�[��vT:��&�5�/��0�^td1{���N�f��)Q>��ҜMn����ֺJ�h�����8�W��x'cS�J)��J�v���eNA[- �4j��E���v�ւ���`'x����W��_�n�ܠU-0��Qc[���Ug���  �/H�tz9�G
�9]m�t�}��`U�뱐�~Ӻ*�f���.<;�`�������]d�X4u�=2$���2|�K`���J�;��9`_��VdZ�i�޷��J(f�nN%;H�&e���NaS����|�")�ՠƟ4��T�;X9<�u�O��R�u��/������Uϓ?_��:�p�Xp��[�W�^�acػ�X�]V��~1�o�5�y�����w�}�f��b�^����Ph�y��Ь��>;�^^f��ҫ緐�?
C���{];"Iɐ�xiQ3�8@�s���ûo��j�.x�m惥��y�}��:[=�CL��Or���8�,gz�%5����bp�!h�<������X�
kS%��V��<K�Y��c�u���;������O��]x����Cjw�+�K	�D���/�QA<��}X�Q`"���c^C��Ә���5U��3+g�G,���f<U��+rn뗔݃�МU򪕡s��^�v#,#J��׏#"�4��[#`L���+u}�f��$a�<�a��w��,a� �@ET4s�e���*@hj�
@h�M�O�l��zZC�)l�;�TӶ�^�,hz� ���㫡�j�=�^:��^*<{
������1�u] ��%�f�������op�X�7M����a�ir`����^�ʇgqm�w/n*��Y�!�N�6�d����d��@�2�!C�0R(�q��t�K@I��Ϛ��h!�n�r;1��b��	*�1E�������T��o[���A��ޠ��u���2��ܑ�����Z~�hH:^9º
3�u�,E��h^vO9R�Jn��c��?��o���H![����֛RGO�[��oJg�����oBG��>�ߨ��0�3x����k�xj�N{���r�@�-�aT�b[��r`�'���ٸ/�s H��oN:��kE *=�~dՑy
��x]Tp��gx��Gr-яo<��_,q�T�����,�V��7�%7^�ƶM�KknVAd�f��1(��l��~b�6L��C+&��c�	�j.b��7�!��|��)3J�@�T��d�LAJ<=�����Dd�T�w^^����󦼒K���g/<w4jS�$t����9ǘ���$�݀vZ]&ds�(�4���?\˅5��=t|�Y�3�5����u�qA�P�Q�6�~QH�30=������1���m��_r�ǟ6 *x����~�>ߓ�]0u��ZVa����IUN�+�U3�
�'?:F|||���sX�ΐ#٦�v	����p#$U89��r��a̙騅����2䲫`u�F�_�Aߒ����<�X����[Y�}P9�_iL�$3kDk�RH�A����>p/}�!
ȸ�&�΍�E������w�@>G��GVZ�Y{��V��ޥ���_�i��,�Q}ݧ+���44@Y=�۰�z�V��>�����k��##Ҧ*���}�v%Q��K�5�ZxM���������x ��wB��p�v��"z���
^dH�
��`j�t�v7T��'��甪��t;;m3�H�Q@�Ă�4Rm)�~�<&��?R���ӽU�� ��������a�P��o��4��Ӕ`Q;����c���8`�G	���@M7!����3 L	2̓V}�h�۬��V%��<���7ch)�e����8S�βֆ��
�Z��	1x����WW�� ��
Zz��\4Ҍu%t���.甼�K��Ѥ�/n0���(�^�N�2D~��M3�q��,y�)�c:n���F�6���eN� ��p�8-�I�-i=qWX�	
Z����z[�A�����r3��O��
`�c�a�\�~�h�C�2�/'�.�NX���9'V'+�K����.�v�X>!3�2j�dp8��`����B��P��,J���f
[Y�L#�ᢰ�`Xv"�:�c5 ��e����>��w�0Z��|ei�E�`O��qT���u��"_]�=ZM�.�ذ�2��\�`�^�ྎ�Gf���7��l�o�M4�� ȴi
�z	��t����|����ަ~�vWWCNtC�N[���{�U��	��[�
^��\���a���G��K�㟸�a�D��W��~���xo��@P�#�RQ�|R�#�n,g���0���\���ԬNl��,A�z�k�޽,-��,�/.��h|y�M*�
հ�a-�-�쓻`�^�,���;�8/WP���(As2�Aq+�[A���^��&�|� :��x�Ī�Gº��{e.�`�0�݂��z�A��<[��M�Z�`M�G�.XzGڊ>
�c�����K%�$Ô��vf/�����?�y������Ѿ���X9R1~Wx�j�p�M>�13����|��՗��Pv�K˪ǰ����j�ӈ�u�;'l�K+Ҷ����d)�$=Q��k�y �~S�a�_��"'*�m(|8�/�V+�l�������4C��h�7�Э�y������odےZfkA\����wH/t)����6��I=��vp� ���:P|;�0�.,�݉f�uXﺸ_�J���q�MgQ��i���:Пv����L�I�f�^�r��G�|f[X�w��n���H������D2��o�q���8j%�֤%63%=6�v�;���2����|�כ&��x�&�||n#&�K_(	��|�y�+��?��5"΢=F��?:�ef}�4s�ygvH�3p���|���h�Z�����s�?��N�z���QЪ��K0j�/����r��G�<f��]'iAւ_}�|×>GA�u�1h������/�U���V���H}�)���7����:��tƇ�$��n6��
����.C��cXtޅ
�f�H���h˚j�7Ո6纏��j2ɯ��j�T������3�V�ċ�U��#MP������֣�S��U��[��k[��P�8��V�Z�G��7t�E�ʗ>J�~�pd*x�CDT=�Ѳh>�����Bz[�D>7�ʇ���
y-���Ϩ�C�;�5����`G �c�`���A��������
W�B��6���=�Ǻj��S{瑭��폳��������D��#l'^$���*ϙ�1iAM�
:��3ɹ�S.�l!��V�W�� 'i��dD�w�*p}�c���Aj}�q�?���V!�!O�i�S���f��	���I�&{>0�g��U{������[v�aZ?��ƈg6��W$fN�H.����]�:�23M*hެz�#��ْ�V�G�����ں,4U��!W��s\��ô@sߟW7�����GV�=��m�t(OC~�D�i����"���c�G�VfI�$7*�g �UG����e �_���Hi�ɠX�P��=[7P�Z�&������:�� ��!�&~���'�F�j~�f���r-�3���g���<�Z!!��}v�ģ|����L�j�y$�T1V�i;P|��u�*<��-��-���<K6�J�֛u�hu�|`���
'��lפ� ��.�����K-��+;��IE�hN!��\��<�=m<������x�Bc�j��V��}HDi�ؑހ��7��3r+r�T�#�5Iw�Om�XY��!9�ܒ��L
��=� NQ�K��Ȫ�V��ֆ��.XM���Tz��.v��"�׿VL�e/���}<���qH���kH��`�g�]�d�����Ԧv�c/ë�֌�q*��{1o�`帖j���E�-s8�k���"��Ú�{�a��>������k}I3��aLe��k����������G��S���?��̤Tn�+n��l!��=t��(*M��'G��ۜ���|7%�"p�Rrm=������]����y�k�z��6/6�h�q�$|˒�]��v;.hk�os*�a�K(�	��oM��� �	}
^�w'U��̀�dA+�$f8?w?��%O\h/k��#�����Ҋ!�#[M�pX�6����&O�%̴�X�8���Y��ϵ��rM&PW���c�~�ȇ�:�A�`<L�=���P39F�qU𘛆�=�c[�0l�Cv�ap�_�$��H�����5�L��  H���"v��Y�V)b�xi%湺��x��d0t��Y0g��2��kcյQ@����Cߘ=�fa[�X���(�h>���%n��>*���:����Z9G��z�=;(vB��@��W�Bi��ʥ�R%
�;@VNU\�3��߭u|יdI.��6�6�h8솽���(�R�#��5Q�l5�y�w`�,�#��������s���X��c9x�Z����=�Ѻ�RG��m����SJB��aj�4��k�v��U�u�D���(���&����j��P��R��?X�	ܪ�@����N�w:��ܧV�������$�9�6#�Ɔc6@M��:5�q/�1A`Kq��>w`������!� UV��c�)��a���k@�C��&��U���!X�X'A��#h+dM�����|�����m� ��^+�V�yI~��
��ɲm�#�����S�M�*��Ӭ{�a'h�����{_!7[��3#�l�I�ؙ�A9Cq��[q٪�)}�8h�^�EIDHVV�;������췪NnXT��o��D�R��]�U��bG�#�z�&�C��|Pb�8�[��M�8@�ix���ۍ�݋��&Jpu��J��T�蘵S-����d�7es��N,��jK"?5��|\�!�
3�z���~��gL�P�EcP�>\!b��MYD��ph`n:���tN�w�,;4�����o9�k�S^�}\���E��l�[v�gE�oϚA�ʪ9��g~0[ëbF��]ѻ.���S+0}�Pn&�JF��� ���!�!�C+%�A=��k� `l�}�I�4{�T Z��}d��k-J����5{:,�#}�$E'y����Ǟ��/8��C$퍬����;n�>h٢(i�
�i|n K㐡�s@Tvjn��V;�qplG��áC��cIu��	�g��2��|����\>�$PG�-N4gQ���XD��<Ą���ʎ�Ab��%t��Y���h��YЀ����%v�ʹA���7����\��f�<���� `� VS	}Ֆ����~l<�b��ADD3v�j�j�V�� ��p�f��n{~됡Ҥ�̱��79\\���#�1���$E�xiS�v1��pͯ<�,�X�Wt�����HFQDM6�K*K�c�4�c��l� m�Ϛ������I+t�o��ʶ����܉��L/^�ݲ�=Q\��"H}&��E�+�Ӛ&H �M�;�]��UmĠ��9�����>�:��
�՟��$��|]J�o1RG"S���u���^��|��V�Vv鞙o��	NC]�0y�w|�^H	'-�q��C R�wE�՚���E䔠;k�&t�4xxw�������� ����Yv'~.O�#4��Z��<&J���j`�˖h<H&����R\�%�g�n/t̚��ȍ+��gy%I���@�H�|P��^�+FX�`<Ϧ���Pn���Hv�4 �W���h#̢�+˽4#aih�*R���ZU%j�&��w)A~�S��<�pw����A�#��+g˓$��3䠡@�g�{�&���'�j<6ж�2}Ը�����b�y/}�mh�ݡ�0��`�<6���Jjj��?L����)�!�%z?��^Q�������W�U�M�ʹt�3pޛ�S��̌�������0�,����_6�d~
��ϛ�d"G�C��x�����`���*��D��)d�����^n���c�0Q�Ȧk�;\�0�]g������u��̖����c�S�������`'�m�(�yi��լ���ÍY1�4�� �o�	��`�2#�Q�:��M���<�~A�)��/ESb��X�5s ��Kj�I'���s(��#��"k�%C{��PR�B��^ڌ-[����s��� Q���GG��+v�Vɇ'Gn�à�γ��ؐEf�����4��7��}k~3#�ަ�ޝ��}G������aG���OCV�)h{�;d�9Y��ڎD���y��5;�~�k�!�����t��`�KN��k��9fKT@%�ύ|����������86u�I��Gv�!Z�!9XjˮH=?����@E�����j�ƾ����|�=�`^�4eA
��BO��')ߋ�f`�pX��^�3�jy����5����$@��uy�K��j9iA(WqN��|���t|��CG.�Xvk�Ճ�b�Ƒ�w��x4�gl��Yt1-	��ٗ Y�i�*��%OU���߽�߫ۜ����E����p�L�c�%>�kdB��W<c��4�cu�Ҝ!:��e&⤫�CxVI�8E���T]+c��pXOJ�c�w.�)0j��6��4��
�'Dk+p�M����6���dp���F:=�
:qY�=Z��ԪuP�Z{�H��f-%�����fs���w҇��x��2O	����l�oq�i�^�G����C�!<wA�;�yX�Jn����)����p �����S �����=JH����P��jq_t�]+��\�nTv��,�@������O˭�9ORk�4$�,���4C�(���3���[���0�վ���H�r]2y�Z*����;�a5���T������ݞ�_����%z��`M�G7 �Wf�P����er��[�p�[@����_f�,7J�`vV:�����m��9#�W���/���YZ�+��������m2$2]V��W�'�vʗn'�ykKq��@�w\݁J��Ϗ�m�5���
d[A�w��piz5ʼ<���e	Ād�Q9�k�������γ�;ѳБ�᫢�Se���N�F��^�D6{�
�rǖ�L���OV��
nq��e��0Γm�G
Ι:�3�H�>�knrGO���WC�6	JƆm�\�F.	>ܑ�XJڙ��Wp�H[��_�>;3(��ݰ�CB��<�A�l@�76
�wǪ]]����A\Iok�Ƈ$ᆝ��?Y�t(�uS\�����\�	�Sn�'hb�M<������^K�uA�9�˚�R�ӿ��~*Qh������K
_Cy�B���Q����m2�.I��?���g��I���3~��y!����_�;��x*/�SՖ�z�n[}�y�#1"EC�i�Es#e��uh�F���-���.Jz;���p[��2|bk�(�^w�.J����v׊N���p�%�H���JՍ2�<�B�u��&�I}��5Re����hPb�X�N���Ty�Թ��#�[R9p�k-ēUFu�Ҽu1�T��i^l;X�����E�:�^T�.�P��։Iѡ\ޜkd�/�G�Ə���%�ts����?���Ks��m�\�xz����&����!aQ�^k8p�@ʨ�Nc2}�Nf�����u��|;�6Y��z�2��;d�v;[�"���Yі	��VK[���7)L�����D��ų�a��x;e6\�?�١����@��H � ��3e�͆I-���]��O�H&�MZ����V������/\�����ɍ'����o��́�~�����1S+���1�7g�K5�d������.!]�ߚ��}�k��Y��J:j�W����&���=x��\b�s[K��F#�6����;m�6ڳ�$)��й�X�#��Wp��f���t�\��	�yh�Q��e}�yv>uZ-Cw)����-\�n�q(�od[-/ufo �M��)������'���2���gsr�wN
_�^pKF^;�y���V[Y���~�y#=�/��k��Xg8�&a�Ŝ�?�K8����ĭ�և����<,��<���;u��1N�N�����s�E\�Z��>��Pi]3T	M�91�"h����Hd;�c4���>>C6���7�K0z~B1�U�R%-w����r��[�PUmE�Q�lC�MRg?�mt����{��\-�1vh1��[�Ha�?Ś�Ί�GG�.C�W�:jpH�#/_h��E���b}��_KM�ߤK�P�x�h��CB��\c�� �g�UrU)����e�8�ly�գ���Y�AU�����Uq�%+.��*몔t�+���rFx+ �1='1#"�6�!�/�#\>I�?ozģ�U�|Rv�YC��߬G�WXR�_���u�Hz�Z�
�X�h�{P5�U�ĦڈK��\�6f?�p��vp��u���{��8%��*-���~gi�J�m30f+@u��!���
W���u��ا�;�%�z�ǻuI�;
Ъ���xiJO�u�9b��]�a�òev!~�֥�ó[��*�Qy��j*�oe�밉��Yz,	�^�ͼ���߮l�`��<�5n��u0��q��r�XZٞp����~fmIF�/��^�n�y�*Y���El�)��,#O���ޜU�>��r_�{b?g�-�Q>́��6I����k�bu�F���*��ׅ�?�xW 6��ګ1��
N∢R��I��+���)Z��>?".Ñ*������G<C��{Ҹ*������%;K��IP��L>S̨�	�d� �a�/F��"�[�ӕٍT�2ˢ@�o?��%�u��c�^�񗞲�zOlĔ��[�|ccGh=�㧝bP2	�6�F\��)��>ҿ�M'Ҕ�2%��)��=����}�3�G&!�9f�]�a88;���-��B�������pp�:^�5Y0����v���aS�P�w�!��([p�Ύ��H[����w��8q8.5��?���S��X.�:�n��y��}��H�u4"�ɴŰ�bP�̠�J�^�[��)E�׉��`
���4�e�,�~;�M*��*�D��qO���5�!R����a��qeb�R�+���.%wq�g;!oiC�ۤ�6{GǠw �(�Y���f�~�������E=�p���c�m��ۈ���ד���9"�5c��Ha$���rpi��7\�x��t�ߞ�ۑ�V�s��6�6�b��k���;��N"�����L�$z�2E6KHwO���Zґ�j��N5��U:nq��z������la����U�K��!�rq��7�p���tS���Ti2��J7~�85U��H]N�'|Te����T��γ�r`Q(Os$G�����qi�LK{}��|����a�L-"�l�������������xڳ�fY9 :��Yv�f)�QB�F����+_�g�\�RP�
Иmh����CB2y���|�!Y�)��KQ̎7���Z���ZmzFN����k��}p��"�M����1�� ��T�C���/�!� K�ێ&�
��RWĕ���
f��{zEC�C��֨��j~�{�c��Mvވ�@�\̠��咰�*/��/��FE�lq
f���������ٖ�~YN�����WD�������jr��M38��j������?�e���z�"�
���cSƿ�r�3\J_����7x��
@�R)���A�9d��o��֝t��AiV@=H8^��/�Xf�(�tG��x�&�r~��8o�Ӆ������_E���'��;�}�i���MԖOM65Y�~2� O�\�84��u��sC�(d-R��gy	K/���~9#8M6	b%iP��)�����>��(8;��^d�T�UJ>E�;�[X����I`�W܊�0���3Q)��B�v����ld%z%�*�1�A�R�#�6�[T��:�0/[⃔m�qb1dMY�Y*��k���l���g�������v؄���Y��G�o5�h�+~L�G�'(��u�-��^=��B��"�R�Fl2i+�_
tts��:�s�y��1�?��o
�fgޚ�^��D:�4�˞`���p�뵃�KoM��60Ӈ�A3`�b��>�p����J.�+��Q�2���a�;�7��c�%"#kD8Y&R=T�#}��X1�$�nw��TI9�w��uM�-I��0;�4�B��.|+�Q�?dT`���Z��x�A�P�<p�3���F��1yr�1I9�Fr)��#0�N%t���_� ��J޲�!�B {A �r|��N[�kAA�� ��R..6�Lt�C$ �[;r�;�%M\�s�-PΙ��YS�%�+�0��'��s� �Hn��%�ft}��pȾ�����H���b*sSr��'�C�Zݻ'��0��l"ˏ/�|�eqW��8A^UlLh#���	���Jq���' ��+֐��m������Wl�HJD�+۲�TZ{ܨjS��5��h)�88���V1�?��B���'~���ɍA1hpV0���S�ho`;ڈ\��'^b7A�΅���M1���^���,��J��%D1C��*�g��/q�NN:M2zQc5�r�`�<��=�'_
��SX$p"�7�#	f#��(Ys����#Fp�6��:���5��M���
�3|_��W�S�1���BSн�;��+	+-�Hz�}�*�8?y�Q玖3����R�5Cyi�D��!���ն�Z��Ԟ���{�Z#�dq�u �����Ր������<��� �o�R�>RJI����+��i�E��d��V�4�m�����o!�7�"�ر��ˎ��+T�|K���H7�V9�k�%�:!�v^�����xQ��XŌ��\m�d��*�,������}�?������V����-4��	0�U�H\�.#�S&cn�@�v{v�o��)�S��s��k���B����m�=�\QG������W�il*F3���� 6F���xh�Qe��l���ь8�HJΙ�I�s�"�ܐՅ�߳�w�fX�?�ͥ3�c9K��ݚ_�ڙ�p��A(���qA�d�=2�rC��[�%6+��'��h�2�'����Cs�ĸ7�N+D�
��h�Zm���O ��F�˕�b�5m�7�ۏ~���Z�߈���.�x�x]Z��S�Қ[Te.����(RR	i{������aɪ6�Nd�E)i�R�&�VP<n�wd�:�����4g��{��{l�ς-b�u�_�\��R���r�֤2�$�")'�Fpoρ�]�͕CU�y*�b6Iˌ(�޲�Z;#�+�[i��K��|���X�e}���%/U�@ 9._�N�cWS�b������aA lsѩ�����Ǔ���xࢎy*���.{��	���!�m׺��nP�����Fy��+3��3d���Fmr��xz��yz�x�9ϖ�q.:�q����O	 {�?"h��f�����V{�V�0��S��~Do�?�>��pf�yF_��ףM�(g]X��P� ��2��%uZ��=�Uu��n�-�=?��'�\T�1�a#��sM>��6H�z-�>�ͿG���P�tw.YbӘ����T�9:�^)eRO�{8��~�y?4H�E��WX����VV��A��Ε�'�����=C6�F��
� �d�j����]%�~��-�1�������#èE]����Z�q��q[_��v�����SKM�Pm�5�zZ�j�����Sv�F���9U?��a=B�o��g��!ݺGzWg�� (�SM{u��k~��&s�bu ��OA�ow'���욭7J鼦��m@�J��>bM;�����8%��؏�h����*�X�8�j��T�uR`�bu�G/L}`��|~�S��R&��г7y�ܡ@��(��0w�[��%��Ɵ��vf$jH�b�%'�,2�W$��44_R�CFԉ��|n�Vy�@Z��
~ъt5�֜#�d@�{ŵ,�
��4�8hqX�OTv�q�rƟc|��W�HCU�h��'���Z�Ј�AQ3-�����~��wF6Ih�QB�O���Z5.W�J�eKOUq���%�)oT�pB��*�pŕ��,�8h�/��	��=b�j#�"Qn��;)п��Z��~�\��Q�K�n�U�L�A	�R�
�:��!B�>t�ދ�.A�7��ȫ%���8.p�`
�{�4B��{�5Z��3dּpń��L-�.2x�P�S���q���f��_S�iځأ�v �A�h�@�bhm�Ju��������w�E�pE8_��^����%JP@�[i�k��~"A"A�eǞ	���H��.F�n��b+��#�� s�ˇ��ࠐ�W)&}��z�Ҍ��Ҏ�a����!3��d�؛#�oP@�$��:wc��ܦ�:����Q���!PTP�lT��"�?��݉*��m����"�n��0q�M��c�ه~ȡ?�h��⦾�8�m�p��UX+��S�?������"m��t�6��{��Y�_�=�̮ߜst��P�!^�x��L���;U���������1GȓB J�*r�ða�ӯ'�SU����P�l�C�6Q:����� E+?��b�6T�+Hͧ�f*�MڠyAjEE�E ��UAE~o����㭠�g�>hb豓��]�	S�� ������N#"�:�����3�V���et������'��d"L)�TJ�NB������j73���
㻑��	�B�/����1��~0ⱽ�-�#ѽ& �s%�r�B_@�����?��,˂��V������BۜȐ���	i����gU��ʵ��؈�h@�x�����7ȯk�ǡ�
��z��_���1��՝���u����+$hU)f���|n;2mY����[`�]L3�@�?mU�%�C|4 |,��S�k��Q�l�U�NP��E����P���z������Ϭ:,{��C��F��o�H�e�0��T�D��&���q�@��T��#��Nn��� ���%�h����OW�I����~�#�W.�Ӄ�q0�GDƜ�R�8�#Ÿ���+te<peɽ�1|�g�j�,C�/��6���G^2Wl?�����ϡ�X�W����h�kw��u	�{���%w���M3R�
9�9����;�V�L���+C6����g������/�5�SCB@���\��,�|`UƔ%(г-o+bl����L��O� S����=��6��`�jëeK|*��l�D�u�{9�0Z!V��ݲi8���T���	*� ���͉� ^fZ0B����ʅ�	Ј}��2�;��-�Bn��lu� G�V�.�E�j�"���ƕ��L|U�t�_ѥ.�̰�*:��[P��m�E��ĖĈ������V/@�7�#ı��̃X�8/��#�nhN%ץ�dl)~�05�f�g@��j�	�����!\�ʎ��.vk�"M ��JH>O�}b�y�"��������!!�eT�>����L��x�i��3a���X]_[om����uE�� ��j�2��B\Va����P$ >�`P�O�����3�g��fsCTڗ��!f7m��H�?��ߵ��G߹��R��B7���_-�?1(��Ȑ�3�`ۊ����m+��e- 0��π5�by��<	b�����ܣ�Ou-��~��|/�MY����F�B�!��Ȉ[S4l�h�h�a�y[SS5F ��[m��-67� ������x������ݣ4S��.2S��qP6<f���o؀.�(`���4h�޳ 1�ԭ/X�G��z�k̍��Z#`��F8�;e�S���%Q�Z�rK'���- ��Zܙ��,QE���Y��W���aN��{��
�`p�̻�KU�^@�@U��mc�����ݿ�gj�e1��� ]� ��:U����.\eW����s�<u�t��4N�Ha\���*�KY�*sw�4J�#�e���=��3�����?�Z��(���ݧ���$)���9D�%���yt�N����W��=Q�dd.n[�t�p�V-�Xu��>�S������-n�!���x,�m�Q����Q�"tC���) ������)��h��[\:�wu��1\8:J��}���=�y3����I�0Zu0[��8|�G�$Ֆ��5W�B��bj%ܺtXMH��S����m/�*����YhMk�KO�����pe�[S4��zB]&�O3i�,��Ok�����4aM�x�#��`�����
<76;����p��K�U&f��\M�"U�|��з����;ɸ���+����X3�ʣ���1K7q4�~pE�є!���U�A�-Γ1iD��cm���h>J��=	.�l�b��*~��˃&ߩZ>UmÎ���%Or9%������*�����_�D��CK�A-����U����!��f��aL����˽O�UA�z8�&�P���ϯpd�Î}N��(`C1b���p10\�;�u�9���?#7�����2���a�RD�\�(�ވ3��y�c&>�Sz�p��O�V����n�8�ޤN�"�
��B�Xe�'Ǚ�3� j�j%kw�/�v��G�\�(�aI�����u�XE]n.j��Q<OW�\�˥�b�������P���a�����أ����mQ��ә��ع��#;��l�LN�]�)��ZΡ��ǿw61�|,U����1$컦B��ッ�s}V����&ͤY�FN<@���o�Rp�Y3h���	/ٚF��@<)�т���D�0��&+��χ����aW"V���+Ή?w����c{'K��L�����B���H	[�t�$�t�D	pm�8�%��]�߮��+W��mo���M��8�SZt�3���̠Fd
���?��Ҷ��S�ԣ��<��"BHHН=12J��.��V3�Y�n���?`�$�s�{n�y׻%�Oc�)>�*�<�\���~�!�p���w�z-���Y�~��=mf�p��ċ�ʏ;\���_:��"&�5l�i�9�A��(-X�e�He�$α������2h,�U�nʸ���(󨇥�>��5�0g�ܿ&���C:/nW,��W��5�ehЯ�C���3���t�����x҉���0�f�a]g�ց� �0��G������X�����Iyx}���Y{s̔�����犻�pX7r�'�aU^�Ē�������UM9�((���e�II��U�>�o�/���
h~�<��񳦮���7̷�$I����eУ�Z�-�'P�$`��0=���a-��q����3�G �Β�]~Wyi���x���4��X����1��JSH�4�(�f{$f���'���E�Hm. �����p@�i��?*�#�Uq��\8e�xo�����ar�$�K�G��p�h���]I{1v��T��XA�'h׊�ēE���6:��8�H�j�����"��4[]�	��Ұ����Ui]�q3`a��j����@��̞����[��N2 �'���˞���\('�O�"�����~=��>f7���>�`���pS1&c���ՕÕL�-d���Z�^���E�3��w:I;ے�]0�@�7�+�N�
�;r�@c`n�޷�Ѭ�;[�n���v4���_qÈ2��7�]$��e��t+OIZC�A�@�oE���N~��
�pқ�	gpK#.�&[��C�*Vop8�x�P�@��e
���g6�oe�3	�G�����s�hV�t��/aO����p�E��+s~��ľ���\�~�����S'�mVlk��� L����̹��wml)�ZF�I�����!ʶ�#��?�2Z����/
�w�||j;ȉ����'��].!�_]���-~��$�ϴ�I�Ǹ8�?��ߐݐ!G����̴M6}����RQ+ �|�d��/�K�-l���Yo��'�z�w�3:�a�ޜ���2�˖�������P��Ԕ��l�;��T��	�.���F��,i��xY�Ld��S� �}����J�-5��;����Ko�%��U}_#�����'�fm!�ds�K�P�}�b)A��g4�^�)Hvs9�MZ+�0�����p�*�����B����~�X�[�;e��ʡ��G��#`�8�5��AyIz�x�YIj11��`�֋���eYt��RWU9��I��/�@�pX�$������J�|P]=��?�6߽A���P"���G��ey�	,W�= R8F~���� ��y������Ǟ2"f��m�X�#F�ڽ��Q�ꣴ��[(�vݩ3�1��nc�Kzv�$1e�( �a�X�w�2�^��\��$s_�g^胢֐�~"ހ�S����aW�
y+� |]���%{T���h_x��x'��{�¡���a�/���{N�����c-�{	S��yW|`����$�)����5��`��<�f��}y�/NEU�]!G��3�~qF�D�h��O&�#��i�	���Ͷ"%C� .��4��{Z�pC��o�����k��� ;8
!(�;s}�&s�����a���S	r/]�Q�j��4M]]|��XT�?\�o]ue����؀>���JY���� ��"���PЮvi*�a�=�_�L��>�#bI��Q'
�,�|�yB������PQ��s��#�+E����*fM�d媚��tS�<��HH.������Ćy��$~ڸ	J*����Pƿ�2�̽�q7N���\~E^ޭVe����% �\bt�@R�]�,qϻ��i����a������a2�5� Rd�(Z���Zx�b�p�>��m���7I���C�����\��p[�$�@�����&g`���x֤��0�ܭ�	Q��̮��cS7hQ[������K_(ퟱ�$ƈ{|n?�$�M�;���	& �d��\c��_�>����\?�;#~�f��	�e 0YwT�^�ۗLCxn!A��#�3s����O֝�#F��2�M�>���ajʽ'���,; �e��-�}z\�,'.�ZPlh�~P��bx�. �oS��m�R����A���L'CrD�t"���{E�����R�s<�Mxp�����Ed�!���������D��蝵���$�5e?�g\}������"�/�H�,P�:9�{n�w�_Xu{��#q�,����<�����u�P����ఆ?s�p�/	��Xº�Q��ѩ�IG��編�\`��}fh�E��/A�"DV'�Y!ｭ�
yt�@<+���D[�qcd�'�"�I�n	9��oV��W�ЗJ�}��@��2s����l�G�i.�笓xW@�`�vc�}�biU|�K�/N ��j�����>Z:�����?�PI��:B�*�<��M�؇�'��,~>/�����
������&��<�٬Q�ܭ7�%h
�u·od�� +:�̋
a���,j �'B�{�ϑ��BQ,����v)�� � �^ �~��lİ���Vf��-J~A����L]u@T��vX0 �DRR�t¡$�K�Nghp�I���J�J9JI+ �R�1���	�?��}���|���n����Rʺ�B���a]`d�9W�l�9����-�qr��DQG���_~�oXx��(c��%ٗ,BӢ�vP�� �/�f�a�#��h=���#>7�|�>�l�/D���{KvP����L
�RI��[d���bo���U�D~e.��Zwy؞�{�A�����;H�H:N�؝� ��-Y��62Ia��Qu���ٜ�t'�)�	���S?Q/b<���T��WV`����_�L�U�m�r�4�˕ %��<<3֩�K�w+g�s�Q�?A~
�~j��؂��&!X��.n̘��ӿ�X�9q�m�� 	������Q�W6�l�H����w��jNk�QO�h�PXe(B���/V��B����P&���Ax���{�*(������s���������!g`�S��q��s���%1¯'�	a_,8�Hm����"4�Y߷-m;/�����R�������C��y.�D���Y�?�E����P�؂����|*2g~j�2b����)�P�m[�t�0DFE�';a�����U00���o�9�a�M\�YS�&�-�C���Dq^~�/�vp��!%䍬����C(#ť��3C5@c�;������KDo�,9��%�_����Im�E �/�1%��-W���|�a����vh��~y\�U,���|�k�E��ge�R�D�Ll�;�5�j��֭�>��0��-�����:}?!]�X����e���6� �Oӌ���+�?3���C�ߞ��S��3�J`�z��D���z�?�L�L/��-�$��^͌[�/��c0�Y�U	f�	�/��o��bo;/o(���D��+�Fj�OR��0����c��*?��f����� �Q9b�\�C1��l��wz�f4���!0�QN�j*�:�s���"̤��S헛SR:��9��}Z�&��bA�i�$��m�W�4��q�VޡKꖗ@�]�F����������Ì�N	X�w��cCܠ���τk:��8�5TTOgf21n*]
��7��6��V9�BUM_�t��kG���>��RX9�8�Q�Usv���[�Ч8s��i0���A�:�~��߲��B<�[�g�Ys�O!W�Z�� !�/�
)P��A\C.mO���fec�3�ÿ$��2����Rj1�&�u<� ���R�&��	3�iĖ*��p�� M.��)K{����ɴ�M��p�?L������+On�����ު
���t�;�A>wД����"�@�/'W��*�����h$�{؟V���$�gc�~������"�Tf��b6�|�,��@�'y�����V�+8�u`�C`߃0O8Y2,�U��"`����ŗ�>_֍�Dt?
$��v�"�/��oA��&
f_�8��H<�ޝ�fq��j���U`��F_�Z�i־T5����wP�S���/�O��ւ��a�~�1�R�����˺^��=�կs9$#r��_�@t�W3n�J��̏�����g__8��t��{~&&��"ࣗ��O��6�)W?�P��\���G���G�ɑ;��
��?n�ɱ��p֛(J~so�S��vn�9�
8��!'��!=�Hz�*B�n�jt�*pΏ�'Y�9a*)A�o��u	oPoh�a���"��KT�;�x�=v� ���X����9�cf͌,5$�������K���/~�O�SL�|��]�	��	O�[_�xs��\37�(hH��܁�vv�@�����p���W���7 ��9"����FO�Tn^�[�m���~���N���'�,.Uq�1v���u���;M�Ф7�l8�ʨi���A���7`!q6G2�%�4G�6qW�m����~���R@$�=ZZ�Դ_�Z�<�.鸀� 
L�y8vX1����<q���Nz#羏��da&)�~�&��O���{.}l	�WaFP	��p������iPM��C%�O`�p���n_�[Ҍ�$x|��Y�uj��bm���ė:&��g� ty=$<��S�LlnB^��&2��Oc3��������t�_�]H�D`0QY���gc��ܺ���́� �X����$8l;C���@3����
Ǻ���Ӽ�4~�ơ1*%W��YR� S�������3e�����4B���o-�O5���
R�.9^	���5N	��M�~���WYW��|��c0V̚vi���$v���#�M|��Lv���7�X'ر�ڂ��s- @��]��~F��N4���W���0�IY|`���O�m� ɾ��\`�M�`l ���`G
�[u��+�B3�q͌ǥ�g�r{���EL9�&���K�F�rr?+mKmC�(�OgKjAH�\�5�>�D���$NJ��]3
�6i�6�mA4.ǟOs�q�&*��ۀ<^q�>�yJ �;ks�b7Wx�p�� ��/�М0@��@���$%t����uzv��7<�R_(�+��H�Rf{2(x#�b]�rNKJq��W�D��a~����]+��!�Rc��\��}��`��X��b�Y50ޠl�D\��b�#��%6�|~�W�W�P�^
:�� (K���������_4��ȬK]�řH�1�1ߛ�<3:~:S���!^p�e���1�6��r�b�?��$�ucB�d#	��Ƴ��1�3��fu>���D"���wnճA>�d�d7(r��y��e���ݏ��Zy�oH����*�Siߐ_f�T�����?{Fw��D�,;�]Rm,E ����b�O�ϕ�,m	nঌ� �sx86�{� ���#.�-=ҩ�о�I�+��aﺤ�k{�����@�c���fu�a�?��P�en����jOpM��=���A&���m�I	@�a2������Wx�_�������`����g��	�U�_�IQ����,��P�'���r] ~��#!�։��[E��dn�?��IP�����_�����J15�ҳ}�OP�1��_�fr!J� a�Oi��ro�R�8|���y�O�&�������j���l�!����3��G��U���w�M#@�	���m�L�O=���)Yۜe�Hztu"-��>Ōq�m�)t�K�t 9�֖~�Õ�4���.7Y��)�Z�2�><�wm�v� �i蚍�7_m_XW��U|\Nx���9A��2�}�f��)$��?���X!���G|��������ng٠%�<�[���W�V�ߑ��^��)6�}�L[��
yYy���`6����"�[��
ӛ���O��5R��P� =�Dr�|��'6e��,߰�?�<�ݲ�~C�=+�N���_
��Z1#̓���_���(��.�Cϱ�^S:����G�Խ}8�q�-���!2(hq�̄�y���qi�@�S�Di���`����߿�x�K�p�8��}����OϿ�L�ކpp�i��2
ZR�]=zUwh�nnM��;Es/һ�4�
ή��p!>�䗻��"���w���R�,�A����~��i��No����S^�Z+f��I�C
�qT֘^^9���*�t	`[; '��s�g�hx��,u8t�9�0u���_���=p�}Ph��`����d�Z�jY]H\XuR�da�����#�u���ƥХ���������BЍO�����E�K�ߗY{���`���[G����eZe��S��%���y�-���&�,���ss�=��gC�!�ҭ�j��8�H��g����F�9�R��و�i	�<��g��h��oIIP~h]�B")�����b���1���I�b����s�}�2��b<��IV�;MBc��.��)s��с�\=S���b����́m;�)���'����u�������Z�c�I6�!1b�Z鶲��H$�J�ѯ�cV�eĶ��S�r`da#���-�v��$0��Xr�W�N��NIf.�:�̼�Xd����!{^��V.y{��6O|T �;��l^�,e��]g��1������n���y�����|��C���	�W��W�9�����U�b�����p��
����d���Њ��Ί"b��G�pq������n�3%�D��zMI�
cZ�H\�$��Չ��b��EͨS�	��5BYZ�Z�*u��U���2��ᴕ	���O{�i�S�h)�p0sCG�����𩍚q�9l�%C9�&n|sd�_��$�:+ځ�eo�D|I\JQe�&7|�Z��t�0	���0y��і�.� �=�}���LY�/xx�����{�A��Uj�\:5�w�V:(�x�LW���|�7�-d���{�/�Pu���$��6�b��b.d�C�ӣnb�U����}%�*�5���[�0Ã{��b��,޲�v~:`��a]��W�J�Kѵ-�0/ר>c=�a�(e��%���qӵ7�|���O�F/F���_A��L����P�ְ����XSM��13.�,��kJ�X�=�^�Ǵ�u��`]+�N�U��\5��{Ey�,n�=w<?�E2���JK��},{��;XW���xW�����x�����Ɔ��"���v8�,�^�(�ޅ�Α)٫V��tt�V���y]>�Ar$T�$l���V=�i�����1�|C,٩3^�������V彩X�0탦����?/E�GWs����v����+ޮ�t}P������a'n� �g�z��WPH�)G���ٯ\�c������ԧ��M�#�m�B�{{�Ge"����V&��\v��6n�H2�[TZk\;��Fd��G��祐���_y���,�Y0�M{{�k&���/N�,���Okq�۩u�q�����G_
V��$1fKu�J�4�˝9����QE-o���d�, ����
��OW�/7aQn7e��O=�ն}{'(HmQ"-�`����9�Y�H⛀m٥d��Ecg�l{����Cn���˸�a��'�.րxt���� ����3BB���h�w�VHa~��YD67�F�~:���}�Q���ۂ�#"�Lqsz����������Ci�����տY�;y����-��H[I��J��N�	��&����5�c;�S�ʝ&�C�d~N��҉M��C]���z����F��0yb�i����H���s��fZ�'��1ہ�����˔��[e'h8k������z2N�(?��!��`���<�Q�MS{���[���e]��o!3��I�����c7�!��G;.�� �*�������o�MzN���2筱ԇJ�2|-�<4v+���󟌚Ǔ�ͣ�<;���'+O/ϔ0�!_H�~̶�j��n�"��6�<,��J�L Ǯ�p��V�z�D*,`FeZu� *��F~���X�I1}9y���Q�D.�V�v3���zdb�i�����f��Aj���bw�H%������.A�1��ei�.�N�Z��/�6�4aI�`/�fwV6X졬	f�ae�"�6fJ�dE�dV%�o�;v��o����e�6��n�0�̠s�IVo#��N�z����V�mm�33ҥ���^�ܕYv�ϝ;�4hB|,��o�`�#��♙i+��*[��1���s���xo�9�%�{��5
sα�h�;�Egp�[?`� |�1��|}�HJ���?���w�J5<D��:���,�����2|2�� ҾQ�$}���H}oޖO���AP��%V�Ud[)���ze�S��?k��p��=t@էp���p�>b����	��9[�؇��o\��H�(L��}�d݊��o�#�!�sc�s�����i���r��~��%�%�4eK5�z��y�EV�k<%��P�]�k�>ǧ��3�% ��� ����Ǚc��Ŷ
�	��z��M����3�� ���D���n���\)p?0\���b"���:j�_�����v7j����?5����#6k����N�z��������Ԑ�<��8
}�q{�sdax�5�^���U����jքӊaoV��Ɓ��|�<:F}=*E��=$��2�Ԓ2U��&�߱��)�$�]�I��o�A�<u�x"}�}�Q\��BtEjz�`Q�����=�օ�<���VX���w@U&�V�љ<�
��-K�ו]��؛��c�׈�;I��~0��'�z�7����B\�eҾ����Atc����S���祈��f(����u�=�1��������j.�5�}*��p��@��7��2/�o�܇t��IVla,���>��9	�w�7���|�T[mqAEk��`�T9� �%�4�X�S��\�1=�����1�@�Ȣw�T$��b;�����ň��Q>�����z5����}�����jJua"1�)9a��<��CS)S|��6��N�՚�AK��MG�d��er���|�}�e9z�ক��7��߹/$5HND*�j�I�l�Y�
��o�/S�b�^-���⸎:oU�h8�K!�|�1j���>��)��U
;��|�nm$����̣�+��*`��3����u�*m��D>�z�;�bcm������#'��u��aoR�L�M�w�/���t�}�Ƶ�݇��2�m��y�ɝ=��H�mjߍ�t)(��{|�v.�$�s��h�R����D��,�l�X��yO
�T��~�A�U��X<M���v�/W���5@�+u�
*H�@�F��U��:���P�}�t�0e�u�������o�Bg���7nSK��!� N�*O�m���I�f� 3-����5F�a�J��)�=�����񙙷�70��F�}�k�����у�E�����X�_�OO����-Ҷ��${�<0�����s� M{{�����|�T-������"?���)=��/h�kKm�S���q���n�O�طy�,9�u���d^�Ǔǃ<�\��d��9c[I�j�J�El�i������#P0�@���DRC$@�@�v�o�U��Bt��M��Ӕ��)�*՗�MK`(�6~��$Hċ9FU���A�j�Ȗ����� ��C��6y�6]��qn�N8�Z�u�fv&jɿM��V���ci*��ذ{��ٰ���M�t�I�����KΫx.��`�F����Wcp6@6%����@8�DӢ�@���?t����xO{쀿:���-���?�ȜE�������$���������J+b�F�p�8V�34UWw�c���sD��̰���� ��~/�t�+O����M�\�v�^P��]�R(���G��a�64�(n��"��t�A���$&���̹J凗���n��sq~�p�L6��8l��K�����Rڹ��2tԽ{"���V�5�y�PG] p��%P��*�]��_�tyvb%e�l2,�4�nz�J�H�����O�Ɂ�y���BS�lt{���{�W
�#�()�=B��!����k��7�	� ��϶���a^�ߓ��:��!���`[�k�o���'�㊵LÞh�j���
_u�f�	�fF����"��!dB_��X�m��M��>�i�ݲ&l�1�^�I�X}�2�2%��U:r�����'w�om}n�z��D��;�e�M��U@@s _d����͏+)�wJv������3�i� S����,�͖)��5�{��\b��*(��Sv�@��&���%�ߕ."@�.9�4.� ����I��TS�7f�v��&��xp�7��w�!�5L���Y6�O� ^��/tH]��ur�q��0ff�"�f��n��h��.x��W/�����I�>]H�TM�Z�IZ������O��nMD�8��n��K#���(w��� ��t�z�|� ���ľ��U��/m�;P�=��_���|���2�w��b���+�i�v_L���'<V��9������]�!��x��n��T�5��l�G�z��c�_���y�w�������|�}�,��!���F�L?}l��;��=c���Q��LS��W���^2�6'�M\�F(�t3A���\Վƀ?|�S���p͈D�����lI$��_������ܞ�ʌ�ݮ�#�b2�ko��{��I�қ��E��Cc�'s��n�m��`��C���I{��[r$؆g���΍Nik*f�Pg�2�g\�Ūu�x��2Ew��֎�������wԟ��V����5���nh�U���ů����ly9i�����[[&is_�g�*Wn�)��ˑ��Y��8o�g��:��Ԫ������7	=��-������f��8�����i�g���#�ә��E��F'��^~��d� 3���D�(�WTaBf-���;t�+;�x�V?Ih�����AsL�s��ڥ�/��YF^ޛ�&E�2��`��#�ڣ�o�2� �0nԔ]�U�9���k9F5�^ǚ��6[V�
�fU#�-ON_#��thY��P�EB�S�J�����dN�J�ч���=����"���Z����R���2���a�<����'��$:����bA1F+Wu��n��h;_M?�>�u%�����/ q�U��Yr�%�r��OZwȐ�#2_��C�4�3�F�[ /��E���{�wW�����F�Kx'y*�^�;sn� ]v즶\�go�	�+z�٥k���`=����_���!��N�S��{��/&�����[oR�z�.g�t��mp,���*ն��$=aA�i�wz�p�ra}G�p+=�r�V�;��V�8s��%�Ǜ��d� aS}W��m]���d�1g�;-�s��n����rH������n�PHt���`���['�nW<p����8R3A�������������4]��[i<g���T�����w�3����[11�d�}��mϒ����=5cg�2�g��*/7��$v)���"�B8\�b�+�txl�H�\�j��^�j*�]�h��eC.�� �2�Or!���f_�\�"�h�r�?Xa�����i�]�X��\/9 ���3��,
��R�<v"���a��kJ�x�&��5�UT�
ǹ��9�cQ�dݥ2��D�K��	�h�d�;���	^��KVk��>����hIx#�a:����)�m7��{-��+m!u���c�Au�		���,Nɪ�@J�`s�y9�g[��lV:�H���qj7��#���,6i��w/�*�1oU���缑�?H����x�& uK�ɗj�+?�Qƫ���=�V`�]-´N�K`�����p�6Z������	�PD��D�Z���d#-���c��eco���hM U�𬻊G�c!"B��=�_`i����xH�X���^.i:��2����*C~D�F��MO[��3@z��I������kݬ�������Y�t�>)�
ͳ����t��U�YVȭ���ο��O�>�ok�ǟ����S}U$}���`f\��s���"���[��^�8�Œ��%���eKN��l����"8�V}��Z�14e�K6���"�i&��E�<�	�6;%X&(�/Ye�4��th�P�����µ"Y��DI�p���������=z���g=n���刴hgo�5���K���9�[�9�-s��Y��P�~��"S[��cN�kI}��	R�)gU_��,^xlw^	t�T��;��_3꛳{$��:@ċ��r�{����mz6}];�6���#���5ԈW�7���4H��D'�A�=��~��&��M�T��l�4�/�~����T**�~{Xd�!�z���MR�h�k��\���	ګK�ު��*,�/b��(��'�.�b�Uz�����l�	Z���;�=U��`[?`�]8$�u�}����Bz�9��
;����})O�C�]5���5�1u7n�+�;No���>��tb떣̿��C�V�S?��6���q�Ր�� ���}r���Mኼ'q����yЄ�.��n<�6�?~,WcI���a|t��xw�]<i�Tl�(.�	4:�@�`w�v���p��=��m�r����O|��k�1>�����ȁd±E����i��@�Z��HU�ܲw�D�swγ�0�'/�uו0���s1�ʌ�>?�[m�,���	�jeM��wT��$-�G뮪×ɏq�o�
}~���0_�]���;[Kw~��V�N����%�Ծ�O'���v�d5�����R��l7'�E7�?�z�M�wG�N�В��ho���0���5�x�e����΁]c��EHºɛ�k�	���Yp��o�I�����6��ͼr2I�#�D{e�ޖr:�j�B蜜�N�i�#{��o�:���v�q� ���y������|�`W磴�U�%�?6�.���WR���C37�����sA{\@�lmR�@´+�a�?��0oVDk��.P�\�[M=K�hY����xix��y�H�R�h��s�>x�LI�f���Q�V�;h��J,@Ih��בx2�.�9JJ�j����?��G�~��2蟲y�<%�䔅/	��am��!����S��c�U�w�n�.p�\8D4�G���k�� ?������*e&�e7���_�Hz�����b�\+V�.��=UE���(������c������X�;�L�^7�|E�X�i�6���8Qf;t2(�[�T�2%2��(��w>|:ڞ��]5xZ@�� I��X-��T�����R�Ʉr���gLg���|��BW�ܪ���cP��	m��'I^y���bP&K@�t0��:����Xh�����F��ٌX�p>9�q��c�j�j�_Kŧ�u�����Kz��f�{M���'9�b���̹b�2Z'��3�:��I)�,����cE�0�-�:	.'b�`$�ѺqiZ��	\tZ{�0�r��,��Y	�+K!ǂ��L��V�%#���(§|��eo�sV�����������3��[����5���br��c����Hi4`�ד��!Z�K�%<���E�Zc=:9���}�h�c��	�l� gv��Y�e���6��-3����'���bRg8VE:���az)�����i*���z�1�:~B�)���N�6��,�i����iOc��Ͼ��E�]�w��X �qy���R:q�� k��f�0�ܣ��Xsϔ	�n�}1�����a����K���� �.K�tզ��v�۪��3dŤiK�a��ǥ%����a�5����k� 9����0�p�[L���-	@��O���2�)��1rG��a� ҂��~��
�U�'���un9B�%I��٠^K��6���÷:�	7ϖ��:�u���o<��nV��ô6k�)V>�i%�?�m�W҈�V]��ꔘu|��B'z���s�D�en�q'D�Bn���83�_���z�,��S��=�������s��sb)�M�*�x�)�E>a;�?����NU@0}&}d��.���S|�kί��
�5=�"!rv����j�<7#��x�#�D�o����7�ky��y~����rm�����x�|:R��?��Oe~r�� �I"%�2���Nx4�ѥ6DDFz��I�\����ܜg.qK!�
��3���lМ�t
���(����p��}�qbz��W��-ۛ�C���W(^t7�a%ÒW��@uC� �jo��ѐBB��4f�ƽ�����#����v�#��w�,L�֠q�{���	8AB�&�G�kl8LT���Jp�O �x�\U?�*/bK-ʪ���cD�G�|�{2����:� ��s.^�ȏ������	��m��J��*�!�S5{\7<,���zb�;<��<�0L�� ���?u�ܼ<�G��W� ��FD�8)U[��h@����۳�_v���/� T�./�$�h �z����#�?�P.�_M��]�#M�2dq�N]��{T�5��|�?Ȥ�^V[^+a"��*B�l{���ح���{�x{ ;���=�B��T��c(-����Ӿ�~	�Im<��h�q	�
Z;�L=2�be͜X�PyS]��d��!߳o�	��B�29S��𥇩[9VZ�'ۛ�I��ԯ̬�'�#"�.�k]F�8v+>�1! =l�oW˴�;Æ�G��3Omv�]EC>P��kC�xKUǠ0��x�sNZk�*����+&>3U���E�K��6�+ˑ�����p�
a����Y/�uWk������d	wqaB���AO)1�*Ջ��}�1��Ȕ�x�66�`�� w>/�I�����y��T�"XR���^e�����gJ�p���U4}L�C���8�͝�q�]	�Ұ��ؘ(�?FX?��~hV�>8Ь�@�0��A������T]W�-0��K2�� ���pA	(�����כ�F����ן��lV@��-�\��N�:>PYI#_��[��sjo�.fj�i3�Ġ���ZHPGw?zt�d ���\S��:�:*彍��۫���i$l,J�%�a�_�)B�Qf!�o�KQ�m�~0Q ��Z��DS@������!�B6��2%���+��ª�\�T:sk`ux���l�Cm�8nW����q^�b���$@Z #9��1�Yۜ���^"�پ����1��R�&W@�j~��E�M���f��<z����ˁ��h����򍊑��sɓ����א�!�ֈ����������;d���rD�-�h�$��!�l__^3r��0��z(�ʇ��>4k[�9����E��d� <br{�������2�2�TIj�Wx���V.T�r�X]t���M��<������^odߞ�~쐃|�,=�^��A�Xn�{�+#+��S��#��q@u�#��� #��A+��� 1�O#Em�W�x���t\ĈUFL����X:FX�1��D�Jq�H�FuU2ti��%�V_H�]=z���+b.���n*ׅ���8�9��P�_��O@b&4��:�+̭4�&��c�U ��E q����N]9T�m��4�Qv��UC�j�դ�!kfY�Qx�;'18�0�)^��len4��>��&�]���s#���p(7�H]�r�1m�I��Ğ�z�3b�M9�(�Պ��A_����5"VWwـ�%s��x���ݹ�Z��-����F��"_.�#�NxpЈ�x[v�B!'�yp1Nl�>hJU��}윒R�K^�����D�s����q�c��qo��-+���T/_��m���֌Nc�B�����mBL��%c�AF� �������|��^
�U,r�����(\ m���!{ӏ������'O9X�����]�z���ݙg��{|����$�I�S��D�� �a�ནGK��'��-��3���8_yEp��3�/��q��Bg-�9KL,��>�O�T�l�+���g��l)g�$U�}��rL@�F~L%�M�{�b���=�C!jo�����Z���1�=;��I�1{%��;*�����钆"4E�\T�=s?6���t�>m3\�sG"2稛� ��~�3�<o�"�ڷH���ܸ�� ڊ�MG5���������������$
�+^�	M��k��Ȥ�3xKnߐ�@1�Ft���{.���W'��B�Vʧ].���Q��j�ԯ�8*��YAn��}m�AG�1I�����Wށ�a�^M>3%%pJ��2�;�B�ǰ4��JjS�b��eѩ��]K"F|6Tq�s���k{�xо���7��?YI�& ��/�'ܐ�2-��ۺ��[	�,{�mݛ�>�`���%��e^;��K��|��e����&33"V����~k��x}9�͵}�m�H*��lHP���ݦ��؍L;�Ħ��[���ޝ0�Z3��S�Dco	����Ġc��DG��u]��J�V��I<����jK�^uM��+(�G�E���K?2��qǸEFK��և	(pp�g�\�R��\�8�80v�]��[��HRp�~�E�������ڲ�C��q�3�GZ����)�秺�y�:C5��"'>8���EM��YM0 V%c���ʭ�����k�����DSE����j�"�va���w<�-��.�>�+���^�>�o�1�k^�����GjG��l��6� �6zQ}#�F�X��}����T�z������"_Dk�CK�v�q�6_����F�F\��s21o�d7�]xڔYP�#���1�՟1D���]Q9�U���c֌⡽8^��9��(����\/��s�����0���a9���Ps����r������U�ZA0��o�ോ�������|�	������q�v:鯸8*]�2��Q3����*=Bp;>Zb���͂NM|����MXn�6,�<�_JK6$��b�d��w'%8��Ob �?��\���}�d���8�A�=�,��T�l� �iۛ���7g�k�˭��o���"+qe�����Q���~y�SH%8��"�]�X���&'#m����B��_�+�\�G-9�0��>�$�9�3u6���k��|u93](�/���;�p<�@�eT]��]�*��?;�g�<-^��I;@�rwr@��M�(��X�[�E�F�SVT]�m�v��]/�$P���D��5J3]{9�5롋�ѾV3��*�J��{=�~�i�B���u�7r vt��_��n�H��O9V��̩�f�݆�Sۣ��ec[�A�!?W��LꋖӄP�z�Auz0/{�9JC�8"b�9�6>ի�3���w\bG��m\K�	�}P��?�t�f�;O�N�F����� x�v�ڥ5�`�Rz����+@K]gJ:����4��&��I�_ A.s�{6&�!&��-�Ȕ��d��i��#͛.�-���&�f�� ��_}a�3h����wE�,�3j�d;)S��|�&W:c�T5���1�̳Z{�š�ʛ��/�"���e��E־K�(��F���J7Jl �ʈKf�t	^��o�B������ �yt/�Z�C���R�Γ�h��نF�ˋ�6�`g>:w��i��o,*���N�*�*`ǰ�Q��` '_���������{���	#CN5�>=�N�ex�\�7j�}�AD�:}ѷ�+�2�%We�7Bqى�RW�]W*M�(φ\��oC��������=wƉc�X+�fbZ�z�b����ȓK���ס�N�Ԁ�uM�˘e�G���l̷?�U�mL�����y�Z�L���-�؏�BV%3�*�ѹ�a����u�0q�0ޟ�<�a���˄�/���@�#2/�8�X�^�p�0)�t���y�yq�`��9dF�R��3�ڟ���	��=�ʀ�AK���6�@�E�9����Aӱ/����l(��ᢙ�d�:�\`>	o�A�U�V$Ҕo���tj����g2���qT�h��:�z'��l�fFd -&�y
R\�8e�?�9
J�]�4����o��W��#r�>L�S������5��0D皼�S�	s�Bk	��Bw6�v`��B��c����s��%����}}��lzp)���b$a��5d�v����Rz��Dv���O�?�3u��Frf6�kFx�l0-�*�'���$���znӇ %�^�ɺ�[(C�o�����i�h��c�{��iזu>���?:�6�z�"g:�p.\���=F������ȉ��"������ƭ��}��;�<��"�)7@(բ�$����@*V��m74ᓅ{=���I��@�����3QC�*)�مU��G�_c%�����1~.�yJ���U�?�͑���wE��-��8-����yR�j.���.������5�UR{�SbG���l��fޜ��ߣo+~n]ٶ���l��qYP��w�;���o�W�x=r��*�%��J@�C�?�𧅶�caj���!֒#����i��-\e~q��Δ���MV-QP��;ϻ_4�Y�-V����A3Ci��Xi�0�E_���|����Y�U�
��@7$�AD��j;�lO$��=�%�?�M.��ɑX
RD����^z�32��J�77?2�8ެ��R�.��PC����֤(q)옘<_f���r����].l���Tg	��x��I)T�K�y�M& ��Q����VBi�x॒ޘ�N�k�/�Q釿�N�C����75������X��](�;���<�Vn�v�?�;�ٝzWәs��������'"Ld�;�Y,�l���ˉd��\�`% U�Br���;�4��`O��#��Yg5H��Zu�"2S�7v`�E��΂�A10`Mj����"uG2����j��{��%v[��j;�g }���?;H�=��0��j7�J��������?\~ɢ(5����r�ٓ��4��<�
V��Rɾ�=����NZ��.2��lh���]N�!�����C:H���$i21s��}4Z}|G�_ܲ�]����?Mg�i�N.��נ{n5@��A����ILu�!�+;8����3ˎ���#�'���A�N�.W�Ճgly��2Ơ;�u��|v�H G��ʥ���,X�1\���2��}��	�$Sx�v�͹ef�8}eզ$p�r- �嶷�����s9�^/�9�N*�����A���x
?�~�f�x�V`n3y����+���ǣ�ڮ/_���F����^�������k�ǩ���;U'�(�{{�D}����n��C���M,�:/J�V!�@�h�i��9OY?��;�����O��'��2�8i����'��+�����L���mU���+q�'Og�8��%v���Qe�8�pK�ᬛ=�m4�����|N	m���ԋB�Fb����*��f�X,������x���8ƙ��u��U�W���f'�JG�:�G�*���F��2u�F���a���芔̬��}\�MnƲ�
�Ik��ݶx��Q�[��d^�|b��;����I;z-���2�ti��sѱ��p����0��6���l��)�A��>:��ѳj�n�fC��6�~vzi��KH<��[of��R�j3j�h��Q�Xčn���L8�ǔ�BaX[��;ϐY
�]�s�BgF��r�<Lnf�p!3�<Q�z2�mJ%{?QJ�Q�k	U+�vs�C����Ǵg��%z��:����M߲�2#�`A�L����$횑/���ma�@?��ɑ����!ɪ�r+9�0jKOUEl��Ą�^|�5�؄
p�;��|�����)V�Pe����[����x���d��O��x��b��N�R���ﲈ���P'G�a���f����	5��V�����+^q�*���tu�� �ϻ/}�ۺ�D�����nNk��1�jp	��Ț$_��i��y�n���zl�D��_1�r�ܲYT��%�e(9K��^ed����x ?w��ӽ�t�^���	�u/6�C�DCܻ6��Xz�q��ڼ����,�đqs�=|$��҈�[��W���W�k�|��t8�+� �)q�E��g\iu3��e�����!���F����7�7?�O��DU�jW ��J?�M��>�
"zHlt'�Can�
_@�4�IA!W#�9�\to�,r�+N���m�����P���'����6U�(C�10��q����%$v�Z�k����?pIv�|�g肃�`�3�q`;�c9e QQ�9n��׍]�89�o�F&ȩ^7��a��,�Dј٠�jP������*s��k�-\:�F��Vz+] [�-k��!�9]��5�||g�=�������ug/��=��`���Dr���m�׳��r�L3A��Y�� NW���T��MP�����Y��K������@�c�j��h�����ч��ϱ�qhel�ոV�J����;�
�,2g���z?���R�m�����d���| �tj�Afr 4iz1й�b|�9��H9
Ci�9X�'�[��"Hrʁ�D)��[���'ֿ�{��EN�s�#�nmy���͐U��G�>����� X�s�)�����>�@�jYf�c��؃B׭��*5�LP{�j� s�	j-��j�Yf/�� J�Y����>�^����V�Qбi��_��C����[��8	 �V��0)��W4gG�|����v�Y5����.�K���4����075�x�yn����M=�{��G�
*�HIa�/Z-"� ���VОY�Ym�LS� ������Qc1:����b_�����N��i�	(�<��J`�Xs���l��+��lk͏;�,�T�u���T �W~�S)Ӵ n{�����y��W���m���A�nṕ&��
�����ʀ����Q��*
W%���5�TRD������(HHw1�PC)"��9��s��{?�?�E�<g��Z{?�9�Q���m�i�3-�/����p!����ᾲ�!��Mԫ��;fq��N�?�1�˙%/���z0�;���д]2}��ήH���8�۳�^[�xWAK����ٟ�:�d��'gC�IX�Oq]��@���P/���~��Cw��<��j@r?}���qI�U0JG�z7*�u�8��a��Q<�I�\�r�3��"��TIG���%`�^Z������f��G��'r�;����~�u�+�O�v��g<"no�P�QC�����P�KLDx��F�W��Z�-w��ɻc�����d8�����v-":���aj4��Z.���?�U:H{]�S���&޶(�����3.�\a3��>���N��$.��a/z6�t5�z�EN�XU��&aY3�tC/}�_�9�+����)F�uW��sU���𹃓�ZanE��	�Z]��y�0���� �=<"%�Zk�����Q���Q=.�h����,��Ŀ��?�:��g?��� 
�-���Z7�H[�C��>���<�2�D���d�
�#/�ӸS��u�W��ˤ�T�q�G��$Ao�z6G\md#B#�6�l&S�T�-Z��A��`V�WD��+�3���[�.�y�X�#�Hl�"��v����"�8�q�"z��jk?��~�.�f�f~P��-�*y8BY����m�E��(?�L�	%��y��%��d���s��]:���CkS �v��c!�����rn����gF��2E�J��5s�g2�!Wk��A8���뗿�'�^���=�8	\��.�|���F�S��u�֍\�����,�UfE���&�a����Y�X)�v����_$h��w�r��� �-�u��{��Е��ɱ!��~Gn]2)�pټ�]b�Йi���q>��Q���UN�	Ug�ɱ�3���nP����}�(r[��9����¶tBx�������H�P�� |�#��h�<9+P�l����(]���M��6<�&���r�R�8+��cĽ���<��q_�"B�@��KMOO�5�+����KX���ݜ����,xG����"xZ?�_�v�����P�1�L��'t�n���G
aM��(O���q��\�����z�6#��������f~�-q����'R�G�w���3�`��0!I��� �����5���~�)��y��ێ	�Z^#�E˸��%�_��k�x�B�̗��C>T�~�rogk6��������ݭ��ǅ��Z�yp��G"[�i��0)�(%�4��ZB�]I�;jz&]�5	���m*�l$���ź��{����і��0�����i��H��?����@Ka;���Z�$��<p�V�<�������>q2 �J��`2�.���N-d��ҥ�t���������.~��uQ6��G�Q~ 7O|���7ż�h�:0$_��]1�t�`��w��_	����Ec����g�3��[*Ą�fb�Ib��O���(�z�qe�B7��1���1���!��D 3�a�������/�Ϸ�O��a��r�N�/waYt2}�¬��(v�	� o�Ϳ�r�Hl~��dQ\\ njA�����2l�0z4�р�y��_P��c����(���,��Wի�c��kss`�2�����K�$y�!^�����|":E�n�>�b��g�>=1:x#ۥ �ـ���x�<IIY�Ŷ��-8�PԻ�ט��.
9��RN }�)ͩ&1��F���uօ��n�����1u�b��q迌~�����h=�u�i=��,���OȢ'�Ѳ�>+��=��Y�x�ey��I�7;Vz�l��t%=����Q���|L-F�%�:~�H,�[��%�K㤃��?=̀O����\�]'}�5�����nzL\m�Q���=�0��Q��-5w1X�b5Y��ʶgpi?C���
z?��I}�g��_�;{� ���w����Sa>�B K�s�oPW�=͊~��CL{g�m��~AC=�}/�f�����np���i�5-4}|Q��pG�g�d�jZs^��ۤS=?��أ�+�mԨ��):L9�~�>:W��_��	$�}�WP܍|`zu��s�%.Vc�Lt~���lH�K���[a��Za������l#�qOJ׏��cdl��6p�
��l6����V=���dE`kq�W�v+���F��ɗ)/��-��W:�ˢ>Ua]}�=��߈����. ����D�G�Z��P�Ѯ���dMv���[=M���3����@��g%���~��Z���{ַq)(Z��
h�#����|��R=�k�J��(���*��d&fR��}������a{�8�5���R�x}�%��˸)��=�×PT�<��?�F7�C���S^B�*ب31%��"�i����Ti��J�c�nw�:�1c�� ����~�	bt�7�M��,���z,�7셁��3c
 )���3�|�������֕S��XG���2���8�:�L' �Vވq���#��8c��ɋ^ױ*Y h#�@�K����c4/\L/`��~~�@*d]'h�V�������@��b�ź��iS�^�N��z��6�̄��I�K�l;�_湀*3[Wvc�b�:%��*Mu����gg�C�T��s�|ڨ�uN��1ʣkG.!�'����}b䌇�\�f��I��sZ�ɧ��U�{$�a�͕�R'����_��nڹ2��~���ie�;�7<� ��!�0��Ԏ�*S��-��!��8n@�>��R�	��gip�+�4���N� �o�3��c�=���{8y�h*���*������e߿�d� ��K@��KF�r2��qE�(���f��J�P��&������#t\Z�}��Q��[�jx	+�AYu}�m
��;�Jd4�S��Y�:�8���>|� 4L:�4�y&V��y7K�A�F���Y��_�q٫����-uI��uLr��=FJC��7�����P�u(��7A��j���Z����м��!V�m^Ȁ� �F�ٳݎ4���~V��Eb3��x+}ǎ�A�=��_�/L�(kӻhxX�p�'��F�1��3<'c*��7�|�1��*�+��;�l�˿�}Ҹ��H�7�Uă���h?�i��gû)ᕅ�\���Yz�ߛ��t�� 7��qp<��VK�]tk�G���A�x�K_nR[,;�y�a��!�� ;��uȭ�S�!��]��ǁN�ue ���9 �ЏM�_�w����~Z�U�F��E�R¼�$�|4]�l�)��hV��cѪ|��O�j��x���Wl��;�o� 3�M��~�:�}���^�����0չ��vs����=�̈́��0f}�*�<q5�[1�-�YFUd@٬���ˆlʌ�Μ���U�^��.ܼ�� ���yȳ����	�y���'�1�}\���V?9�p6wqi}����aw�+_1�j�J֧�n��UU!�����<�ɧ�v����FW@Lf�G<��Ak{9�!�^�� Z&����g�P����<�zk�(o�ӿ��3K���
�����Y�^��Ex�������
��q)Cݞ%_l��X h=,��	�h��5���7 s��!q�l��v�x 5+T\e��c)���J<*��E6���z��\he~�V�X�H7�$y(�����Ou}1�΅x(�*���ڜ�Ax9и�4�����5���O�
q�8�"%�m2�~��'�om�M�ߍv�_}ոg%��o�3U�m}?�Z Z�X��

o�w!��� ���Ei�@A@`�������_9����ˎ�&z��5��)W���G�8G
�r���_��᥁<�:�um�� 5������Φ�y	��)RB�~�����f���ӟ�\xs&^�����1�A߉^����"�N/K웰��2���Ԋ�O�5���y�tqyM�5�S[9�=�N��٭�tm���h���2NK�~�����8��ׯ��.9N�i�#ݥ5+VK�7:�ê�`p}iw:��i����8���B�K=�5����
��}�I`%�C�
��.+洈[u�zJufi 9����j���R�槰Ӷ�|����Kz6�e�"5��X�)��X�zm�1�F7��|V�A�R�NZ��g@�Hf@5`�l�3_E����3S�O�hٱ��}�[���=�4?�UU� �Nf<�mVU��|��������т��J��ZW����Hmb�A��y���)Ν8a<�4�5�Z�iH[ɦ7 @�K��	�����q��!&���w�r^]p�|8����������'��p v�c|������W��6x�_���_M�Y�TN��g��k��RX���$�{v;Тa�u�{pH�G\���U�m��a�ݴҤO�y�׾��s'�䔥B45�Ϛ���<I �J�� U�
��0��x}읏kzdh|`drfƷʶf����½� 3�Xx�
8l�>zY����t�����@��z�3N�A����Y�{nFt��@bFU` SR?�1d���;��Z�!8��p�?̐���5��,��j��7��k=�d�/~��� n�RA�����*�������>`r0�lTQN4��xb��p�� ��z��k/OJ�Q:�Q=>=�v���i8@�K�E7��ی�..a�R�)e[R��B(�1�����)�����bk�\��_����*�+��61t���1�e�%� ��x+C��`t�������y2Ӹ{�R{�'����.1�扰�����I��~$3���2��]��K��s�Bzo4���ח��w�P��|Hb����6v�Hd���#��0���f��|x��'ʫKirc��۷N��e5s ��m7�aI<�'���$�9I�9�ҺW糺�`O�քJ.��~�x6�w���g�����8_Z,��ޢ ��y@�!���v��(.��7�|0ٳ�����t3*@n(�Eg�)ݱ�j{�׷�Ք�śI�e ��h.[��?��A^{|Z2�c-��I#��[Req��t���EP�<����d�>�jF�
�^iz8�,�,Z���NΉ3��ss�D̥�ENW�W�ͽ�~x�!��ؘM���a��䓎uCQ���ğ�H�|�h�K9��ٵ*͖���� �*��ݘ��*��=9�mѯ��[YMD1�a��?����D�7u���ݞ�g	:��)ҳ�d]�˼������\�a(�ߐ���Eb��$:y���ɟ3��dӃ6� �@��?"B�iXu0!��Y��$��l��Ѐ.T�.z�ELK���E����B߶�8��4!�̄��ՐCn�Oݗ�	'�9���r9�wȽ�=��|ݎ�}������
���i����[����j�cyx��-�m��e�I�j������a�
/Wg4j���8��8K!2g`�.-D5-���ժ4�T��5�[�&)��@�>ݎ�ji��m�/t���5G:H=�����pog�7��϶p�&4�H��V_X����s�>�~���I$!��l�YS� 2u�`�����v5~�?}0:��j��d��]�W�u51�w�����쌄�"�b�y<�H�Rey�_�1Q��q�dɓ)�#�3yfx�6#"��r5+t��̱��f.|�o��7�a�O�GRނ���V7|��Y?�u�$����]�g6E)gD�k�̿�u��9Ȣ���ޥ�+^W�f��I6$d�XN�e�B�,��g_P�Ud�{�����w��g��x��j��t(,�Yh����o_���k��mg��.ГB����E���}zF��`��<p��-���I��2iG�����L8��Y�¨ƽ\Y���4���c��qn���p���F���u�_qG�厀Yz����L��8h��MV8JD��1��.���=����Y����>_�����p�Z��wN�'��^�tΧ]�BcH��52-�%	̰z���f�Ftʕ m�ĳGj&�1J��R��g�;-	��p~h臟�?}j� G;��E���=bae>x�\^'PX�@�c����l�ŷZ�gǇ�<��hZ��e�)E�V�<�ϑٯ/�J�|�P��*�����'��ߧ!z�ٳ���R���:��)�o[<��~}�VT���ı�0�0���OIO���'�R����6��V��E����9<Ulx<W�����~T�f�fP��{��X�����%`{Y��\m�X�0��MNw��`A�@#`�f^݊xм=�4�hXʆ�ݔ�S�Ef�������&��ieIK�%�u���K�{��������Op٬�t��:�RaJ��hN�����Y�A˳���~&s�UE��DGOm��E��71���A��R!�r�g?�<OU�*fg�Kʫ��^�1���5�v�V��Bx����l����c��^�P�?���`��o��:M_�0r�l9�*B�Qz���ķ�(P���8����j%�~V%�|��6���zh3��b�ga�I�;�rt.Y�Tw{��q�|C���(�$��Y� _X�A��;|��M��v�u}Tߜ�q!#!�Yd=%�l?���kT.�e�x�I˨�"2���=�]�B�S�N�K7j{~��R�Js��{��������:S��e��iDK�#c)�͞����*7����Q�6�#1�HINFx:,$�9�.���	�j`�gM΀S�YF���u�oxQ~1���[QqA꾜'��=�O��͍k�On k%JNu<���*WK��M��c���.��(�cM������0���^Q-GR�Rv핃}l� �J}�^d�U4�M��A�P�R}�P(�dF�e��.��C�Т�äXV�����Y�L-��Mx�s'��'!Q�t�]E�<{{��GxN�^��BN6Q4�\g��,���1��gg�lrP��=>�,	�<xP�RWǐ�Sq�%yg~������x�y�,*��iD��b8��<�,�(���H�nL�)���蹞��K�̅�BĽ����k&�/��8`Rh��N��gN��ͻR�u�\K=��:R�x��̼<�P��#�^&����>$ �HG`p���/}Y��r���#H]�$ [w!�Y�%#�������0�
 �);����C��1�#�ao�
�~��.2%���n]�\�2h>�Ax{��n��4TU����fL����=;��o[�^b)�VE�	a��������whʹb+��f3�	M�f��$LBu�,yRBL"@�I<7���/Y�/�=en#i�'竉�~D��877�]�M+͖��;�!H��q�:���[{_�U�!��q��!��iE86���?�ʮड़.ʔ��1������!6|��$;<gNV��x[D]�@�fy�I;�����W(�$}ヨ��ȿ5`��+J�r�����qJ��>����\���7��B���L%18�f�%�������l��ɭ ��e:�.�?k;�^_�a�d0�]�5Y>���i_�B�j��IGl�t���v���p�-��Kv�(�j�_ɷ�·!�|Z�/�+�^�HX�L�W+��c�&��Ck�LV�:�Ph�u���@���ډ��T��F�D	8��
���˳J�����>��o{FnǬ�ȩ��*�y���uʓ�*���������~
X��p_�Jڻ�nc3��df��[K�ҰV���G�*�2^��S���cu��b��4�q�����@&U�AwK9��S�<��l�v�7^k�>լ&�j���e��.y}���K�)̎�����z�K����B:t?R"W����T�S�Y��aqB6p�f�u� �E��ܓ`��%�d����������S�i5� %5K��t��{b��꾂�s
z�1�cG9�G�H���u�P:�ILd�^/��+}�&�w�⑴�����76Ny���_�G�D"
���{cA�����)JHe�ښE��E�Nn��4k�7v|(r�~i:
A����͝¸a�E>�U�z�O�)]��f���d�(3C��F�OAu�Hʀl�ա��1�0����!�ooh������VO��rs���d�ʢ���:(��&�'J/�gr�c������Q�*-����H���|<}%$���>��PQC1i�<����*k����[�{	����g�d��1�C��\�*����M���S6�P��b\^���9�>�~�c�̫�G�Ê}�1��W�2��OB���:D��S�=�zt"�$�{w����.7~�H#��O��x�_��kУ�S��ګ��ԓ�&���L� #88 �|��:߿����'�#tdƤ��tb##7���^�9F�ȩ�h��'?A�Á�Y�3� �� m��ϒC�`h��^J�+a,7.7�[�6=���
_�r�1�1��6�a��li>���~kb��͛j�TV�ʹ�i�nl������̥�H�(\�k `�1���/�2ۊ��?�ؕ��=ü�Y�*]I����X�V��<<��o:�=R��ɥ �w��qm:�ž7CD�Go���yS�`]"�Uޚ�}^����5F�R��y�-��}9�`�����M��#;p��\9\��zz\�6���p5/1Lȉ��gNDjB�C�G5E^95�䔁����q��TW��dC�32Gnf0Hʎ�?,"��.��c��44�%���SG��g�'��_;V��*�g�$�>��>��������(U?e"�T�'
M�ì�@�B7�u-�;dVR��?��&�m���>̴�=�yɒc�V�幋phy<�>�����g�+��Q~�K�f�2�l!Ʋ����bl�ni�Rv����>A�:EVh���n��h�[�܍*;�C��h����Ͼ/r����TP�{T^@���I��:`]\��?�P�
eT�G�U�~�����L��~�.��! �TК���w_�S�ʴ�J6%+{��=�Lc���"g��=	��; 2N�O6}�N9Y�I�e?�����AhFG0��9�]dd�ڜ�z��n	�*r�}Cc)����R#��_������KӸ>��4泆����*���PA$Yި��c�@l�YQ9{J����k� z��US�X]*���b�G���cS&�JΟE�Q7�����(��MB��!&TPM$�>U�ďT��R@Q1"��������'Y%Ś�46�0�-�=����� ���ݓ�g#o=���9X7���Nj۸�O�'�(�'����ě���9\�����o�x���j��b���������5��P`� ���Xz����y�k�&ʵ��)'�Ŭa��ù(ޔD��KN�nT�K햋7�U6FY������s��`D�l,��%1`�R'N����|a3��Z�.�v3WkBg�n�V���%2���]AW���]z���Z.���J�����T�zO��H�����m*��%Ge���@�c��<�,�b��P�a���}��q~� �7���-��MdvJ�/b/e��H ��M�?(Φ������Q����Y]�`��k��p���K{>��;��<+��n�E�pu����>"�$�~�r��p/��I�Y}n�R�B�s��j
W;u�z��X��|�/�����O[2��;U�H�p�����a�V͠ AV�S��}��ۓq㮺jI����+PT�:z&�RC`��qL>a����e�Dx�a/W>2~�_��	��ڳʯy��>c��V�O��H��;ߊ��� $C�bo6� $́�j]�Ǭo�[�Sep��|w����MC�LM�EYػJ'���2u�P�c��⧟I��YY�,ڙ�R�B����u��6U!�����w ���E�|�q�59�!95����L�jj���a�	��w�a�Q��D�W����،��H)9��5	�9[��c1���ъ�.��g -��D0Zs��3�Y�����#JŁN����gWD	A�m^�Ī
�o�Gl�w�=}g��b�ղ�ћ��>ɓTd�U�8�?z�c=�&;"v��������|��O  ��Ж��MFe���}��Ϲ5�T��xiR�cI�:b���cb��J�ԸT���'<����9TP�x��q)���D���o� E��(���*�v�/uw��0���t��p��P����Os�2� �k�
 �U�٪��'GR�(�X�:V��3��ʆ�/��i]��ɏEY�hx6���3���Җ��F٣S����ɏ�B����o��˧̤a����z8�8�;�|����� կ�C��cDB)��yr])� QXu�԰E��?j�$:$�6Vݧ�w�ж��������'��@��4��5h0��
<\s�,�"�=�<�%��{@r4���5�N������H�.�ǐIJ ���.�lһ%?�͵��|��f]��Ĩ�K��8[@�Kq�Yl�%�ɂ!8϶���g�:pF�
��
о�Zw���3�N&ԕ�Mt"�a�r�#�0�P+�ME@�}��Ia=�˚���4ݟ�~�u�A��YG�'=I���@%�+Q�h����,�O�&�B�,ε��#����t���)��������~|h�^J�4���.Bx�MR��!���i�o�<�%;�K���q��d��>�T���,�
�jX4���}|+����5OhAb�񈷥.�@���4�G�B�u�-�
[�ξ���e��c%Ph�����)�T����S��홺Ӕ�/������4���c[��}'���Z�f%�l���\����彵���C9�Ȓ��`�x�c����kc��x�v�/�,��k7Yq=yņ��}S�1��t��C��f��^�o��J+��=��}�g~���T+���?�C�S�a��t��r���&^ۇ��Q�4�u�_�w��f�>ʯ��	V��f3|rJ���d���3�R����a�{�e���9{�E�����ܑo[�@�,�="��걺[D��]�Kk�]�Yt���S��糇v?m��{k�[�A�%f����t����рZfa�iyZ{tX��x�(=y_7�^����y��r�� �V�d�Z�.GIAQ�6C�(勯U���^�g���h\�Ҝ��Pg_�l��4F��mɵ�b��%�����i��jy�aQF����AC� x�I�	�A��U�^>�+�W���P�G&64ꂠ��&���]�����&J��j' �Φ�lreg�!�Ks�Md�Z='�CPK �E�N<��:�٦�`���]�nfc�&ﺥ���|�{Ub�4Q�@���j�%/���v�~bk�A���/��]:�S ��e��4}�B�4,�xJ��û}a��k�����;��j�q���K�5�^�Gw7�ݻ�58��g�w�h4�n�(���-���<K�C;�ˋ.u%5��:E�[���Q��S��1��8썵(�V��7��rg��{uKC�����+f3w��Re�k@_�����oj���)vtZP���w�+@n~��E�5Au�E����]�s2:��|� �e����T�>`Є��t!��L��4o��WT Qrm�h�^V���<�6)�M!����j{ud�u0Kf��bW%���\r��� �@�=�|��M������YC;����G?:���VN����
�r��>}6���XNPY �4���˓����(J]THs�zN��{#�_��w���Um#d�X+��-� �:�v�$Iw��\a�0m��!�]���
���%_y����C	��a`kSF�m�/l�8:��!��9����2�I�������]"�?��"�)����"i�j�M����l���]7S�>�� �r��� �*�] ��_���coaܯ܊eiʟ�,1��Yn�c��3�����gL���R�%���,�z��r��0&� .��<Q�~��@k������y �Z�"o�n�C�yqHŏ���uT%@�n�T��v�G�'?�Ss������N�x�D ��� 7�*�Vg�X��jILt��z���׫F"��aJ�S �T*��yz9�WkC�Y���l�{!K��w6��nv�1��U�R��Z�]Uu�]�^X�I��[)��ݾh~�&�!��#@�so���ԕY��g�Ϻ�5R5�1��]E�l�������H��uH�t�5�=��R�rs^���p�h����T���61����i·K�B������n�Q��,�qҗL�dᰔ718��ۛ��n~�K�o�.`��>�QP�j���J	�6H���m��Gk��߆9ǰ����+i}x��i5+W�"gΧ�TL�	�
�gR5��/�K���/�"�5�(Q��'�������R1p���/�rL$3l[*2jv��$rF)5n����|~��|ﵶ4hx������޻���h�L�P��M+� J�����)1T&���5h�8���a�z�QQ��(rp��Ɵ���I�)Of��F�����ĿIU4g��.������<x�l�x>�s�����/Û�f%eo��}f�'/�E��V@������T9�K~2n��<�th�����H}����ܙ/y�b9e��c�H���s�����0Zꡚ�;N�|��^�L�mh�~�\�'`䢋/l{�ʻ�d�>��N�sPpK4*�3ˎ#��j����G���rɢ�lI�[�����N�đ4d�� :�ڢl��u&��r����� �
�X=�4�Wݜ*ѧ}Bhԭ�� �E��W��0��饡�r7i�k-_G����<����n}Z>��B�0��e�o���p��8��p�'3�J��I���V����+N?�;≭K��p�$�h/7�cs�dvp�N�U���Hb(+I�̙� KC��9����h�R���{8��3G�Ym|�.��,��H�Iz��Y��-�V˭!����꾃���k���#Hp0���P}iJu2����j���/��M���u~_ݖ�\�GLt���?�\ǕL��G(����>/?i�#�5#GRG	�.�Tw�<�螿���R�&]X���r|^T_��&{���hS���3@���f���c��O��R�崤I�)��;���F�'�|�SSB���
^p�Q�p��h���S_��D��;��!�;��s�2!�zߡ��l�;�t����ى���T�V6�p��#|�:Yo����m�>)_kB���k�\X�=!����*��,��ߡ^���	t�֢���kRuu�d 9�������R��w<��o�[j�F�c�����1�P�U릫��`n�<�t"ST��1��`Q���6�L~�R~y*�%����P���&���5�X:�Z�Vqkw��"�S�*�P�{K�!#0�����	���A8����;U泆k��s��)����%`���������oũ������q��ђ�s{rK�F7M�0I�n��vn�4�^���?�ׁl@tFe��+�Ŋ��T��*��>�%�+��n_mn��p��L��ס^u���g�~�-7^Lp�VD|��fM��£��2Ax]�n�e3≜ܲ^��������Rۡ�zzc��v	�;8�w$�&�zɹ�#}<m+H�l%�q����Q�I�����$I�8:pl���>b���ikq@y?�t�Ω�h�i��-�`Һn�d'
#tݩ��fc���HrM�=�1b�l�J��O׻49+�7ŭ��9_�q�&�C�o��+�*YK03�Np�bG.���&\��t+�y��7ۋ�"���PPP�p�����P�._�fc���tݲ�Z0�NK +�բ�����h�(�ԛ�Y�d)VF�hMY���1B�	N&#%mM���(%z^� �`��R+��x���ᄎ����Z��v2�C4�>qs��?�!�~#��ϳm�R�ڰ��/�Wl��V�����9L.p�=(!3�(1d5��6,�>��%�������L9.�o��Fp��s��RdG�$���R�A�d� ۠io����x�\�e�����$��`�ɑ�Z��q��vX$��/ܽ^S���HZ�r�M7{|�>�?$���g��z{��U�a����Ma�5J�yM#/{T�|X5vX�8s�l9׾��F����3���!������|�5��pz��2��˻���G��L���!@� �E���d]�j
F�i\˽Tx�@z?y"#�P'�V�Dr�A�"����ZZK��	��P�Oh�̡�6����s��{�r3��]�㧷��uG�Y��WK�\�C�p��6��)Gb���`w_��)��~`S�D�z�m�l��,�}.�Z?Xqpi�%>2L��6_� ��+KV,#K������o���7�˯Ҫ���n{!����H�ҜU}Bܐ���G�q��],>��F��e������n@��/'��Եg�~4�
������䊥�`�V�u7��
���QF|	?�Ûl���h�����/v�1���ox�6N�<Q��P�s#j�l�|�ܰ)˘�O"Vs�We�f ���Sf�շ�h�r�a�Ks@�3���2�X/#�ܞs==4j��y�4)qimq����	t�w���������p���n7�}��4����=�ᒊ�5	��4�RXZ���h�ެSh6��fʅ�C���;��[t~�Ī.�}���[�AB�JƓ�vG���=�P��F"avq�b��;�u���\"�Y��d���$�l�}sXK:��>Z �bT_b�:窇�F��p��H�?]�_ۋ�}�����G͞nJVX]�Q�/�Zfe�|Z��������+%�M��w�݅�}� B�C�Ն�}	�4=S��r]��C����$��������q��J{�Yb�������Tl�q��\�$V��u����\}5�+�K���uh��+��(U��B�R��Wj-��(�ä@�\FL. 8�vY~��������^����aA8kWH=���� ��t�y����W]?�0.�4]���1�U��Y��
1q���5�g� ����%�Ҹ��8�q�:�����*��^(,_-����p^b�P�e�/C��t���b&��V�kڢ��?��!��L777�iJiq�\���	DV����w�W3��� ﰑa��O,{�I���I�*@O0�~���I��#�7>����Tͨ�h��d��vi�����+���N�֍�%� _��ˠ�Q }S;D^��^)=y��!�%MY�[��Q�Y�)��=�cE�g-��+H\�{.�v�_��˓PZpZ���z����]{�1�����LI�-���]#�fYJ�t�����{[����VM�!@��|�mu�uf>�:Fɏ���ZoZ��+O<�B���E3w	>�1�v�	[	�����K�1����pz��wmyT�F�m�{;B�өׂ'�d-?������i��C�w�i��V�	��N�T�;�$H
J$��cP��3%ˬo�f�\�?]MqyA
���s��-�#��hC0�|KWy����(��#-�Y�� w���)��Q��P�����,��QP���	���YT�,�`���p��;=��?�J�EQu1�
2�E2��Z�2�ֹjR�W]Wm���A3�QZ!�\q/�a�>�HE�2uuX6g�Q���ִ�4r�]PՏ�G�p�qH��4��{?K�� ��T��TQ ����#\z4ׅp�<�Ѡ�����̠$�wV��cy�f�g[����"*I���(�(�>�aj|�gؠ*C���P�,u��_!�^��T�U�͟��?�+&&Z�䚳^9O~����<���`��5y�B_ -<���૨�E^�v�7-%����p��5�,��x�,m�?��	��;��G_b�����ʳ6����4���۽9�%��iCq�,Ν�x�G���$4�Uڸ]D]0ݢ�%z�e#FQR�-��nm��>5Q�rjq"�(�d�P3��ld^~�d#�1�:�9R�c�<.;vjjF��6�{�R�I��aɔE[��8'VBn�
��k�����a�U�#ul�����u��,߰e�M,�����UvO��"×tCk� ���¬��"�;��!K"���:�	c���W�Ĵ�-�:%�HW۽G�0)�����,'�-Rqx	h~
0���I%����k�{8�y]��e��r孲B��K����>/HYZ��DS
C �&�)z�N��l�Zih#�ޏ�U$� ^cmj���TN�'��w T�.y���d괹k<���SSĔ>��L�I�La�I%am4��ު��6�PA�f��K�u�>���pEG���Ϡ�{��H��KI ]�w��;Ǔ��~!���.�lo�3\O�Ͽ3�x*0�������K'�fH��D��	Y�r�S�f��� X�D��:n2W~����=�uBڮz�8x "�V�%G����+K�@�e�x���ͫI��7-H��'�]P0�,���@EkY����7�?��,��0�Qr�����2@7m���n�B����zVm�T)��dQ�M').�k\���;\'��n�[e�fa����,2<A�,uӦY��X!n(o�Pxw߽o#1�����A"P��u�InL\���.�6����ʜ���o?\؅E�
[K�a�'3�������v�289���Y#�����'fI�(C�<����T�#���rԜ"�8 k�����%n���{ޣ��{`�ϱ�]	n��˨c�:ol�2*g���y��}֨=h{֌�"�6w&���2��w>��H���$�k�����c?#��>�����}p���j���找v��-��)�y��-B�QZ��{�X�V�&_��� Y�Y�C��?âx(]mXFr���/{�.R��B)aH�b��rV]�����kT��3��D���[��MU�b��ŉ6�ʱ�|���٧6��׵�����lU��j�a��<<9H޹��ړ��[]��k�K/?�g�W?� �9��<��Rv��u�+k�o�Lx.�X>6��w�5�g9��a%�U2�4�s1�},dZ��:M����&J�E��zlӮbI����7�G�ֳ���7۶�@'ݯ��Ul�?;�ݓ�hl4�"�h~ʝ�4j�q�(Z�q��yXPN���&�!p�}�U���X��ٜ���[�)�/�ӿ���[�ve��������v~^r��C0"I�K�t>�9�����U���i�l�HJ�M�P�����I���dC��zT��@�8@:̭J}���X�c�"չ���o_:7�0"��h�qѶ�:�1f^w�R�i����(!�1:s�5�j��h�)�g��x�c�e��I���Ŏ����h�#Kp�G[ 4��c͡4v!�.:��
����ќ�r�aOs��R1����X�k����\F���v�W��Qr���Ob˷SN��Ngʈf��^��������C߶0a^u1 �6@�;�Y���βJ1�6���5�u���jKCc�	��2�M� ��|���X���(n�s0���0�gi��qE�������t~{z�X�N���U�{�k C�H���4o��Uu�mq�NP��f)p�OdXs�@����E��Η6�F��CK)��*Fџ������=���/ZB��DO��A����}"�{e�	���0D�����=��;3����߻�͚���֜����g?�{�3�[��8@�Ѹ��N�����\;󈈂,��n�}ZA�L}G����:� �~�/`���Wө6�h4�z��Y�K�p!��7�SE�����P����B�٦c0��R�]����D<����j�9O�J��a�蝥8>�iG�t���k��"Ü���ln����AC��M��kdG��L��+��������M'�i�Ñ܊*�OR��i�64���	�.�;q1|͖SV��gM
�ufKi�E)�����\�|ٗ��C��!���My�o��)-_%���w2��N�)r�Q����n�!�I�5v)��O��ۓ%���|췮�ܺ�4R�bm(]�%�ta1;���� �;�{~F�1�v���*���P���g'k���9jAK��jr��l�;�eN[�E�9��9&���x��T�[EiN����РG��b�Hs��-���1�Al�:���Or��L����V�o�l~fx�ὄ�e��UG�����������P��Y�7�������}n����p�����Y5h�?�u.&Ӓ�b,x��A��`��E\&��)ZO�y�_w
6�i�<�� �J,F�9U@Ǚ��A;q�x�j��u���L���3���C)Q�>����=ظ�vE0��ei5�VA2�9b�5a�b��L��
%��A'R&��}iM�h��z@�e��@��@�[�,��#KV;Dd�%+��Ľ�z����t� W�uuUi�y�C=Ck:����sj�vd:-�{4���t�7�p��S�2�R���szM�'0�~��h�j�$�U��&�hA,&��7�,;T /Eq�O�`��k[y���0%`�2�gf���[�_y������w�����v0�\+������ۺ���<̃֠���	Ʃ�U3���Pv�w�Qd�&�E�q���� �Z�� ��"b��L4��@t<��&,���# �ܡ�o�5X���Au�2�-�b�?��P�����¦�W��1�pxXb��ޣ��-�`�BteX�oZQ��Q�87;;G�i*�~���w�ab���b��}���C(`�ؼϕa;iO�O����s!�,J�`c����m�B���Y�� +��?�a�K�Q(Ts���(�����֪m�қ`3A�ȯN�Ϟt�̩Ҧ�&����P]:��X�w�2/ �`��?.d{oH����Q_�Ť���b��q��8m���b�a~�g�3�Je)�
�,��`&�@+�NB�%e}�bu>����_�]|�0-1��K������K#��$�!s�kk��؝���뎏H�/UVZSO�`+�u�n��h�;�-�^�}#6�Lg!_z��^QB��5*!���[&�:f�e�]�%�a�m��.E��C�����|��x��@�DJ�3Gh�}�^�GL�S���WJ��\�[)�<v���&���U���;8`u{մ���c
ω1��6��אs�l����˧B��
xTM���SQ����KS��	�PJay��>�ߟ���q��L4��U�E�\� ��.� ��jqJCy%�c���"mfj�~9��%^w��#�q#�a⹻�.! ���|>�T�U!��mI@Z��Q�|���IB�~o$Z����uQ�ޗ�Fו�MfqsY4���Р�c5�Dw���O*�	E?nb�k���[�{ٗ��7��{��tuU�՘'�ߢ9}��A=�=��Յ;�,"���N�z�@0���λR�u�$����5��h�1{.���Z#��5ź�j���V��z���d�d��++'�,��K9c`�?_��]n俌��Ւ�L�ƝƸ�gu���}c��r*q���f��k�e�u�@[� ��!��S��!՚�T�wT
|�*�;Wx&�.cb�1J�k�>y����f�N��~]ʤ�&�z��հ��P<��i K=�W��{v�{�_5g(9�&�6��a?�˗��|?�kɣ�v��jbQ=�L	��2���׽J�]6a���.��E�v��CP��-��J�v_>�ݢIh����1��0��Ԯ�K���EJ���T��(כg�'4��۝��_���m�"�V��мʆ=f��+��e�ຼ�R���F��"5�K��2�2r}�͸�G��y��E1�S9��˘�T���jR��z�e4�2;G�N]�3'99'���?��gSf����� '���h6�{��t�ϺD�	RIO�i@���CS%.|�M����bL�s|�w����!����s�K�h�I��l��K�}E��H71V>̕��u������E~�(2� 'ac���j�(>�H5���1���OJ�����+�º_^�1��%9���@%;}A>�-7�@ �Z��?3�p�SI��.�n��:Ԕ��*u��H���+O._�<Qo�&�i�����K���>-D��Nr�`�'�V��>ޑ�#��7˖��b���s�ð�����<z%��CΙu'��,yV�b!x,e��+���Vo,�ǳ~Y,K���@��*}�g�( �ȷ*�:�\_��5�>����٦�p��;�[��U<�n3cתE�C��
�ēr%Hn[ոN�/�|�s����E����H��C�USM�lI§%z:_gQB��|B���b)��p������X�[{���3�3Q�U҄���o}�%X�I�L�^�@�l���w�a"#����sU^3����a`;R0!��ٶ�2��+%�5B6�w¬N�4�;<҇���þ�s��-T�+��t����,�%N)�E�O���<�
�ؒd���6�̽��ᶽ��rn�!��:]���W�}�p��6j	5��&��� Bs_�����̃�ً�����|����&쎏�ܼV|z=�>�n^�@:s���mx"���=��U�F�������*�^�,�d��Tȧ�p6sHC�ښ�J�j��c��P��_H7n��Mo�ؐ��m��<�N0�-���()����o�[4HI��Ǌ��L��=Wj�[<|�����	��K� 
�ֽg���æ�tE�R��|������\�o�7�7���}�läRP�0Ffa`*��aǷ<'�H�$��D���}^��@T��Ka�{��t�kBK9���+���`j��JRtm*�<�y��Z��d��uJP0�f�ペ�Ⴍ��L�o)�b��Ht�w3���#x]������dj��԰7lP�&�۞�^�Uu5��}�Q��gi����C��,�V����~�`���xv��;%(q�����Z*���'��:�Mps:wz���	ww��3�kXb��櫎21bJ�w��]&�"��I��VYx�/Kè:v�߾/w��V]��(����뉣o߸\)���*��=�Fɟ�L���.Mؤ���N�Y*����\0��l��P�a�Ob=A��چA��A�<�?ͻ���fU�5_0˷�Ȭ\d��m;(w��|ifc��R3���a�4���4I�K.�Ʌ��݄O�%���q�~� �v�~��ܟL��|�ǜx_����y���L�m��_
By��btN�=¯���� d*��V\5m�n��mS9,)�%�y�alXm2��G0�A�A��b�<ޝ�(��3�/~��� ���J���/`�������uO�T�%*:�E��f��bGEOD����*�B"��7��r�J���\�7P����t�Yk8\W=��ܾ�+����l�r��m�*��ꚟg&>�9�����%&5Iw���RV��b��3z&9X^&t{m2�K$��o���m���ec����r����cD D�����C/���5H��*W4�,!�S�!�Y8yP]}��QV��!�U���%$�w�R���0��-9�$8���)ǰ�����f�ꍹ$�H�����a+��zҫ�s_3J�?�B��==��QJno@K���3��q��̃A��GG�V�j_��;���I�F	l�r�G�М�3���I�Xw ^G��yQvqE�M ��>��T�G���ݕ~;�����Z�Z�^�����'�J��1S�k���Q�Yu�|_иp��d7' H�WT�ڹ��﫪�F��5�d�������6¢��ӵ����<p�\W��|&�5�T*N�v[�b�V\_���O��h�l�O8ܶ- �%t,Zt	�[X+���v�����\?�= �u�(�T������S�4-��~�+^ա��~�����ctO�ſ��lc�z���JJ�L��kEO.v�����#<���u��$���ݚ����O��G�ie_���?�5�|�*��.�{d�[�O0��b���;5H�WH�	1��w�]�'�l�ȷW���kI�0���'�>2Qd�y�����ǒY��y���rD*��<~v�� ����Cd�#ث�f&rb�Y0?�hL�ި�����<f�����?,%n�����ߵ&��-�iAz-M"1%�x��8DV� �m�nJ�F�á����o������N8��f�]�Mk7_R/z��Z{��͕Fx�������b&r��+��U��ǽ�z�ܥ-�'u܉��Vs	˿�MƬ�&�pYl%G1���cJ���L��	����l����W�sR���D������N9J��㬹� ���)��z��=n	r�t6�&|�=�.��n� �ͬw���Z��*�uz�j�"qK�v���M�h��@X�ǽ�׵�o�TV�szZ]R)W�8��,��TWy<��;e8Uz��W':��!�P��0�hgۇ�*R�EI��F�/n��̖Z����K�N0���ğ}�ma��R��at5~$y�7��s��Eq���4��_����.OE�<��8E��YJ�nȣ\�D57�k�W|�h����P��=�J��PV���:Keh�T��6�TS�7 �����/���פ��*��rfPi�L��l��{�^\�	c�2mour�Ѱ���M]I�3B�ϋ&�!?��h#�&!c��e*��OgD�4^�J�����������$�jW��$p�љ�%���ü3�n-��]�mq�IRLUQ�N�<8q�#�̈́���_��_���<~��M
��l��_�C(���7�>�V�0��*?�׷g%re���6������ߍ��3�"��B� }�Hb�����a��Ǒ��z�������EY���&��`��ٖ���}̊:-�LƫyH�`��{C�l�_�׽��e�8�G(�0jSsBto���jk�	D!��=���]��7X���z��9���f?�fw�ɯ�-��B��tƐ���v�ߨ�;��ڪ��IB-�*�I"��AJ�&�r��6������oJ�ZL#�[~�C�/�̕{r{�<�/�|U*���\��'��������j=�@_�����0����ܰ�e.BC
?����H��4i��M��S��X�f�82���̺�6q���>]�v�$�-����X�]�U^�����|��d�z�I�|�}�Uw�����W&	�X�%�w���#6QlˊK�t�[Kƻr�����u��Ԉ�m��F��kZ��t ��E�ʐ_�A�a�AA�7���Ӹ4����~ޑF����a������#7��aߔ�x��z������(�-�tl�7���`���,�b��P���F1慭�b,5�ݳ�>��O�7FڏWV�S���\ZXX�0�#��"*��~��ƙ|��x+���,\Æ�c�K�Z��&׸�jX�]����� �_MԟM2�_��#�u��Xث�ǆK,
�����wO�HmH|���Jw��rf�����oe�}��Ȭ(���xJ�hM�����$J"��aч8�<\�Sؽ��.�9nl1X���@df��o&.���l���{��Pq�6�2����Gx
���n��&�����1(J�0���1Qlu���l:�e(��ak)*���&Q���#_ӁEǂV�?�\��Э��
��9Y�~=�p�l���q^]��~�az������dvT?��,x/!���/��<��1UUcee�v^$*�[��X����j]Xۉ#~-%תJ��I79�պ��Z=�.!�w���K3�Xy���y� ���/��un�Y\���&���X�Y�4E�����cu8�-{�`S9�������Z6S9�����3��S.U}���݉y�	z�^��k�`)��8�
>�ޚ�?��m��~��������@A�k�<�U�5+�1�*�=#D�}���!�,�8�s|�i�D��VC��j�ԞUt����݌����`�^��s�� YOY`;K�pФ�CN&@sAt�%@�5� �;~��DZ�iI;�����Ӻe���g��{�N�S�[^��x�d.��LDkY���M�\��>�������qN���&8>X����V���T@$�٪Ȃ��O�7KJK��Y������
����������1��\�����h���Fգ�v�[S|�J���j�U�����Enf�G@i�d��ԃ�ݽ(��J�^pF9>�L�>�2�eJ�=�<���ka�]�J;l�dK�R�\�Yb!�a� ?Ĺ/__����UӜ<y''ϣ��(v��j�є����^�O� � �)�ég̚��g��Q)_/�m��y�]u�mT�A�ˡ�	bQ�����u{yޞN�|�mS�d���꾋SP|H�0AJ6<̴��Q4'gpP���nj��mL���I�`�=Ɛ�ͣŖvR��"��`Z�n�M�v��od\�fS��0>��<�I'<�����I��� ����#��<(�~=����w[Z蒰���ܳ�a_��9��]ɞ���wr���b���^J�,���l}��z��:1�i+��t9��qdq�5L5��/*rk�ЗdhV���(�d�@�H4XLV��lQZgs
bE����>�}�=�����-��ѿ�F��6 ]�'����?���Nv���~W�tz��֛�}ˋ����'Y6���o�Ȁ�fS����?����s����8��r�غBi���q�B@��@���\�;�n,Ɏr\���W��K7}����,�~���Z˛\m%����g��,�Cwsu����^Y�����9�8pc�N}��żN�-[�r�����L�BE�;y���"�
PX���B$������Q.��6�6��+�zi��.�+˙3�g�+��Y{F�/0�� �Z��"GLt�����_����ln�O�Ξy֯+O%���}��[�>%AQ�����ٱ2��L���MI
pYC�sȻ���Δ�S�m�[O� ;j�bD}����6-_|����`�Jû�ire�
�X�z�eQN�`��c/���=X�)�9��Z#�֤A�����o
���zs+�e���D;�0�t.������'3�49K���+t�Ţt`%�Q���ZO~P �f��k��R
u�u�M�W�i./f��4�+�"5CY>��DۉM�B����4g��G����m &�QVX5$~�~|�ָ�X�y�N�)�L�ԂF���̨��n8g�o��U����1�҆l���<���E�m^8O�^��m�i}#n�ڛ���Z1ڬ�9��:�4B�b�r8�֐�7�ˡGv�sT�-(�U���(l���\�
�'I�UɬoO*��ҭ��q��gU��M�b]v�Ӟ[p~�b�@�r� �C�QK�j��X�4q�Dj�R��6�*%2�$H-�/��*�F�����+d�_�fS���dy`%����O�wY�X�ų��9N]�UYI'.�zeE�����ӱWڅ���p6�G ��L@���w�]Y��o�r�(\?f�.t�eq�2�]'K��[������s��%�_~�Q��<�R��nU+�74!�em��Cp�ⅰw���j)}��/ňy���TI�>	��]y��?�(�E�$�pK��ؑ\n�I����[bEyW4��,�z{
'b�Z�╔��z�;5�JԙMN��6�J �ejV>o��&���#]@q���r��6�I���_J��H�{���b���PӍ��W��*�Ӯ	1�4mVz�e��ë�o� i2m��,ߡY���x s�kD���]︪�`���W���*�^�-��0�F�N�CV���_E�!~�m�U.�3��^exU�nA䟸a�C��Qt$em�}�c�V���N�SG�Keeb�K��n��ʩd��핗y�,�O+G:^�G��$Q��s����Nǉ�U�)���(��#1���*��H s5!�=}�{C� Z�Z�R�<d6� m�J h�A���՗�T���:nؿ!L�w��>�-2����d�.î'+���A;M�o�C�'��*�|��m:����a��S��,���IC�����xNR̔]R�n��aE�� +��|�!!u\�wv���2���b����Yv:��/���u/�#v���;S�T���̇�<[�?/[Z�v��@	�����k.�m
�N[j>�d!F�P���`�aܠ���W1^�H�>&�{5�1C�p);E������g Y�\&�r~F���x�}�Kc]ڢ~J�N�X<���Qs��g{�/����TGg����}ӡ7~؟�a����F���M���DK�:W}�v��kpM[�w[�Y��B�&�7����V��)#{�\�����%Lg�$��d����	)gZ��+O.���N�� �訽��\>5�Z>��RG�RYpN�@����mv���k��Hbc��Δ$����(��7�X�P$�����fzs��U���z��CW�ݵ�f�Q��~ܦLE�TV������oUcl'ΧnWk:��$�eq�����5���ɴ��T��:�䊺�s���3ފk&�F"~�{�{����V��>|���1j)��7fP\=���Y]!������y>����~���I����b��=:�s���9�2���A:�ؓ��W�l��wܭ�]�S�i��}��.՞��Q�+������3j�&��Q�N�_E�̟)ڄ��ǫ�{����m�.ͭ���D�]���DE0��"�N�I���L�Y�<b��!��¯�S��y0���'��L��ލ���^�Ma}���5'�j��M�����kw��~����I�M���qg?a���Q��4��|'Lzwn�`�{��|��<;ۀ؉y��C���(��w����YxL�Z|Ǫ������òjֆ�"�ۯ�ϖ;��P��C<s�����uu&ԕ|�6�πƲ��q��P�����y��P��w�e7���`5Jes^�;���m2�T��j;;������b^����I�^�ގ������H,��/z��,3��I�%$?�+K(�~���{3=	@P��ю�� �w[�_��o �s�u>��DM���U��<3j�!t�g���d��29���YG޾�/�=����ek�6h/!����RpNN%��������5N�]m#H1��:�sD!&N��.��pc�?��^R��äH�S�!u��ABϦF芠w�����ɝ�L�o9�}e��9��iP~�x����7��wx�9�9@4��]��5�\Oh�'A*P"����h�c��)q�aH�y钲�Wl����})�[=��zMq��VJ*m�Ϲ�]t|PZUf���.�?ҥ�wb?�&����e���9/~~�faHLAge?�S�
hKZ����^9�":�)e��D@�vr�d�g��Q<L���p�>%����ø��v."��=��A�",̍0��uM¡i�UC�cɔ�~�ܤ������a�֏���W'�൷(c	�G7H2�B����S��Ki&l�}iwD=;栟Q��1���`8]5u�ޤYd1(\�T?�F�ȓRЈv�r�tS����O���1�X�1[y�5������}����5)���+;���Zk1n��)tN"�l�v����m�̧aʵ�[9r������;�ߞqr-��R6{G+Zq��ɢ�$�����\<֟��P��PK��:�kC���&}O�E ��=�[yQc�h��ǆ�]������C�n�O0��qR�����8们�3��Q��j�d�M�Rd𾦲���%>�0��E���]��y�<X�oc���n� >�9𥘱>Q��%���f�����`�O���������b	UJb��jd�VI�4)@�?���0xMo�ۙ%�~��x�
�0�ݲ��-_�\�<������y��J-��AQ5V6�Fs��-�d�U�e! ��x_��U�+"!y�t����$:J����K*���O�u�f�edul�%���o�z���C~C�L�~E"S�����cz�����	�E�/���	z�9_��c,rm-�	��lԘd�	|I��2�IĭǹNb�/.-)�H�ke�����!��b2���`��0{���`y�
�����NDx��s�-��XVƧϷ\8N��p���cNX����L�}sE�I���WlN�8�z�\`�����?��
G���G�ޝ'g�^����.g����|d�z8����}�V���<Y|�����<c���X��bo�$���hT�\���2��M��	y�^��V���O�w���Y",n��ts�U�A�n���m���dF�
��ۥ�.��	�mz��2��/��m,R��_<�m��K��9T�I�ٜ:�������S�-qR��������L�����3(0����P����;mN���U��G��j�o�bz�	�P_I���/�<�}���� X�E�o���楕ɝ�l�23��,f�~�'��<^����:r��G�]�u�2�k�6 �?̬WOl��K1�ђan�[c!�0,�� �J��	�c���T�B_l�]b:PZ��Aa�,;(���7��6��I�7��;<2��`:�:��#�$*����柝�0���ݮ���1��2��B���}&�m������GX�@' �V���gYMر�Vg������=mTe-�8Y�@$��w�w� ���W��I�\[]�=n[��y5)�K����5TrӘLXmWCU(�z���{~���b����?��n{F��b�/u�K��M?�T�7��ݓ3��<#TP]Qj� C����	��m�vCj\�©�F��{&���I�Fq�|��N���Ft�+�̙F����*+̦�i�Dt ��βNg	��u�N`V�_,>S��Q�:ߨ��)�SN���j�Kkf����%���زm���,��|�α\�@���`'���DJESr/��㬸�"e�|�'�����],�[*V!����ͦ�9���Kg��Su�3��F�3�!�-A�bG������O �4�o��� pPw��
�<J� ~|�ۑ�¦$���^���c��FX���T�Dd�U�����)M�"z��C�-��J��:&�0�F�������z�����<���Z��(>W�f�����$
6g2�y��4D���W�q߸�'�Z?t%Օ�"��� �s���2#(��&~B��ͻ�t�Xz�6�8u�����7G��OT���!�.�O��;��G��_0h��-�5��=�n��<�ӦB^��R�Xq�X#�C������@��@;�w5p�K��\p:���ixzy%K��~���=k�6�%�6�ib�~��T�����X��˗�ﾸ�򞎺`��~!Л���Et0n$��AL�G6��IƊ!f�G��?w#��Y>M�?�cӝ?\���ʩ+�M�,@���Y��J�{�m��1�C"e�r\��Og(��96�к�Jo�lŤD�9�H� ׆)7V��w]s�Rr#��n۩꟯�'��8��H�]�Z;
-���ҏ��a�r������������;����GYb�&gG$O��G#�g���$ ��ba����n��cO�/�k�<�mX�	yq�=��T��ә�}��������c�F2�K����bcm-�u�eA-���xD�p�|�-<}w�FU�a"@���4(�^��q*N[u�$�����J$F٥X��=����M�:8x>ZQE����Ǩ),lc�?u�����H拰�N*�a�t�s�t�c]/�2�t�}���88!�����O�	�c��TNn?E�<�`h�4�Yv��m^���h^�iL���a�XlH*���Ӿ�_�������蒝���u��+�j���Ot��O�C�Uc����`mG��w���'N���}�Α�|�R�t�N�Tj7"�7�m�+o5H^`�~H#,B��-���>��7��-1����6=��}Qg�J���]#�s��;�ִ��L�H���SQ'G�V�U� ��>�6����p�l	����X<�B8��7�H�8��h���
4�f�3�m���j��fڔY�c���6�V�e�'ǯ@N��W�7L�cA�O� S���`�)>�)��u��$��Q���C��|7�#�Ϭ�E d������nX�h���q��v���B�3��E�O��u�ylݧ�������S|��e,TZ�zPN,��lw{n˷��Pf&rf���nS��\+��--`���O �=ʎ��6r�0��B^���bb$��7|z���-�3�5��"��H���[ۗ���l���KQ�b��g���<{��y�Q��w^aUA^�׀���u@=e.s��>�o�q|Jr'��re�����B	�^#v��q����Db�K;�J�G�CLI_Xh����b1  hFw���%�dBb�\+��o���f�jQbn>�ޛ�����t@
�����.�g�;{N+�B�݄�lh$�?\��Q��VuAq���N�x[d>�ز�v�%up��������ˤ�.ͅ���ls]�4�mƛ?/��k%�E��T��f��yK� �?������0n\�n��r��!��(���yR����7�Ĉg~���a2����s�5먑�j�̧$-�?�]i��/���eQ�30�.����f�����麼�d�g"�ϲ����M�~{Wb
=t>P|��5� �̎7�ۯ�n0�m��;�+�[& �y`?�:ۻ@S�J��M@�gx{,�9چ�u��k�om��	�)��C ��e��Ϩ�,��҇���#.3��@,U��|@oNf[�TR��f��P>���~.��< lΞQ|�놋�M�,TvJ�Q���H���`�V����mg��"|i�ǃ�4��� }���x�`�gKZ3���f}��?�,s�㵋~��G��u�{d�no�&�wL.q��Rxp��@�%����t����t��2��ϓ#'��4�M.xŴ:�Z�]������]5��x�*���'do���v=��
��q�q�5(��m\/'�&;LB�HM��T`���󜏇w !<J�%���_�/�m���e�l�m�W��6_�x1I	��[�ls��F�e��*��0���?�8��wM� ��5CO~�4�_����P���:�J�����5�0�h-n��W&�>v#CȒFRT���FJV��:Τ 3Z�}�~�7�3�ܡcu���	G��&F��<7��jþ�d��	���!@�:�)İ�r�_��~�ָ��_�r�uw �F�u#ٜ,�(n��|�7I�xv�ʼoe�7���/��w�7{?�� se�9��0Sg6���`�pA�(������G��r���`�M."�g~�w��?�j�H���4�ۼm�J���L2F�"U!��]I�Q��5qj>/�$��9b�!���t|��,����@�Kj*H�4�j�\(����ܖ,q̠:?iN��V����e5��xh�������ve�N��S��߯6��f"�=(S���ӓL��z���3��<<Z��{�s�O5�7k����Y��J��[K�� �oJFL~涹rZ)�a�BL�ۖ/ct��)p֓p+gh�Iw`��+t�<�j�q��A��^���+�|J�;ĹO��M���%�VS��\;W0#:M���}�BF�Á0�
c����;6Co4M�� m/��F�#����:��<�5��KXl8�fb�Tj�4q��m�!�f8M���G��mJ��c|�'_H`�_�/'�OtAΦ6���}燥�����_}{����N.��.h>*�kI§eup���<��+�,�b�.�&~�z���o�>[%nu0���q&ƺ�GQ\^�l���k��N꿋`����,8�cOL>5���������������=��~R�.�Sѕ!��Q�Z��w�r�͟�T��K A%Di�v�ȸ����P�4O�e�)�Um�������A7e7���Z��Q�x���w�4������ן�L�cS��67��/�
o&��=�P��X�'*}���Ϩ���n�ʔЇ�	�v[�q����
cw�{1V"�Z'����=��U+��v*s�Eu,��`u��D��>��-����-<OQA�R���>�w���n$:�k[[��D����{�|
����ǅ^���`~��u�GU���(=�M�d�"����J�o�(e�v��y�6�G
�N�Iz��;�v=��~j��������et)1�,eI�<B�*ԁx`�3
F��PQ��#p�"b��_��Q��Bל���|i_�'d�E����:%��'|2�f�{�u��ӎ�t�1��J����s�5�����l��"�)C�K�5��'˪���M�s��to�D,���s��r?�!&���M��ڕ�_�>5�=�G�.���	�\��'�%L��o�`R���F�q��r�%�QI��7Jk�D���&�w���B���I��i�Jt�>P �mA���f]��^W���o=S��Sǧ3S������J�e��}�ނ�_���; (�M`M���?��?�,:p#j�Ika��Uu�{�� �`�G�xa��b���E*fJ� ��1>kZL�i8��Dr�5�2���;�6��&q'&��u���[�Y�;}�I~�GT�By=%1�����q���wO
]v�e����t8��x�H�^��F/�=9�&��~.|��͆�4�x����Q��4�p*y���(5�6S+Rx9�Yg��*fKp�m�=�����`�jquK�1P����şg����sE�)@'�h,���I_h��p��{3��	��{�"��n���6d�&r�k٭v=��X>D=V^b`��?�ƿ����(�"�ֺO���~��� �,�N2?O+�˓J�bL5$�r�|�}�#����=X_~S��̜ Mb�P�q]���]s�]�u7��������.�S����UP'
;�h"�M&{��}��Q�R�Ƀ�:l�� 
{^gC\-�n�}�F��Ӂ'3S�A�v�D�k���Ɨ�Nf�O�z=�1S-�X]��g���ӝB�`m6�6�C��S�}��E����NĵNoԢ.�z}M[�0�v�ݤ6�`sp�T�I��o#�yWB�&>rw���V51�2?t#���,�Q�Y'[C�x\Bn��+=֢�H �����~�}CD�ݛB�h�'��Q�1������_��v��Ф�������s37� ,r�^H�r)m����������Ӛ?������>�K���s�nr�޷䣈W�xő��v;���	�h)8�rX��Z��?9��y��U�OX��b��0�F�lF&��	n��X�	W��jt�t�`$#�G߆�	�]����=/�h��ʲ��]��fI[>@Pz?�:!�bF��ڍT\c����
7bm�$2��;��|�/������ș8a�U��U��*)�/���G�B�,uQ�s�H���5T>�5U d��!��Fv��/�0-�"P�{����$� ��6��]B&�u'+��)�����q�X|�Zxo�Ԋj
D��m��L(�`�.V@����5g�_���^�D؟��m���%��g3֛D�H#dWx~h��6ݼf�.\��v�W�c�-��,~�EU�>�WWC��0N0Co�sx��l���f�l}rI\b�0�l�,�&�AW�'�/`՛� {�*o�i 9��8j�����_�a��lJ+U���K&:���VA���<�S�lҴgB��Ƨ���l���K��k���N~y��D��5 W����6I}�@i�y�x�xŠ_ �L��x�^�U��˨?��HB�+zs{��̓�@�����~Y���c.2��Y���UllY��s���զS�<��=��xt�"c3����i��^Ƌ�l.�'�@T�p�������-|gެ1ߵ�"'��)n��V9�k�E�@d~��Z%4�=��_��2[��?"?1���Xy�1#����~j);�nV�6���ߎ&�H� ��r$��X?�����'�qҚ���v1����e��Ԙ�_��N�Ժ²�����[�@��~��~�s����%/���0\4m���C��khb�*x5�pR��	�י;�]wp_4h���(��VZ�-��������3G���-�'�`�*�(/W�:�J7�2�\�������[�<ֽ0w^�E�`j����랬��t��G��������d��p�yy�aS1h�_b|�ox��;t5�PE�n>��Sx{p�j ������V����f�5���ss���'��i��`��py�B��41�	oX;%�A������֥��I3�I��pv����,w;y{���0L��ؕS����'�w��zWCan�z�B����+�n���Ƒ����6K��=�o�u�Ko�=��k}�����1xq�R?+�E�<��6;���M�������}A���EGe����Ȳ����#������w��m� !A���&���0����z������R���b'�ͺr,m�8-s�������b��&��6��m��#��iA՛!>�D��mL�9�3��h"�Z��.E����n�����Ƀ�����e��^m̀h�0C����yB�G������h��q�v��q��ĩa6ԥ"u	�8-�A�rv��x�X�+ewE��W�����^�������<|'k�����%u��λ&i寂T�
{���Z���ƭӉ�23�\���jK����P����"�c�dR/=�ߜ�6T�6����$�%���ɔ���*���Aa��pY�!�!��)�K�ϟo=-bwf|�t��n�᭦�α���<��k�ʱ�c�x,��-��1'�����Ԍٴhu��G|�����ՙ>�>�A���h��FG�[���IsC���7��S�飭�ed�e��=!:?��躛�)����C�w�5u�m�Z�V�R"�
��"#�
����
**� �VA@��T�2e�A�=��V�����|���}��O��Gr�{\�u_�sN�3N_�M�'�[����Gܶ�ͤ��b �M�����Q���Ƀ�C��ov!��g�yt}�Q�sxo�oQ��;�˰���G�������8��uKFS;S[}����(ë�fPh���D��/��e��g^5�5.J3K�~�AP��P3�1��Q���gY2UVkZ�5N�G=8�>��]TXK|<��g}
�B}z$��R��{T)
|��7��\��o��k��-�c�7���P
j���[��vd.����~��֤��?����H1����2���8���]�kc&dwg����O8�?�:�(��/����T���v����7�����?Ӕn�nu�3<z7�SK�O'ӗ�"��&3���l�/�j���ƺO�k�@���'(��\U�
4W#	T���Mx�g�|zj��4uR�im���=�/�O�Ĩ+�}WMb,=n������*f&y=ƒ�]�."��o�ٽ��"�"٣����e�ј>�UU��'��o�k>0[�,8>�Rx�z�z�� �3v9�>:yu��|�.�]0yw��Mn�\�����X�7@}Oؖ��ʢ�?l��ڷ���e~���+4
�|ha>�Ac}�f�"��A����+`�_�:l�H'�'*�?K�GW����ڨq�"T��ff�F�*�.$.���a���?+nL5�p�OɌ��U�"�V!q�_O�����g����?��
v�����a��p���� 7��V�s�
�{������XI<�_�Q��-�)0���*Q��W�{��7�N�H��QP����(\�N.p�2���9����i�WiX@�6n�U��t:�BN�N��}�a��ċ�z��=�6�`��Z����|���&���k��`��ƞ��N�<N	��1�د�~��B9lDN�q�W��%�嬠A�e��qD�~��ÖW����[���F�\
���k���D���5������11�Ig������|�4J=�!*� h�IU�c���Q��4�B�`9���,��*�"�=�C�5,=c~[#���r�Av�r�t��-CPJ�n�!cqjG���o6�dV�D%���'���e���G�9����ŵ�	d>��~�0�u��k�M�Ŧ]]Z1��t@�$�8��Q}/�\'��ɵ�� ���aa�S��#�I�kl`���A�&���E��bY��
x�#�Dgǩ	�98+X�6=l>p�8�`�{�뾕3���m��R���AD�}˙��4)DP<Iy��S�W9n�����J�o0��4u�M�PC��|r��3l��br9�{I�	��·�~�Č����O�����HO�	TC�>y�o 2�X�����(|��W*/��T���/�����k2����J�T�=���m=[Hf�NйVX����a�9���	��"�]Y��o��{��UJ0%6C'�������>>z�S͇?x�fg�z����}�"�g~է�οd�;��>��( ���3��R�PC���~p�t����T�,9�^�}��B�x�Rp���.k-֐����:�m�;� �l?�600PI��d����_c���Ke�c뱜�����z�<@��[�d�`J�1Pʞ�cpG��8!A�+9��J�n-�a��g
��9g�jT<��U�_r Z���e�����+ފ�?�S�ey����X�|T}2g⦱Z���ӗ+�(tk�,�hc"��y��>��G�{Sxs��(�]4yc�;�>C��w�=P���p�93$RX_E�:r���+v����J!��wx_��آF���;X��D�/�����o�%U�4�,�v�����v��eņ7�x�QL�	��~\ �AP&��&gv�e��1��ێ�n*6�ԯ��������a��[��{w�<t�<ZnL}��|=y��Y�	~$��\�����+t"� 3X�;M�m��t;��7jS)y�v�k�S9q{-% �����g�}d�,���[��6��:P>]/�}X�P#f�V�4�ZL+X��w���� .�&�%�C�����W=UIp~�	�+k��N�I"ӆ��/˙ga)_YL���i�������s��u9A�Q�sG�7�s�at�{�&G&&�10������{��,@�����?�~��Fd�b��ẀPT�P3����{���շ�Ru�|��gzh2�,1rY5q"��M�t����Q&~�ʯ&��B���~���g�>�̇O��e}V�2'�YW�A�{���{�`ZI�F��ӂϢ��U����ؑ
�*�Ƣ�n^���~wh*��9��_��}���������o��ć�jnmF��:�D|��We
�D�P��w��:��*"�U��2��%���U�nc�MK�ح��^�q��I���uG� �^�hX+�a�������]E��$��<�6�R�ɫGz���3|���K������֯��`=]��mD���i�b%�ͩJe���rM��Q=ޅ�;Fc	M��kgO������QK��d�J�X/��x�P�D������T,/�*���%H�ϰS1?�wpC���c$��.Z5��F��k��7^0z�@��i��� �m�ZOH�s���<�do'H�8�{h
�+L���l"���UD��mp��w~�dT>O���}��΀�t%���附���Z{���Le����w�t��e��@3?S��U+KtG��jHY-���ihHb�c�Y�#�ذ#,�/i�v��و4�\ .�z�uE�
��q���T��v��i���}�q>���5Ųg�� ��Un쫎]��l$(ץ����:(�2q�.�?�D��	{7U�Yļjji^ș�i���é��s�)M����M�f�O��}`��܀r���~�p���#ܩS�_B�'�B.�:���:h���rz�P�3r}��Y��2��)��vJ��ЇVǹ�ꅺr/�Q��ca�o�ԙ�M4���ҝ���y�wʧ�f��֖�R���S�^�%<�
�"��v���}�T���q#�5���(�Gk��RB�ڪ���k�>�O�� ���f�	u������t����ky|@A�U>�IWe�5�b��JJ,�j]9�$�w�#�6��2J�Ŏ80�#ԋH��"���%�B�P���6���U�J9(d�˱�V����6�}�.7�MJw<�3c�I�9rKպ|FWz��wh�Ц���+�Ğ�i��
�toF��*�W�ڴ�@@�F&��aT-V�h�!(%��X9�lp���I��l��"�f��~3Z�UM��%4�(���:��N>=�h��{QA�Z�K�8���0�x�A[��d�(��K�>�Ğ�)�˛�t]�,԰��@�˝��~ܒ0�p��%gil�]C�Q1p�Ɇ�F�k��H"�g�%�!"��N���+�U����D߉U�^�yAk�}΁�z�dj���F~�O���\���!^u�'��0���^Ԓ�r�� g�8�9^UEq�D�r������
����K���<A��CWA4��ze 0Y��zw�fZ�
����[��c}�&�[JR�Ry#s���s��w����4��4�S��H�t�U����	87ŗ����c�'<�Yj?���o�;Eo�O@�P��z�Y����,q� nY�ǘ��ۯ�l���kM�(P߰�����d� ���u�K�]d��Ʉg`���I�2��u�m��O���r�py�t�#��ˇT�=T���~���Ь��?'�bϧ]��:�� W�)V���f�5�����cxfbe���)��Q���˩�Y�8&�a|��o\��2f4
|�,�	uǘg%f+M�[Z9#i �Qvy2��䦕b��:A�`?����ѝLW��(�K����`�>�����uos�,}�܊zHM�� rE��ruHN�2ٔ�n�y<��l"_��xd�S�����W��=�͎�@YC�ƨ>�wl(��<��Z����Z,���qA�����Pp[E�h9�[Y  �O�����fq���{$�����r��|G�U�R��z���p���a̕A�+u<yF�|�e�imoF��9�0W��]9v�'=�Szp�~�JG��e�X[���;��HFi0��C 5��.�$�	����a�<�?�~ �J�W�8t���SU�������H�W�<kӌH>V�� F��U�X'����qb��]��w#�z@��f5�����%���{��O��d�ꛆyL��ZD�u|����,'I��0�l�q,F�2Û�u ��&���kyR�ֲ�ˡ�2@j6s�r`��ﻻ�z���,a�4u�<�E��E����]��:R2:M���]]JN\��I�h���^�'�a}����ac*z���oMmq.�H73�j����dv�)l����?,p��k�o%;,͊��Sb����p�U�G��r��&~�Jl����G?�D���W0hvs��p�&�E#��rh.�%�g;�`�'^=�;�U1�����Ϩ�-Pz�7=� >�d��A��c|ZB��I�e`����uD�/�����JƼȜ�VO�U[`���	7B��Oϸ�^Y�*I��}w�޿����޴����&��>*�ޖ��;oI��+�UW{-L��`��D~~+�R�~D_է�	�'��E7���[�*�j�˧5=��R�q8��Sl�zOĄ�wk����5"c���y��-�#o���C>�|��|[�����[F��䅓��I��r�jߏ4�Ӿr=KB�8P���S�I�h"�4�����V�MU��c�;��3�/q�9��_ }|#�%���䷩�8���^���G�b$ac���rN��RZ��L`M����dUTx���֐��R���JQ�D&c/gtٷn/N<g�D�e�҈��{�Ti�wM�! ��GU��9V�ڪDU>#%#
��9�$�暛�D�XZ�����^P}PCWHw�n��Q��|����l�Vp�)���P���{d�!�'��y<R7Υ�E"m��]-����t�o>�]gt3_ڛX,�@
��������[�ڨ��(��(à6a ٝ߯���]e5[�"w�#&���OX�5Erͽ�C N�Y�g���]H�������Kɟ��+W� o{�hY��Qb]�a���/c�~����,s<4�1!�9){8	��YoE>r�n���T�����zeJB�p��#&ng뢈�v�q��]�����z�-��Sg��iBl�"�Q@)���gU��f$���}w_��Ŧ��(b��g�H�X�%���V���@�7��Jq�N������%A����u�2�F��+�+|`?���~ĿN�4��5 hb���(���^���h�Eߡ�\3�LS�3�|�?o�!z���h�H��.?���7AuwX�#NV�Y�,���|�0��	˪��Ikau��������#A��O�d�y�+,]S^]a�%y�&�)R2�z�r�(�#����Z� ���kA#��m��BC%�2�V��P/�X�t�l��O�G��sE�Xye���ҁ��Ȏ���$�i��Ώr=i�{'��v�Q#
7Y��:w�cѧ���8�=b��\^�-(um�std7uA1��d��t�MVD_�N+�Nq���k���XϖL�q�S�8�>�,:�cߥI��N��Q�
������+C}gT�|i1���|5@��D����:��#�w﹙z�!�*�*��`�H��x[��o]�|���l�
�+�!n�� �{B�|I��Q��@$S[h�fh[�ai�>���B���:���u[a�)���rh��L�6ϭ��9���i�u�7�+�G6j��B�
�+`���-2��W�����z���؁B���lp%R���>,L>�U��琹�윌��(hu�4��툶�ӕ>2bҁɯ��.�68f���>����gͯ�[۶�A	�]�ĐGk����\�p#u��Q�D? y�_g��ܖ?�����(@R�i�k�l
5��
�
c+����|Ŀw�P}jv#�U�7���m���/w7�q&W���M q g�Ip� �OcC��go��V���	cum-��$��K������8{.�F�����L�hϺmk�8X����چ�+Jq��|�O��D a��6Y=ۆd�?���	�.����
�����}��u�C�3�N�	����C�
y9p��þŎ$ܯ2��=��J�fK�di^����ƹ�c��� 	X��W�o,�X��ڝBF�N��K�x�|�X�<&��>!�_��+�b?�.~WZ��N\���6�ͬZ���`$�ѹ�X��4�(�X;�����B�`&��N;��^�acԡ.�Z&��������Z��T��dO��2�Iu��<��h�S۲ᡸC�-���g8q�M8��w���΃�0���+%�c�����e �V��vm�[9�����i������Q�����V�I��� �w�9�s���˃D�����������]�c����?���e�����c����dtO��:o#��	�z�������JQ8�'IGe꿙$v*.a�x����Z����D��:L�-+ϸ��ʹ�l�LPp)w�	{)ly'�/��C��"e���797�/�N�W(߰:��u@P��h^��@��]g�7�Đ�9ŭyQ|�f���sKM4M��w��t�n는��݌Y�-o��F�r��p��N�f���^����������7�8�J�IkcۂD��������"��}���-R���FCC(�$0���\�_6�*~'zs��n �/q��̣���?T~��E�UD�"�>Jt�?����L�4�nuT?~ ��Ð^���u_�Y�,��2:�uѦ6�+4 L�,�h��y���IM�Ҫ�w����]%���c�8�,�ןl�O~1r��e��L�方��{t���w�Ƿ��d7����X����8u�m[/Aҧ����1*g}���X��M��䳖�uq��H�}7j�/����Y͗�UE/h8|�0��&��l���eh%�����DϾ('3���������Y�u��1ߞ�h,e�����G�HN���#�gá�h'��� ]������h�Z8�Z2�飄�	����[�<jd�>���>����t
>�v_��U��:7�G��Q�o���c�����]N�R_�˼�r�:�Rfc�qaywM�կ��T��Jz�˖I���(�l��� ���%8�n]h�lli��5����A��;�?+�������O��m���VϬ<�N>�ݼn�{��-m��̞��o+��R����VA���WxP���f��cS
qu����8��U�,��^�4�f�x� �-N���������\��[�@��L��i�M���V�B\�no�"c}!k���5^H�ɪ� �F��-8K���>J�W����y��M�����Erݷ	H�|���Co�}�rK[�����(*��#�dAh���s-+�&�F4�X�y��NB5Px
�Dq�'"��?�Gb��L�#����8����΂�J��q�E��� Avj議7xȁ�i�C���a��l���n���g<������#�� �7�%*�0ͽ�[CnKo�+Ă�8�&i��>��M�)�,��m{�-�,��2�$�	&g.�i�0������2&�o6ik(�L���E��d�u����ε�ӑ
��[�<x����s��k��G��cK-X�W��[m�=�2����9P\-�V�� ��Zk��Ҷ�ǯQ��zﰱ���s�q}̡�A�l�JɻV:��0^��X�ndO��6�c�n�1|���e�t$*8��r3!��߲���E{F�l�k#��P{z�:~cN�晙��y4SQ�[I�1�Y�R�m7mo��u�u�RvI�n�U������G7XO��S�B {6�4�L@���nM��m�|���4%Ӗ��h&�4��m��3�.���de���VV{��	�(8���xV.p�")�(�h��e<wX�i���~Y�#8��N�y=86�E����n|�a����������L9��f�I�O_9�
dr��#u��Ļh�����e]r�Gh���2H�G�F���+��!�T��%c�q��ضy�R>�|tۤڗ�v� qX}�4����t����έq��m72S�0WVz�&S��E���2Qܒm�TZ�%l��I���˔�۹}��&e�����d�̒���B��*3�]@��=M!�mK��Ih��qsq#��^�6�h��� R���Q?��i._i��f�}Et@����A ����78C��;�V�b�'��a����`]�*l�9�6�^���k~vP��X��Y�r!N3|��4hMc�̰"M}E�Aػ;b�.���<܉$���x���7�7J�s��n�r�����U8�Z�捣5P��2�V�p�k��N|��N}�J����L��Z�X���6�B������C}���䙊��k�\m~�%O�ȅrO�DʉԆ�;nq������ۍ}�e�m���xb�Ci��`6^��rJ��9y�������,�4��*��ݦ+�հ>���h����/�r�7'a���[	�@�_� {����V1�ݦ�H��/�6���4��o����Fz��j�K[��&���]�#oa�u�����_L�)ڋ�ℨ�������և
n���8���>���!��;�!�嗪Dwo��A����ӷ��b�n����FC2"��t�9���a�0�׼58gZ眈~~�Eҙ3��Zä�I������qI�:,x��>����f�J��>�<7ѓ�Z| 0`$k0؄�˥ �'W���"��+���\S˅g�Fr�-5$��%��#������6f��A���?{�[��e;�Q��0��Z1+�Q�ޭ5x��[�(.z�I'�I#*���*$%ɉ�v�\[}��l��y,$��8�?4v�O&ƽ�p�d�Q�P\�m!#&�T#���	y5�T��.S�Q�0��� 6�E��V�2�?����d~�~��Ȱ��jz����ǯ�XG;z�=z����/�|����qr�S�KTe�8y�����r��l�|�	��:�������M&UU�֐_��3u�U�yY���x�I}ai���h��r���9C٫g(D�m���^��(�u g��y�G#�`�a�S���1^��ȣ�o����8�/��B����2��}^��ϰ��eq�<�����w{���ԴG���=#27�:�57i�v�[/��U��r���з3�׶��Z^��8�[i�U˝��_O�Z��EZ�̭�1Z�Ü:����ۼ����Z
�{��&Q݇����:0f`��X�g�6=W|kr��Dq�Q�^H��\��_��Q��m[U�'���	�O,�Or7�c�����,���/�(:9��ӗ����e�X9�.Y������V
�ܠ�{�wN?\m�Z�w�yp��='9��\��Δ"�_�H^���J�o���fn�61�|].�R���'���n���*KH�¼��jjk�=8��=����S!�k��-[
o35�����}�͠D��ʉ2:ͳ��N�S�N�1����U!x�ݪB��Ҧtc��`��ŧo��A��R^7eۜF>)�u����cKo�zQ�2��P��P� ^N������}�_v���c�[�,�����y�W֚�|iWr�ջ��3޽"'3��KQnS+V����z��J���\�AF��L�٭�l�@.l����ܶ�H/�z�k�loT�X}(D(��#o���Z�~!.��]}���zG�M���|k(������{�����Q��6fd+��3�$Q�����݃$�d��dKЂ"�A��C���c��BE=#[\)12�e.�g����֝;u7Ζo4�`Q�W@)�}���,��u�'q�#��a��[M�3�zȡ(+�6���%�V��Vx;��x��dϠ���o��P���a�.l���?��ۗ.ig	�}g�8kx~&���t�%��֫��lg?�:���jK �^߾�5���r�������b�
�Q@7�N�R��=�
Q,���;��������<�l��ߊ���W��P�,��C����ɓ���&��i�C5^�m��l;�j�C;	fj���@o�'|����2��Zmn��C�H �W���o�$O�sF|��������-1֨�o_�X<f4S�ߡb��ײ�!A���9��S��rԘ��zD$��]��i,��z�4���f����C��Ed/�k�>�-�B2�P�}�Fr��Rm9�x�J��1yW���o�C�J��MѣqK��u�cjPs9'��!\,��_]L�kÃ5��iǾ�@A��&�^kI#r�r���9I��S� �]
���P�j�Y���rtG�.����h�y��Iy����㓇IB�Z;T���S?���BQ�h��h6� ����5qn}�6O����"�;��T٣΀�ɸ/����@���^К�4��yﺏ��ٓ����mL��<����9%�
;;,v����G�!}۽-�L颅��W�/ |�Q�N-�Y���dה��t#��KX�'V.)�c�{�Wdz���%KyJ[���Akcj�J������i������)2�H6��]>��m��${���(��H+̠���Fc�r/s�xIX��L�����ְ�b��D��^�JAf��&�
��������*�O	ޚۿ�+h�4G�Z������i:�6u7��/���M70R2����(p�����B^(�S�q�k��`���Xu q�h��M�/KZ��Q�WG��2��&s�'+�k�ڄ�w�2o���@�/C�����m#�֌��&F�Xi��[���`��fa�um���܅���08:��.?�Z��6L��W@!�j�@����Nd���#�iHh������]��'��@��M�������D1C'k;,�m7����'@<>	&�d}�=^(�U´��"���p�
��:��	�tW[x�z3Y���ff ��PZ⡤��D�B�w��� I��"�j�0�����dݹ:{��:j���������I��_�Mӛy�R|��3t`��X�91<⇳' ����g]00<�Nl�d'��mp���r��?��%乙<�Tzf�๭�V�J9�={>������ ��y'O�j9W�[Şw�������\%A/>u��?�vǻqE�v�Pd��HBWu����YB1t&���]�f/OWcy�ipO�|+��ig��\��"c(-�h/8D�#qʖk1��R���P�HI���u�%�%��!��
��{���)����4��z
<W���f�ڻ��օ�*ۉ��W���7�ꚬ�
��<��'u��k"6w��5��nqg3x������$��*�~�%ry�v2יWq`���څ#�8��7%�U���N�J��3�Y��uy�7kA�#\�R���'꺏���u'+�ߨU6�p�^s�V�E9�L�?�L�"��:x(z���g_�N�<ߛ���'ɿg^�� ��;�'s�n$�W�˽Q��@�$��t�'/�C#��+�k h�=��FsS�k�sAjjf����r]�Кᇠ@�˓Vw�f���z؝i}`��p���ډ8L�NQ-i���,7 \�D�[2Y;tA!�/�4>SV��=h�}®�e��׀�O�-��������w�p ������V��O�[j�L�˄�+����od��F����*�
"o1w��b0�tㅶ���w�/�'�qY~S1q;�u��\ʬ���9��}��+
W���U�/����J�L2�^]�?P����V�Q;��-z��ܲ{�ѹ:���2X�i�
t6���1B�����K���9�}b����%Wj6xw|��m������,�|9Kg�Q�I���4�Q�]�y{ΐ39{�CM�����2�fCґ�d�;dgP�|�B�H�!-<������g���45i�l��H�nri������׀g1U0i��&��N�;��6�&C)�]�ֵ'K��n�Љ�)�S��T�c"&>��|�@�qe�,Aj�kC��/_fk���6oT�9����M�A����RT�_�?xvLxӸ_���hs��ݻE�������T+�Z'߾v�|����Wu�2N�ޓ�5+�a��zծ�lb��G|L �;�xEvǳ�n�`�0l�ibD�o�{)w�`��c~���kd���t����5�y���D��)�g�����[�|�j��`_��D��MK{���eV�H#Y�s��.�}`���.�b%F-����h��� ��Y��('�p	��T�i��� ���@%�>��~٦�����y܊�r�r�N]t���0Hcqv���߈ͦ�E�^,��SR�xW�Q��o�xn��9�c�tA��lQ
�2)��=B�1��B�|Z��f��\~{D�we_��b���XK�ڴD��ֿW>]���>1y��_��2Z�˚����4˷�'������QC�������I��"��ٻ�}�	�>jy�ڟv��ǽz�7��<@]\�O�KW?
��%+<QN�V柚�1:)l��7����ӶO�Y8��,ᩎA���	5'm��ƾ�ׯ�t>������ӭ��Ԋ)�2�����z�Pk>�^�ͨҞ��\Z���ȔOQ��۾kw��$" 0�)�|f$^*�7t.����z�A�Hd�����m4�X߯x�TL���!��I��|�^2��p�����%��vu)x$�|ɦz^���{�\��N��@�u�t�o�������*�"��'U��9t ��5�븷�)�@�@Al��	�mओ���}���*U�5����N�g�Cwl��ulZ
I�c�Dc�(;%�N������i����"��JX����L�@�<�@Z;us�[���E6C �2kq����$+�(�ߠӓ�gH�1���"Xk�MuN�p�&�y��äD?��.'�93�x��)�Z�WnL�M�=wO{}dtz ��d!�y��Fy�r�w�̬��9����E�V���`&&k�p$�c��=�eN�0c�\��s�v��"����/#.~l�ư�� m��B?�3�4k��ٵW���@�x;��8u��ۆA�9XA�W�n��C+�t���>��z��bw3Q��w�a��fQ����zd4|%�7�Cg-�iB_�n��Y�cd b�2�=7k��y����b���AjՈ����T��5�Ơ<��|C�!gNV��5qWï8�s������A�!R�cz3)�o�C�B�KX0owN�(��×��T��{�AK�Åsg����������VI��)#&�V��Z6�[�u�KB!N�i`E1Ndj�$��p��<8w7���Ѳ�^�c~�b�=�WB_]�'���KJ:��.h��ɘi�<���^0<k2��$	Q8u8�϶J��*��|�B����ň�fö��*�����	�/_>��ج*�兔�xa����������7)*�o4p-�|xȱm�����d����H"����@c�u���1��~�x�haXDd�(tZS�>X�?�Zƞ5V|�.:��Gւ�@N��`��p���E��8�ۓ��$�=�ȁ7�q���V��R��(�BK-���C��o~�6Ԝ5$빼����\�0�	9xt�}}�u�u��A%���L���	,�<*�_1�ѽ��hCW�>�<�@���B�T�=��S�-�9J|�MW���ct�OZ��m��������ʒ��>�l�k3/��t���M.�FJ��#�4��
=Q����-����:�Al���W�h�@,�l��aZ�����ƃIX��Sj"i\�NS��%O�rDߛ1�5	뼳 �ZC9�4<4z���r}�ū悎�B>��� �$�a�>E�˴�ٝ&�IPeiyR3au�C6���w�=m?'�8	0��|����͌�R(��RSjQ����vJ"ynz�Z��ۜ���CC~���-��%��C���-ȸ(�P��l�ffGDP��UMɔ���4
A�d�
W�4s���Ӎ���@�*.G�h� 4�T/@\�jX��vnz����C��U�S#��>þ��Q;�j��> �V�mW�aF������7��uG���3���B~�b{�Oh3ӣ?��r�DUD8=
j�倴)+�$Z��w��c�zC�8�aF�'��R���r=wNO:B���E����G�z� G|j��i�{Zˬv�rQ�N���nH	���w36��Os	���Qj6E���	*��i�sj�F�F��{Mߤt?V�#-����Vu~LEX!�]-����w/Fʾ�$�t�bR%��l����)�w0���	�[�e�F`S��C�Jtα,K�S��B6���fJ�����_�TF[_%XX�!���>:z�GlE"P-�	��c�ݥ�v������?�� ˢ�R{���MM�]2Q^�G5t�i !�j�f�d�1 ��5-�6��������֪��zX�Ȍt��#���v2�G�x��R�8�b>`����Tp�C��gdqs#���%�M�����ʆ�c[��F�MoK!�[(��
T���H�����o�&6�1�*}�8��b�pV�q��Mk�V X�_���U��:��F@�~~�cԛ�����8�m!B��x�N�%��I�ii�Ii�h����1��eF�~(�h����hϤ�W;5Ly�E�􈩻4$�9��M��hK=E�NSuAH����-]�α�~'�qx�U�A����t�{�!�)��R�6�x���V�ӌ��-NSZ�Q����ٟ5btN�o�pČi6�gb D{�����<��Ԗ����I�53�9�`��lAk� ���7���@�(GI�3����O@��C`Z<T�r2�,>��$�<`a��d�h����K�]1�*�C\�����*ņW{S\� LGv�Ak��.�2`Ā��~pO�$�,O�ʄ�A�GdXyعk�Pn�܀�#]�9���٢'5�'��6��	|B;$J�t�b˺��,T���#,ĞL�.�*w�P?j��DQ8�v�O���3ɋ��t�
5������x)i���~&�&G�N�0M�z�z=���Q ��:�"TC�9P)��������c�C�T�z��~�����T=\
��Wݲn�:J6��q'�mZh ���{Z��Gߡ���ꈯP��#�S��4�ۥV%�@ o��yO�qxZU`j0���h['eX��+=v-��zo���b�P5�͈��Ix�ă�R��'Fr��\��V>�	���ǎ��5�|ݒִ�"q8�43�0�G^g�$q�zq�|��}G��>����Ӎh�����4�J��P˂��K �>��n!.Ƒ����i�L̟��#�3䃮ټY��C"�D`��!NQ�)������Ѣ$5�HQr��ߟ�(}O��NZ`��]��|t����1Ϩ(��n�~�jA�0ҫ�2� �U��� }y�G�&�;�#6�8	(�[�ux�+)�T�>�$�+7U�d/P�N���>���a���V`DE����ݼ ���Bph���z~����3��U�1,�w��S���~�<S�~�O�#5�m���N
dm�����	4�獀n$�5u4�tt�Rz�5�S5�k|��&��ϖ$1R�O%e�<��D�G�vᗦ_<2_5w�#�g ��ϴR��̻�,R'��,�Z��d��J��H�����pqf$�7�(�&�X�^D�m:zCX�γ3�(Q��(�l�/i3�~��ZS1-E�V8P���r���$��BտOwo:l�D�`�R�ʡ|�Ł�T�1���ׅh9��E��e���]5�ħ#�r�O��{S�v)|�RWs��_����	/��Л~k�����u@���:�UCۈn[�Ղ��F��ʪ.4JGX̩ԥ�d�+��9�h�3�R�hA�vSN�eΎ`l�ڭC��N�tCO5��Ε"�=@ԤE���7?��H ���k���!p�x��Z	�%�7/�6e[
gīU}u���?�Y5���R�Ju����c|�*-�?�g�+�'��R����Y�ow/�-�~�Ԑ�7�X9��q˥E��XaU��0�J{n�3���t?��'oI�ݖf=���Ԫv�%(*��Wx^��z���ϓ�tnI����įCP�ҡUU����2��)Yaxd�_A��e�\��Q�	/>`���М}aKMհv�!i�e`��#(a�' ���+�U�I�)�a_L氚��Y/܍���?�z�`����x�0v��ǰim���ds�\[ �SL#*}ӱ9m'��x��ؤ���@u�OZ�n�����s�_ֺZ�땽=9���Bn�������+�FA�궝�٭�{��6ջ4�I�8�Rd�u
 �Aٽ�� �AF�5�Yt�>���z�R?b�y�\D��z�  ���ڧ?��H�K�H�٩�}~K�4�|B�O�}� u	�_yC�M��"(Nc��о����:FZ�����߹�A�Z�E��[�%J������C�Z1��!�� ʸ�Ȕ��'�#����.L�%���{a��nAǳZ�٧����4c�@�%�.6&+�} �Z����h���"����_H��%�x���2bRE�&Tӭ��#�3lL�pq�D)[���n|�m�ן*���XR �}���=��s��R:p�^^����̽���p�{A�F��n�'৬2`�����B��i�҃��y�׽ �����Rb�D	�Rŝ��SuKǕMf��"���I|=��%X�]�L���İ�т<�ه��c��(6�"��.�ߡN���\�cX�MJ��B��55B�d\�y�a��WZ(��{�z� �a1���9��U?t8��=G�xk��ZG�:�X�.T���r��KkR>C�4)]ТA�P�u�4�9i��i�����Ǫ�5�15�`5�g8P��
v0�8T�]@�#�����3i�3�/K���:��PLEE���ao�=;��/> U?$ט�d���j�v����H���K��gl�]�h�ŶwYaVq��bү���Q��/�Ɯ,뒘F�D�Q�_
V�%���W"dwcJ�Ӌ��$\�߽"8uK��bPū�1W"375V�"�VA$L-�1(�[ɢ���r^舻j�4�ܗ����͍9�7����\Tt�\��FU��W��̝�s.�3�w1 �z���J5�W��L��W߶$Y'���{�C���)�^x��W������A?~����)� 'Ѕ�)��Bω�K�j�qp����tD�0NiÑ~��^�O���w�G���m�Ì�R�~�D��S����ғ�ɛ��f��oA��n�&��9ո�k�Q�<��o��¬��{i��q�*��H3�EI�$!J)[�����Y�K�	�s�2�`{/����
#}J3�83rM_Z's���HJD;k��HH���HQ���t�!A���ם��C�g(�F��>���S��Ӽ-iZ�pm���� ����@(��MU�����]�����)��^�e�"��]l+:�u���.�{Z�P$���Tl������aM]��hZ[m��� 2���Њb+�2*�(c�A�[��(SdT1PQ�BPQ�QE�0	B ��a��O����������}�+�Yg�5|�g���I��?�m���4F>%��ܜH��=�Bh;�ejmY}����7/��O�[q�됪��
n�lP�ԉS��m�h��ڛ]�7w�dk��׽|\貴�Yd��U�@���-j��C�e⠅�й_u�|28�|y��S�}s2���smk���e��:�rvHTy��g=�/��(�ʬ��OŊ.�kyw�ls<ӫ��/m͇c�Hq�j�EG�Z���lֽ2'��o� (;:b�� k�p��@�vߏ9�#G��rx�6��	=l�B�'��'aS����h������8�s���M��`hQ��J6�J�J)�1��l�D��9�c�qv�L�����������ϭ�/v�/�r>��i����9�F���bi��%�zƙi	�������f�����,fgm��F{4�[�$����wD��ԭ-j�Vv|��\��ݦ��.WC[���y\��[��_p�*߼��ě-S�����ܤJդ-�E[��Dq�X>����L�;�ې��W�<N� ��U�yZeg�ޕC�[�
����T̏���7��h�f?3-|��@�~뒔v���L����e�s��=��1�{J�Y��U��AZ�OK`��0�i��EO^�������l_�4���ͻ��E
:m����s'ֆ������ZG�$fc����O}��{y1)\�%��{0|��&�`�y��Wɜ��6�:�z���d�o�8s��0k�k2��x��s�ܵ����6-Ky� ;4SS&���,�^殝/L�����{�%jߩ-�a�u:��ȑm�ʛ♃>���9���������^%����T.���,¿O0�;���Ж��33EPĞ柯z<?�2�=s���v�Ѱ��<U��"��Q*tXlp�+۫��4?�!D�[�6�Ŗ**�}_w��۝��RO�ދ�i~I?d�Ie��~v[2כ:��O��i{-�Ś���}i����u��p �_כk�����O=����/�&hs�ν���}jA��p��@Q�v~j��h�1d(9�;�nBU[��T���nm9��7��`���#�ˬ��]��׾�������pq�Hv�ýYy�����	�l�W.�E�8;cWMҽ�of�w	9{~�DŰDf��~r�~��!��y�����u	�Ԥo�b�;͹{�_�7r��{ʾ.����V��Z�t���]��u]4�^q�`70λ�og]_tF������Ӆ<��;�.�m[5�8޽'ӣ��2���o�.O�jf�0P��)Ӎ���C��'�L�~j(k�}�}�77�:ER���~���;�s�����ǜTr䷩��F\J�T�ޮ�����-yS3@���+cͮ��S�N�8�q	���5{�G�Ή�,J���4�j�T�v�"��U���xV ��N
\���R��&l(��Lz�hUJ��#���;��O�+�3U��Q��K�yX�|���!-�
�ڱ�'jS�g9���>�{��̥v��q�J����Ɨ8�֮��`���_u��d��>���gpx��+���\�l٫޷��dC��EL��5������g�n�����/��uM��ph,�S���+o�B����qM���������vA�o�dR��K��)���;�|���t?Ns)���p���;.<��z/��i.{�+�}y;�7���~����<�bx�^�H���r]����.e!����Z��4�8�^�tk�I��r��v����mZ��z�K�ք�}ג<���潡Nm/G��-ͷ��o	���r��hΖr�K>o�s��%�ʉ��-�Z�g��l��q�~�K��ŭ6���s���Gj؄����)I���Ι����)9�)<14��z���ӷ��}i����]y����H�H`^H_E��D[H_�&
�1���Ɉ��iZ�;��o��~%v#ʚ�$� Mя�2����oP��m���K��\���/�~��˥�w/��qBO,P��d��OU��|;���Ҕ/��������Wj�7�Y��/���՗W_^}y��՗W_^}y��՗W_^}y��՗W��yu�w.dK!GdJMA�KS��{�2O���m��K���.�k�����?=PY~�ǻ������!L�����wk�����k����oB~:�����L���Y�~A�����I�Vao˴�̷Y)�)m`�]��qj����}y�˛_����7�����/o�?��?���&?�3��x�3��?z1��]�$��#����X�/o�������k>3OE)�-z"���g�������շc���|֧zr�����8E|�Siy�E�vI ��	������2�DԾI\JO�<���k9t�,y�����p�h���s���Ѓ?�Q�"��C�R"�PI�\6�(�<"�=���g��ѣס��m����z��OD��&+?�<5'���[Lb���;i��Į[HE7�3{S�<:�^���i��m޼9+��f�\��Ku�&Bۜ����N�/�8�$C<xO	]�?���"7��\��g%2�Se��hk2�������n"��ۻnjj�[�siR�C޶�:2N�Nh�:�?��c����+n�W��}p�$�������������Θ�����T/
]7O����p�4鈕���F&��@�/��Z�-K7K�}��.iߖ��Hj �t�M��;c�*X�l�~�\S���ay\$���br���w�����c�}"�1A���8�����pKb�[�1�R��M���J�}��t����oi$jW���g�E˒���^��[D��Ik�=������AcHl��U�Ħ![E�hS���h���2�g��y�s�Qe]�(hI�1�1�q?7���W�g�Æ�>��W�|��pV���^!�m���yMϠ��իW���5�˰�+z����n&,>D���FE2�M�pd	s��1s>���<���tK�pw�@ø����4C^[�*�~ല� ��Pu��}������"�-5 D+w�6T���X9�����ACiP���;88l9ED7�w9,[�E��E��2\�Y�-�sr�ख़,~�DTم[��[0V=K���z?`�}u������-*��*�ΰ�.Y�c�+�M���R����g���g��/��u�~P�囦�2D�	=��,�4%x#��f�<�W�5�K�|�2�y�񨻅��s��!�_�f���A�`�/iPAN�^��ж���$B~��P�/o��L �B�b�m�&��q[kk�E�. �,y%z��U<Wy}�3d��eFKK�VQQ��	�����p���_^0��C:�W�V��߫��<�E �Й�}3)��?/ ���\ ��2m�֣p��D�U��aq%Ae���8����!e���A)nO��2÷~z�����������/�C�e�9ro���x;��t�ޞ�@�{���M�Y,��k��̹�*/J%l����D�����nT�Bui�Hӂ��|Ցp;&���KH% ����ew�SN�*����-(��!��K��Nu���.#c
p�uIII�	i���pDn;�&�Zl�i�71�NH�W�~���l HЍՓil�v))/��B�4���(�[JDK[\���m�oVf���3_��	8 �ն����7�.�$PR�����ϻu+���D�)�%�
�]�?6��;*�T�\��>��!@�CDn)-����@0����gW�^m*��,�#h)����p��❽3sD����Ÿ61+�|�/%�8�ŏ�E�QT�B�܎)� H�{co�-�%�����'r��3X�O���(77^� +��řC���g?��&�q��DW��g@��h�P9�)�-3v{�;�mZ��v{5튗�ci���UQe�D�7^ěj��ڝ���`V���Mgl�WDk��R�j�cuzL1,�+KO��j��}R��g��sZ���ۏ�22�#
5�!�w)� en(R��f��Гu�?��x{-~�?m,�v�l���b���p����ɪ�ʁ_��|�r|%���&�}b;����:X�ܮ��y'h�_�݉���yB�(�����񴰘G&6�+���,�!B`c$r��Q�W��Zʒ�y �bD���V��+?��͡������7),) Ȋ�*{	h?4��$���o�=+���޶!�o��8j��k�!��W���S�� �} ��[��m�����
kjfP����x�X�;��Yb;����I/@$���.^�i�A)��scN����̘9������"D�_���9���/�-�R�[��r]l +#rǵ�^5)�!�V�,_y	�L�������N��>��ծ����;�-h=�}�X�R��x�Xg@4Ʉ�N���X��!��*��M���DsCh�^�Kܜy�Z	r�$�4J����B�22vh�g����U�"Q;��X%��5��AU�e�9)�D�� ��k >�����z�F�N��u0��B;���� �ʄӕqT  ˣ�v�yg���"�Qɋ�:��ٔ�Q�E��c�hY3;�n~�F�^�<9��K��4��u��E+�5�5�u�����)p�d�M�)��׳�3��Aa��W���5���H=7������4�؝�O��>}*SUQI�D��a��iYY��tT⨶��g�H���jK"����f�0��P�ξl�΍k���y@d�|�ȉ�_���IM��=k�H�r,��	<:�<�,9{$"}S�����+-a�6���Y`�^���X���
k^0�x��#��0�1�����C
I�~,�l�%�
���n��	E��Ak��1Z� g�.�����PbČD�4%����G��NĮ}{�X�����y��%�E|N�l%�"�)���Tu��ح�|�O��bQ���Ot������������c�&��?$���[��XX�D �WOں������?� ���YS��3*+�EK��� *+1**�sx�$���&Q+��2�$�W���i�풱���ʽ�!���^�F)�����m�P��u��G�$�"#��+��(���BX�$��>�z�{� K�� ����	�BV�j��ت� x�2��#@Q�o����`e����xG�:�Y�Jeü��	է�#x[K�6�.�>S��X��m��$���E��%$�猱�����ߟY�C8���ХK9|F�j�@~˽�$,
;������l�M|W׿�.�������&�A}����زjϞ��2���p�a}i=	c��o�v��>�X�ϙ7I��Ą�QE�٩��k1���oD�w$�͵Khx�Oi?��ϟ�8yYY��;�x�}#3p}�J�tn}X�k�����п��HƺW�Q�_��%���)�������f:���)I���������r���LE�!Z){��p�X�_�r`)��4T4�������������K�u�@9�U�dm�(�`��i��4RY ��3ǛR~�ʙ�����ދ�p���x�;�)3��,�KU���@`#
��ƅ"��}a��^��˭_Q��3g΍�V����~UT�&̰�> �q&����7n���,o�Q�o�3p(ח��Z�c,�E�^��x�ňr b��m��>h��]	����0k �V����y.�?6���޵�n��૓����y������0�	r�.,�Z^^�.��������l�v��/�����	��e�a��v���(h�\%o��9ɧz�����(���tJYRkZ�1H��j������9 $JPe?pL�M�@�_@�\� ��6[;9���k
�D�Q���3snu�����%b#i��c|�q�G� f�N���sXfN[�~���B�� �JtV���|N��q�?9�xɥ�˨�p�v���'�@ǟ"��V����ʃ�1��· $H���k�5�U�s�>�l��Ǌ�8B�K�^z!%�!vV���BA�#h�^�i:���s��5Jr��_�e�X��!E�w�Ct��t���:��1]x'����8w�1>�:r
m�*��x��/�BK���KIl0M~��f���	+�x��g	��o�S����	cbtS�'_+�!��$^i#3fsH�;���j��b5J��Ή���"�C(|��fl��׏�:�DԠ�?>M����Ud�U�!>G�'3�x2,�� 2��!S������W��Y�X�V��X*�9!�)[p��ݡ�i�SB�YgB��8����WCͯ|��ٳ�V;��2�xGGo���ԑi���d��J?R�� ����2s�B/Y��s����y�JW�X�?x1'M�T!$�m� ߬A��O���y��R�f���ި!���z���Q�C*�i�A������'�S-}m}�"��B��=���<U��o�
���ȡ ��Y�F���h�x�3/4�g'�Xi)(SF+�F�K�ĩ��8����  �`���Ϗ=��%�{}�@~;-X��������
iT���2��]��cn.䭓��ݲ�-PMޢ Ʃb��Os�i��
C��|���\& (���6�*r�m�Q讁�:-���9id��"����w� ���X�7ۇ��كB�1%�J"�g��R��:	�yj�T�Yy �]��
��$��	5�9���J�1Cyk��;�y�o"�M��Ӵ�p�]d��9���O�рG�'I8�I�-��A�J�`2���ƣ���۱�L+�?��t������)۴�u?GE�q@r�¡0F�K��y0�"<ŭ �13�ʼ��k�Sf���p���b�#+q��r�� TZ�f�O��v� ���3sn��\�Y� �.����s���[PxӮc�\j���RԐxPN��Z�k 2uE�\��v�VE�vKu(6�z:��F'���L}�WD���l�Ӝ;Ϙ8�,��{���
�����o���ݪ Oh�u�^�n��O�'x��}NA�~ϤAM��7��� 8Ib8-{Թ�b��c�SE2"9	-�=p��
_
�/��4���-���E~�\�Y&xdV����"
Et9��^��Y�e�u*��6�Z�	������j�vN�0J���g=<F���kP��b;�LM2&F�C/�����	��6�D��{D$T�
:��#�i�s��Ȣ a[�wk-��?c[�#�5�+�!q0��������$����o��.2&����?\�z�汧��~�ƣ	��b�K�H!@%��$3�>&�X��fnȼ���IǍ���ޭ+�k'���S�ⱄЩv���HF!(J}�GǾV�ZM��>x�ђ��;��~�Qil��1,|�����`$�u�K򮙹�'��J�?∝�{$I킶m���`����#wza��~�}�&	�����W�q�S8�j�8�V��S=�y�vd�|�d�$2��̢�R]�cP(u��|����'�q�c��g\uYcӳ!��)����Og�+n�ZT�_v6�%M��Х��Qb�L�~E<�au��ߊU99�!95ɪ���a���8��m��V���E��S���� ���I�{�ә���8�>�$���E;h���a�OTYW�ObBMI�\&*��u ���f���\x*]�i�#ր�YV|^��-3�geI�&�?|���'�>�Ǌۮ-E-Cb,�;��]\\��&�S�r9q�[��Y=�:ۊ���Lԧ#g��d,�4X\	8qA�TTY������qMd޻Ȯ��
Z��dyRR��2d°�Ȅ_h?}����c��q¬��A�"g$^i6�
��K'��(��ޑ�)�����|,	�@��kwm)��nP`2233�P{;�ǣ/�C���uH��n���TUUec礈Z��2���yYء��$1?��YL����U����z�V�Dab:�^�#\¹4��be�m���R��@�]��(hF��JD[ʔҕ&�h�ÒQeC�);Q�$�����,�9uD�u�f̃:������� ���w�7oN[�0@l��������H��]sXy)��XZ'�𡶟.�����T��N����J�*��?{H�v8��^�N�"��=��h�>�F<~sk�ʂ-ʞ�/^���ʚ��W.�
~)�|Xgf?,�)���e�8� ��8<!��g��1��̊ �1
%�;�
�xC�U{4��?��Ђo�9�Og���C(NwJ��#Gޅ\dp+��/̜l�-Z ���J�6���a��d�� 3,,��1��5і���o���'�Cv�梠��?����$��Ц#x[���Y@ouT��_���\�R �מW�,ʘ�m�|�Q=�\ҿ�T��$/D���,�u�4��\g;��Q(��)�QjE�K��W���tf�%F���_e���us|�}x�����Xm����W��b��J򠏘�4Xx�ر�_Ѵl$������D�S���Ř�kʴ?,(�\G����i�F�㝌����L�<ʚ��k��dD�u_����Z�%d���c�Eր. �a������ أo�|\ǌ�b��G�Nt6���b����ֿ:ˌ�}��#|ׄ}�L���<ب���t�/� z�i�m�F���~0܈����z-w�\N����T�{ǧg?wN%�1���J-?Q�`�G�N���FK�����7b<�P�M�A������^��\�C객]���*�v &�_[#ʺ��z�����1q�ݻwU��ad�}�+�qX�}�I<EGIA�$u~��װ��&(U�	�<�H<��_�>����3/`	�>Iq���_����3��[3!8���C!�U��#]e	�	UR��U��nD~	q~)��
n{��N l_���u�9�(��x���K��wiM���o a����T�5�+��P��}��	V�-GIk�툫z> �P�z媉�/��%�!�-(�� 0t
�����GQ���O�+4�Ϫ�A�C�a~��몪*E4w���е CE���o�I��!4���:+�� 0�~��d��(c�9�&%ň�-��Z~��1���G�t��m׃��a7�N{8%�5��R*\%�?��+���@�}9�gb61c* �x�*/F�$Q]doŸ6���ǎ
+��̭��:��\��:���^�ԾȐ��U�g_8�
*��:2��AČˎ+I<*��Z�"'��/j�֏���B�2���(n�Zch�|�*��K�x���D�R��#��4M�d�#��kkʄ��b���_`h}cu�� )�߫����sEd1<�W���OAg��v#�Lau����q�?�@Kv���i�-���)��ege��[�U�`������6��<m� vSq��֋oUP$��lK�ϓf���V��Ȓ��#sss���A�[�7��#���/,�ӳ< {_4�������Eʭ1e0V7�[�)]�=�@��rUh�.�:�!�Vy�wK��D�g8����̜3+��-pe����`����� �A����QQFEM$%�`'��<��'���u�D��m�W��}�0�mѐ�����i�ԅ��`�%�W%u�̐~V|B�[f���I`��8��\�h�H�[�:L5=-Pd9 J�=�,���`pʥz8��[�>LV"BO;:NI;�����:!��,u$Z�-C��}���+%JXt� �y��2(��Q�є�h��B�R�1R��須��׮���}�ە���3ێ�I����3 ��� ��Գ�
��<Q:���kx�K�;s�LinhJ�[GJ<xp���쟌�0�a7�Xz 	=B�9�=�픒Č6u����Ð:R�����'"t��[M��
ނ �L��K4�"g�XsΙ�Z0��p�m%�R&)wլ�Os�5c�j�>R&w1.�F$P<��_[S�䟢��yk���>#����~=%7w_��O�ʡ�]y�>F"M���a�T^|�>��8�RH�~5/3++�ִ���uS�$��`��)��1�:�E���?2+l��Șx����3�܀�������bј9��()�߄1�9fD���v !�׹�	C^�n�;4��m��)�����n��t\��1>EdV�����P���=߇!{�G�������.'Ģ�W�t�s!S�Q
����cd{n=�Sy��Ր3��uT���`'����������D�y�_�CJߋ��?��P{�]�*�Py�L�t܅'��@}qR�����Z�i>�r��;c+�G���\2�$a#N�G	���`���9-�y,��/�1��v�'�e�*��
�h`�X)�����</+�����Q����>ϒ��l���g�����!?�n�٧V83� �'���W(~��Z�s�`d�u�A^�
���,>گ>B�Tr$�L+��~)<R�GYp۹AAA�(r��E�j`����?�T1��k��[�Mf�5�3����;��A��.)�ּgfК�P�Y����Ϡ�SYrvY�E��s-6vo���vx�絎6���T7>��^��Z��{&s<�c>��f>�y�PUEE��;��(��xVC��:RhU_P0A��������$⃨G������.�)#.B��:�Q^�l�
��c����9`	��cS�2?e�m*K"������`0�>�?��:��w Eb1f�*<Ƞ%�s*B͖�2�]�09�|���
l[�X�q��}�����^�z�F�t1<H&� i(:�������E��P�4�S����z�f��)N�{q閂�לɵ�.���*�;����J��Sr��0Q'�r�cA�bG VsQG���
����L�#�ŷ=H��2})zC(q��uf��J�ݘ�b���΁.k����J�6+G-�f�e�3y��1*����JD'���uFB�d:*@y����kP�5a���^�\�p:�]�o]�,��ɿH�o��6�#�\���S�6�X�.RS���d�w"1z,�V����k���h�1P� �\F�*k�w�ތ���NK���z�6FG���~,؂���QG;�Ӻ���T���@��Vw�@7����;�7��p�2v�=
���a��ۚ:��������ف�X���e0>���^�da,����u�9���� 7;k���J�x���t�,���sC�M�݃�s�z��ix�Q%rV�&uɹ�r+~�mì/̗<
Qހ�4����r��o� (�H�R�?��񣖆�F�jj��U8C��G�Mq��O��e	�M���G�|�/YL��ŀ�2�)]L�<��2��N�梓x�P����T�B
t%�3s�H��������7b���>p.����*�6�otLcYr�DR���~TT4���2dI->�@w]r�`��n�(Z�斖@�V���RKU�pwI��ӤqBB��ȞF����,<���u=���;K/&��F���~��.ߝ�ؤ���R�*L���8��nd�]���q�1��Τo3L:ۆ�cH9[�ܝ�ױ��"M��:��a�y��<�)yf�������
���3��⏓y����t5>m�6O��� �L�ݧ� `�_�K<Me�#��d��d{��"�����M�w�f����0�����M&*�K~$�[�VdPi�/�c�@�_dh� �2s�u$w�]�w
[g  �:i)���Q9bLGÔ�o��D��9�q��� k8n�x/j(��Gw�:���A���ۋ�,�\]�c�mD�t��o,lP���Tw��0��6���dצr]=]��5S����$Ui�n�w�P���_��H�SO��x���7�%�K�0�V�^�����׫V=_��ę��7�ތd��~%�����"��{|jq�Wl�����ĶA�#]�4�	���(��61M��'O������8�ba1>� ĺ�*t"��Y%A�4|C;�c6�t�����M0��]�!|��v�-xP!0G�eX�i�g�?q���i
}�Li������̪8O�e��A��X��g���Ǟ��F)lݪ����q2�^��l�)06j��r�J�y�s�o`T�1�׳��JSG� ��b��bv>�ϟ&�p5[o`a��L�JF�.l82!3q7J�),��*�}\����y�hzv�0�"!}��Ҡz8����ݷ�p,�KȜ &#c����&\H���0Nr0w���"=�VVw�8i�b@
�m�݉Y�q��X�m*��O�5��VW�o4�F�e��r �+���$=�����
��3��έ���ȥ�Nk9aSSS,3��	��f�Ns�86����Ү�����1�U=���'��rUC����BG{ߙwӓ��s�:�!���%��[�-W��2ʰleUUfUuu�/�@�����! u���܋��L� ���j�Z�P�`�Jy�����ׯ_'U�$�=x��^ۄ�ȟ��.��k��ڙ�;�;5�_JQ�ͳ�4%9��]ۗ����� ,Iwuuu�����(iP}�����"��p�s��eJɞ`$��
�d�bU�3����35��v-�ٲeKe�OY�]�么"���[����j/
��B��5��o"	}YM��A6�rK)BS�P�+s^Փ��S�E(�|��
gy/��g,`��o�1	;�/�a��O[#u:��D��<r{�;�^m+;��?�Ճ����/%�u���о�{G����(�eUT�l�ښq7�j�q�^В���8� ��j0�
�a�0�6�K2q�q8K�����K��)��>(HN�%A��v��)^b�B�[M��,TUPPؙw7�ϯ��cV�iu���4�>�~}�%�D����� ���f�{���>��'�0�:��)�:�25��G��w�.a7�}C(u'w��E�z� �,�z����e���|��G�)/Zt��0��X�>ۆ���W!5�
�$��l�?D�}�M�z��B����T��I���8�'*C�����z�Yb 
u���"c5����s��ˮ5޶\�ޙ�����jqpq��O���G|v��mk�LP�f� s�U �P���;d�0��ka� ��]0���?!?�[p/�ӧ0ȸz���aH(>��m���Ͽ�� �^��0��Uc69���	AE"|16o�Y���d��h���R�^����W] .Q�В�-� _��qP'�E׳(�nI�꧌��e�̲�D��@�B�f) *�b�����������O)�12��󇰨�d��2���T\-�J32��̙�cL8V��q���"C��F�*	����7��t��tC�tVf��M�|�"G�377w�-�G��5����� 8�E8݈(A���x�4i��vڡ��}#7G����Y6�����N`>r�ǎ��\��S�	v���~8���w�(ۅWm,_�N���
h �q�4�/��F���t/�3	e~����[!3"Qҡ�v$U?�i�ֹ���716��:�$�A>R��SC����Ū�5����W�ԙ-}T���o���|�����z[6#dk��O5���"����H��������sĤw�E��oC���I�;|�5̷��ѧ�ڳ��M��k��yI ����T@y���K�c3}}}��U�䩅�<�ga���Ls���Qg;+++��r��8_��pX�~=u�л�D��C�XX�w9bd����.A��F�ڰg����`�sc-Θ_--�6�:�e���^;������r,��>��y�����VB��y�LC}���x�eGG��1&��Rv��i�7���x��;����?�,�W*�FG�Y���l��y�
�1��;>�8zX�)��$�{7�L!%O�J�s�ςjbz��{	ƫ��)��d�oI;���,���N�5��BAp����\�+�:��:VB���D�,i߭�3�ԑ�gϞ]�:�Va�Sz�1$v�"_&B�kXs��I�|��h��=�`�Z�o(�VGO�z�q	�OKZ������o�������:9��,�%z�;���ob��3� �Cǲ]x�"��d�Zd���}(xE���:��ͣ��;J@�}�$S1����9s]z�z:3��A�7]i��Y�3;̉5I�X���tP���#�Ģ�I�MzP����W��R��AR�333����L��������x$�*�� ��^�Պ)�O�w��Y�����`!����^ŧA�姡��F~�+���M� �����?�c���CJ�W��h9@�7����������d�c��@x'���~��u@�E�M���ɫ�_Q�-��Um�4�!�Z����\�^���؍�r�@"���ȃE����[X���%2�z0��-�}d�8f㎸\ޠ�~�a�)Z�(��,|��07B�0��X�_��1�
`ǟ�J���;A�<M�>���;���=�+u�/l*��l���	۲B�<�������S_��	|���^?66vU�� dD~����Uw:H�w�?��b$7�4�[`t|�͝P���U�7o6�`l���=@�7��*�~#'�lG �Ӏ��VO^A�3��>$A��L v�sF���YFՐ;�O�ܡS�����ɨQ�üN����Q!�y����kZI���	�i��.�/�0�ȋֹy��8\�UQq�I9�:��:�
�b3C^�#�=v��E���mca�R���m�9���[��*����c��K��JKK31�g�������t͑g��H�> uX���<h)�ؐ��d�z��aB��7{7��M��A>C�xz���f���Qбj��hx�<�W�_dh��?Y�}R6��6�{ hh�W��, q[�㗜5�To�z�� t� ��M�	��Ѧt ����3�:RpP�����}=>L��N�- �{QR�9*K�����3J1���0VOޅbD{U76�8p`2v��B�7�N��?}��2u�:4�����ZvVm��V��oA6h�w<��uv�%�N�<ٶ�T��K^Nt�q����,%�+Թ�U��3�$W�%0����!{�@]�f J�R0v��*///'Ї��8���F���6$�=0:�+\ɞ��ѐg���A>��	7W�JK��h����	����L7X��3�L�g;�O7����q@+���wyV�ú�t��@,)>�������H�򧢼��uK���`a�ϧ?��D?؜�ρ]@̛�v������c!��Y�3�<�\f��.� ��o�# Cμ��dx�����㉊��U�j7�pQ3]�\� d��u��"�XvTvȹO��H�$a��!���ܺ�7��eCrT�"cc�5Z�*�"�$F7.����ʠI��,0i:�6"��������r��B���S �::�i5/Շ���6����(�D�T�U������ZdǇqCCC��	��_��?�w�)�{�Z�J~hʁV����6z۶kjhL?LuC�PZ��`�L���)�DUP���!# ��h�>��V�wf�`@󥺄�����:�a�\s)q��dBF~����X�R=LDpx�����L�����6���o�ԑ1o�Q���6��6��S|3�B�j�?(U��1���|�#G޽���DCf�mY�o1?T��4�Y�r���g��� ��Y
�����8h�����Ti�I�x�u�!�&�e�����.�V��a)}of�8 �΄�*'	ŗƌ�s�C�iK�J����r��!g�g����,~�Niu$�r�u٫���c��-� �y##CL����i}�DYHd2��v�� �^ja���9���\ZQ�Lڷ�i;4�<F�Г �q9�����0~�e�gj���A}.�ǙZ��V��ToW��� �O&߯�~׼�1����v-%?�tN�Bۉr��f����D;#L�(�#uO�K�'��i�6��)�K��<�8�cf�;2���-̱4�1�+HQ���n`�9�Ȅ)�oZ�} 7*�qG�s(��7��&)������GR$�����������O���>���w��r���6��i���u���JB��ώ$d��ǀ�����Ԁ����PRn�In?)*�E��	��p���=�x�5	�Av� ��/h]���c(U|X�aw�r�4�O�,+q�&�wy�S�s`N�&���e� �ƺΑJz2�y)L2)[��n�6@���*kj�O�4in��=Bv�-$���F	��� Y�8��Z4�n�m@5�̡�H+���	�ԓ����n�L�t��[�i)��e�ھ{�޳�����h��t�Q=�EG��U(�ZXx�5pT�-�����m۶堺�Y�<�u�݉5��!�Є+��O��A�E�]�'����X�x�aH����^ۏ�k�;5�jd�1r��w�Z�MO@CZȚ���P<љ�y���+��h�V��. �%�[�I�5�DQC�ײd��&���z�A#�	�K.�#���3Ϟ<y�vp�;I�R�q��,����D�[�y�:it�՞d�c�b�uf߃��(�򤚢��n�Tt�#u����b�����%r�
w_X���w�2r�F�ҫ8��5Eb����ڲ!3#������70�ؘ��{I�*h��Uy�ŸzrL1���yTsȣn��>��ֽ�Ej"^���p����vD�K��a�\gcB����YWt$�ğ2���gd�l<�,��jg>�?`$u�V��c��ܒ�V���,����9S����f����h`�`��Q���ͩ��)��<0�܂�Ў�=ʱ�Y�usW�^M�+]ۊpF6�nM:�ҍI&�Y�Y-���к���u�%�Gl� v?ǎ��-}�������D�mп�������)�$�g��>k�=M�ํm���dD�Ni{,���.�;@����x ��%�u� L��
��|>a���%���@=�Gy0���ݢ��]�ϸ�)������	4��!�-��8�ˌ	M�3<�Sr$�{�,YX�j�|�Jo���(��Ͽ��4JH�|���E]�<��8;�Kt'����e�WѯH�;;��$���|(Z �8���H���r���{,G��2D��tu�v�r��e��,u��� ��0ژ*��Sv�Pt���l�2sKصI�&�;��n����$ Ey�;3��|	J�1d�����&�o�]��(t��TQ/FO�n��f���_�
�ԙq�>r�l*3��B=�Dia�|{J�$�����Pj�BKآJX����=�J�}��CY�=�Z�ZE���3��뙙q��^Z'�<�ɚ����vm&W>��	�<ˡR�Pȿ�*����ɕt���݌���a�XǌIn�W+B������ఈ7|<��4R$�I����of� N�B��vV�B;*���&w�4��uf� ̿M����RR��0����u��=h-�C��C Æ�'K�T�BB��&�j"Nn�=�N�L���T������mu�֠q`�8k ��-���)�q���8mI��`f��r�г��������u^��[L/������F��RFF�u����9T<Wj����"D�>Y�d;�����S�2�y�S��KF�
�Hw$c�b*��Nh��2�r;��gz֡�ȃ��>ة���g[�h���@B�")�0MC�����zw+`���B�!ؐ�'%O��g�#ϑ���@'�s~�k�F�`,?O�l(`'��_�R���r��ݷ�E?Q/'}*M#��慰Z��{r�q�w��^��9�c��R0}��4 o�P�:Z$�y�1a -��1����+v@RdP����xĩ�,#�C���w?��82�w	�����n�d�|�����T��S�d$EB����y�f\�+��|a�^{��Q
'�{Ӭa�jZ8b�c���3{7$�]B� �Z��]/37��d�23�gg���1��sR�@t��T�5D;�u�dNJ�ϻ^5+����u�y���.,�L�"[� ��B�<Cܨ̾�Y]�<-D\6ɼzXX��km#:�ƍ���vn�>r/~ރ�Sd��Zm�x?�s�l3���d(�6(�Q:p,ی���e�/,!��l"ET�&���϶�
{�J1d8�oñ�d�\�9Z���q����$ _ħ��w��}�����U��"���W@�Ői�0L��!�Ts�t�^���PCN��ɑ�E��A^^ֽ{�W#�Tj�Ni�����-�Gӫ: �H*,�\,
�tm|Lʭ�����H�WF�A�n|C�l �	<sn�ؘ&�d(B�K��؝��fLu�K�f!BAkԩрtD��<�����f�+���r��nZ^��R�@�n�NLYN����ت�����>��h\X�����E\���?B�JI:/P����>%�K��9��ƪ&G跼�ϴ���.���g��7��n߼J�F��ʯ�j�?���U�%��/���~o�����ħm���V��vm����k���S��Ǎ�iI��S�n�3��������} ���/Z�(�ǧM~�+��B�/YQ[ŌQm��0��r�|���Eb酐����D��4|<:{�A���62O�N��n�rwj�\�cj�+>�KKP���;�y-G�'6�z�i�D!Z��X���=���K4R�A`|��GJ�OL��:khh�U���y)��H��ce���d 5��_��@�rI��� �Ϛ�t���D��O�}����&�.�I<� B���~�H�~wn?#����������bb�ҫպ�ۑ��a�(��z�� {���5��Y /���Gs�� ��!�ai�W����w�UD+�_?ņ_Q1N���"/�MV�x4����s8�v�A����2c���rs���3�Ô��wa%s���N� ~f1_;��������)�C���b7]xE�'�S�-����M?�Iou|���[��W����]r!P&�4��$-��n\�(�����~~�߭��jL>����k��j�Sz"���X�u�4���	ݯ ����W�:/@i4��d�PB��ĉ,S�6������r���s� Ȭ ,j�i*%���d���6?S}�i3/�Y�+�\�3H�<���c�^i��V�imZ�#��	y;���t|��c���,$���uw�H��;��s�u#�K��ў�h7}�W�wHZ�6����Z�(|`M	�<h�豈�F�>%;�^��/�?a�o�9�wEj� �&n�,��~�h���q��u᧟��s�U}m�R�V�-���H�0�{�u& g�nbjz��3����d����s�a����:��X����R��/���w���v80���9�)�Ȩe?nf�����H+��X�bV�l��$W��I��Ͻ��pY��=Ym���!�.�0j\�'��f�������p٪��U�5���^=gq������T�ﾁ�����+5&�R(���0�*T���@TΘ�p[�	�=G�/�8?��j���~�=͊>�kw]��M�u�L չ50gw�4�8���C�e��j��i�̘�ͳ��y#��,�ԇ�`>W�q�9q�R_���>ρ9u03��7���wã̘���VR�>��WYW�ԕ��CG��BS��B'Z�� A\�������Qv���T�%�*i�eu	j1�b�F�Pq�@A���(� ��u�	�>p��}��ܳ|�;��{�O�X�P?��t�I�a{�Q�~?c���;�ˊ)��ɍćtV;�.��f����^���:K�t�����B����~d~ӷ8WB����ΡdH`�]����P�+C���qYwMdz@djw|0��6t�իW��c��0���R��G��FP���oM��mf �EY��$�Ō�Kc��Ż���9���ݓ�b�?|�Q
�_��V�:PRb�pH�ڧ4���2G�}*��2����g�������V�4�[ ����T"�n��F�C�36C��� ����ս��k"��-L 3H@8�/�s'S�X�]�"!���_�	Y`�_MW�,���\<�F��cnl!��ʣ;k�GD!��s'�ȑ#.�`���� ��R�=^�`l��~��P=�}߄J4v�\��y�b�Z4��D��0`��o�gI���;gŻעmR�F�;��N����JJ��ΎY!�e8I��è�ą���w��G9�V��_�ݶ���Ũ+��]�e)v������V!�=�n(<�R�#��h}��Դ��䌞�wI���$;���L�:d�<i#Sa,VnaϺm�H��=�a��T{}#�(r~��oo�| ���0;�����k�M%H:R ����GB3��Z����8��Q[�X�W�mh��%1Ke���q����;�.<y�u+ڐ���o����=x�4����.�p)�R�xW�����C6p���uO>[�Z<k�c���#G?�o�o�D��;�*��c�I��_xR��sF"Y�v�4����{�>�! �-_i ���˪�B�4�R�5�M��k�e���Q6�.���0-G._~T4v~�W!���m	R:�)�r�n���������CXMҏ2O����G�pj��V�Z��b�]��`4-����?b��]���Dtj�P�<2]��U�-���;gb�Gr��(����W�n,B�bKr5&=�y6����I��#l]q����R��Z(���-z����	��� ��{��LUe�f`kB����O�)S�*�x?���R�NEW)���^�♼N���ܯN�v�Z���S�f��.b� �j�Z�܏��<�%���r��`ΰh��yUأ��eꖑ\( �u�]q�E�@�h�kj�9��41K>	�n���Ӎ�ƣ,)[�����^�_s�j��`'"@�Wmp�]��b�
(X6z�����՞]?�A�0S�`$|���Vnܛ��8$�I�S����\]�O:1���!�C�7U��/w�+	δX ��Kt��ء
��J}$��!���B��k�bF��q1�UEEE�h 3iN����JM�Ʌ/�2l0��r���FVW�k��L���Qq��l�n<�qCG �7ۡ��?-..��r�g^�u�Ɣ|:O��HP,^����~���P�>Z˛~��JQ(6��4����>�?���zo1��O[���t���$	V̉��e�a��i:�U�� RX��J���ܻ����5�*����pLB)D3k�i��ZV�ד�COq݄nU�Q��Z�x��m�i�,�Aޑl��.��[/�r+�j�|����p-k�y� "Bݑ�a``��V7�E�;(�<|����
�jl�@N �u�Z��@�u���`��s@�by�y@Kl�b��OԿ�ܶ��r��l��'�(+��O��GM�%���9���-j1����0�������Q��2{���Y��n���3� ��Q��.����yyZmc�tҫ��wbO-�A��"�kӚ
�9�+���&�����}��a}�@����4�zTep�fT�<��ď�w�ܳiS#�9lQ�p�|3�*��#7!�n���0�s4�4Å���y�T���qu!hߔ��Lk�}���ǅ�^UՙS(���^���|�x7��U��Wr��|A��(�B������ၞSvEy�ט��S�?���ux�!�-��GW�^$A<�&�Xxy��XKol�A��T��!rFh�y�k�:N���o.�@��1E�����Y0R��H52e��S� Ъ��xҟc�qM4���-L=�%AM^<d������������l�T�hg�i��'�H�	^j�{&�^@/do�܀ :�t�Pg��2 �6#�%�+�Z�s?gDa�����y~�F}���OA���� ~�ԠǷ��J�ہ��]8��k�������u�����+�1�Y��d�����'N�]�]�7։��!������G&L.��!ЬA�b7�s�^/�x��Q�,��"�pߛ8C,�e3����>��kf��FcT�ݾQ��Zz3j��b�z��jv�J�z�)��W%P/Z�*i�iq�
N I�C��k�����7
BS�R	Pc�j�ׅ��""��8e-0�� ���)� ���)�u��eHr�g	ԣ��z{>s��t��\���H�	O`��xbe[֘��x�k��N�x����*v-뽠��n$B4�=�[|��va����y�S7b�V�&98b��%��ɏԻAU�k��m����<�p�A��}&�L�8�[ox�>'���T�]�����V���Mn;R��q�����`(!,է�B7��i�h6d.���/���ؙ\�������*k�0�߄�Q����_�
���)��Ho������Z1���Pp}8�W�ye��Oڄ�2�t�@�Bڧ�rYf�ծ��a�G��B?�8���ě�eL����?��F��#A=�m�	�B"���)�"��=�,B;NXd0���S�m�GO�K�����,o�`Z��s�w��8ԖG￨�y�5R�&Hx�-ۮH559���>����xJ��e�Uea��+�Yꢏ��-�q��������w���=�Y	L�,Њ�4�wG�n�Κ��\5KJJ�I�!d�3�� ��0�{����< %�UC��ȫj$]5�L4h��:K�'��sR!���\�@��ڙ �
�����'v�d���:ko��a5/ca����!I��X6d ��Ȟ)ɼˋ������
Y=�44����/�d��u=����v$����.�j%*�f��%��1g���Bt!��!�UOzw�Z�V^��y���'�v+-t�W�9�[�qԞ�H��~>Ϻ|��KAJ�${}K�cW$?
vt7��a��t<J◑�����Ҕ�2�=�����iҸ���~u����&8�*���yT���N�D*ډ��L���;�F��	|5}�c�!�b�8���&CL���	o�~Pc߯*��/��`�PGn@��I-�ɂr�m�]Qs3R/�n�� ��qM�k>��ء�e���%I/�L�O��iX_[�GkP������K3��Ł�Z7A'nW�Go�ɼq�ShvuԠ���Ҳ�>͏
��e������Sw��� ��|����C*l{�I�FvN[���h<�2'�Qn��-���u-P�c�����]=4�	��T�'<X�Q5a�R��D,@D��t������=_pI6�����l�"q�t�g.(Y������$e���x���p� Z�ftҲ�k{�g(��}��U��gzk֭.�kۢX�0�5}���bh-���݅�����jz�^��|/�vز�|�o���Ƒ������ PK   ��!Y�Y`�1u � /   images/d9bcf815-618f-4ab0-b416-9f611d86ef67.png�i8�o�7�$ɖ�$T�ʞ�[�R��,ٗ�lc�Zʖ6�	!;�ױ�,Cv3։�0��`0�巙��x^<o���⾎�a溮�<����9�y�HK������+�RP�VQP�=u��/��;����)��;�4�N�r��;W��߱������*Fz [���3
0,����������.	'w����廏���Ɵ��?9=9�Z�dl�l��ăR�-��c�/-k/�3x�Vt�k�4K
�1�V����JE3cx��\��E�݉�	5�����*,�Ђ]c;N'�Ȟ3�=IZHͽ���	U�qW��&��{Fܸ`��9s�'��%��s��J:+S�����*�&�5��^�0��������UR^���S�a��-��8��"�������ˍ��D:g��m�>@&�fJ`{�S��3��p�G,K�J.�����_p�0^�VmMQ�	Su�5���@y����?t���%���Y{^>5��z��~�ʕ8�Z��G7��fL���w&
��#Ks�R`��NLF^��n\~�z��D����S��w�66�-V�}��.+-�ۡO=S����	���u��|}O�Wڽ����QE&����Y��'\mJ/z`NSG�Y~`hK��Dn�V����m���4�[L*U�@>��à=hÃ��QJ�:vt���Gu�ƦP��X!��^��?�/?���S��D�S�y�:����}�jӨ���(=��z�n���kEb��[�������+�c�ς�5�#�-�F���6"\��~���/�䕸�����A��tM�?h��㗙��1�Y�h�;�B+Ч����G�����sycė��?|Q�c �0�n���è����q{5A�dk�s	�d�6k���Jd��f}`��9�;~�U��o��.pʊ��Mf�b*�Vm��^��{}��o�X[�[a�4#�BVMn�N��j�����t����:5��Enզ��ۮ�v�|�x,�&�Nٴ�����\s�)�<���"e�_%m�'�_�sń�[�\��B�7>�5�iP]����[�n4�X�4����_�|t3|�ӌ���]��70<�����`P;z��� ��h���� ����W.+�#C��������-b�:����.�=����]���[ ���]��#�7�����"�-��;)3�$�"W�������������ݩ�A1׀���fϱ��`�������ݶ�����uA�t���(lvޕ�?}�X}\熧J� K��5�ͅ���ȅ1e��Ȏ�>f׹�X)�����ɯ�>�7������鬛�֟���(c�FՂ��7������j��y��FD�br�fk�֚���d�M�9#9l/�nޮ�w�R)��Ctׯ0�:�L�dÓ�ݒ4v~ɂCތRG�Se�t֭:>W�u���-����՞d�v=�����ˇ�i}t{�J�8a���"����M)?kC98!M�͞��Hr{|sPG�q��[|7R��>R5�n$_%��6j�d���lGh;�@�5�em�ܞF?<Z'0������ڙ,���Ai>����yk�	jD_ƨ}���)S�ڮ�'��n��)	�7?t�~)k�m�X?uQ6�%>�׊��&�a��7���
G
��X�]v���iHmzJ�æ�ΘJԽ(w�\�j"�!���w�L֮���J�F[��JdA.�P}�.YZ�#����!��f�bf5�&���8��/	�3�|'3���5�.Li.%�c��4�%)�MB�-7�]o�L�,$�����U�n[���\�_')A�Y�u��E,'Ayq��@����ieH3�,�]J���֥<�d�`�ۓ(�l�<����ڏXo�aCkBZGƠ����}���w%q����Wfj�<$��q0*l����>��)P?KL�P��l��D��dh����;��.����x��є����B��<�hU;b:�;�Hl�����{��r���o4��+�M!nߞ=_p��h������/߉N�ňe�Y{�y,^$KҳCfl�p��7��Y\��>��^WC��O�2F<q3��;�8k|���TT�8��[9�>�oǮ���1u ���U��P��I�8Q2��z�V�G�s��\v=ܯ�lZ��u���aJ7N��<�'sUaܪ��3=ܯM��d0߀�1��0���E����a���:ı<��&P�?�C�Y�kL�ߧ}ث����
��"d0gVE����$ ���e��JK0pAl�aT���)�0��'�w�ssR^�ڦ�R�[x�P?�g���4{{Z��Ը]�҃���Ny�7����� �>��1�v���ޒ�Ĳ}YQW���=�V��I��|;_|� �o(u�$u�!�7ӃH�쮄M~P8D�P���f9�0�zp�^@�meE��V�/�Y]C����7�Օ�v�@Q7H��_y�BI���
r7�z�'#�lyca�S�JO���a���:7��Z/�&
3��Ż_&��~`ۗ���'qH�z1熹��������������ш�ܦ�̞x6�( �F+`���~n�Ѐ&:5�����~��������?���d��8�'�#67�)�wՀ�ٙ(���,*&��fr����ï�B�K+�����O�{B,R+G%��	�ݒ+u;̱����]y��5��e<�^���Z����.j�	��&ߩgו4Q����ky4���|9��_���렉���DB�~�j Qѷ�%YT/8Q�57��w������S#n#n��x�O`K����d��`���(	����|��;��n��A7�"Y(��'"M3�]o�G"���剢��z�y� Q�}n&AB�R1Q�,�XC�����kz�=A��B'��r��n�t<؞/5�C��ỊWfv�!{��E����[#��0j5��6f����
�1
��x�l��P������MT��i��_~4��������\EE�ʐ.?fZ�g��}��d���2M�J���픷*͉�>{q�	v&N�V�|�=�? 	1��R`h�ح-I@9�Oa��^?��/��0K��<(^0�{޸B����@�d�$�Ô�V�U�۸
د��E���Xd���w�"2�`k�vq8�㩚e_K��A*��/��Ar�^.U��T��V�g&�{�7����#5���7�I��'�u=��GU�׎'a4��fVy�hǐbv�l�� �:1	3�}�j�x-u�&���#�Jw� 8W�S�#&��>��2��.c;5�/~��Cv��������+�?���(�\b����Ts�_�,��f���� ��bO�DK^E����Jk�oq`�7ト����N���2���k`�$����iO�2��YC��26�\( �����{�}���I=;�������6#��W�7H���]���E`l��sĎ]*5��J�u� ����Sԅ۸F�S���пG�K�t�m1���L	��u9�� ���}�̯GI�]�(�jS�Eh��F��n	$$�ѫ6t�Z������v���?k�3�q�)}�?3��M��_\�
�p�``�>� ��k��<��c�7�&3�ր�r�R���rby�^c}e7-),��N�=�jA�-�����q}�|l;�厞{�Onї�� �	���|&_DF���K�4S Vݦ�LM�	���ӚYT�a��@o�ަT��d���T:�������uA~�ׅ�8P�L	���R�,��`a[�ǅI̱�X7�=<z>UP���h�.6��`�q%H���?5�}��by��,����q(�P\�_O6�\|����e-��L�(_`�AG	 �~�!3�FBNmӾ}�mV@(NQ���"��`OZ)	^�D6�?6 �Ca�˖G��$#��
�	cG���!*
vhԱ��gS
f����ܝ�d	Q�3Қ $q^�׎���T�N1�; ����Od��`�ٯR7��=/��B ��ǐ���Z�l9~��:�?���!~RG�)���vЇ=Zb�� ��X�����li�@3����
E�Ʊ%̇U���QWxS��"�Jj2%#�8�{Q�w2h��vG 3�'�1�E�jF�LF��VL�H�hEj,eʭ?J8]3�Re� 4����s�?u���w���ѡ�H�Y��Gd
���� Ay����ڸ��������u�<��2JH�|x�u)1CB,(; ���J%��o_�.6�åC�y��Ņ��
�鯴�a�7� "��0@�� Y/&g#q��S\L��UX��pP�9�ѫU!��7Ӎ@~/�Hg���ux���j���N�2�\�4��բQ#k@��`�����y�a��p��:�"Ã�Jg|@^	?��������#�gs��$�#,�v!=N�j8�I�������_�}��w1���=������е{:��9`y9>�,�^-U!̹ �G�(�$�8�l?_������Αqʰ�q��ݶ@�ˑ�_[�L�����sB*n�����F{4猸o����B���G,Uw���ŘU=W�%o�x�7�n��s%=�׉�#V���8�\bV�}��6ׇ����XMV1@�9Xau	��-79�՗FI���m �hߎk�n��þh�o���-8�z���;�w�㱔��p>󃎯���vW�%f~��?�	�ƺ��H���)�-��o^��vDk�0T�S�M��}���y>��eT�R�jH`�|��+���K{ќUj��0y ]$D�8v��j4���n}�$��^W#"}�Q����S�$��6nw ���Wu���V���6���m2k[�>�m���+:��JM��l�����S�@��bH"[P	��M��J��rD���x4l4I��M�\3��k��\6��,~�q��x�G����V<)�~�c�[7�p�;_f	dkY�jjD�Ǿ��Tr��Ԇ�h�Cdk�����P��y��7o�橎\R�2��%&�]�r�Р�\%����9PW���T7��F���2γ��Q�9S�Lɀ����0�!��̓������^�e�r���P����:�� v��׃�)�۳H7/��zޜ�V=��&!�r���ɳR��yO����VzdA>G�$�ߠo[!�$�$��;c��7�-k�����,	1;6��V~��_H��Z4w6u@�}ni�o�'�@�vQ/G/�`M<WT۵Z[��M��d
r���z�5���sN2?k���R0�����x3�0F)��2���i���l��g���햓(�ɍ�L���կ}+3��[���H�Vf� A�%Bvg�o��P٣@-k#��o�T�Z�;�@�N�h����b�ќ��+z�N-&K��&�3RJж�����+Pu����-�������k#�EYdr���LR_��Q�>#����Qk{vOG�}�1p�t}�G:���DC�;�����aZ���'y?�P���!p�I�I5oP=�?��T����gf�N&����s��� ��%Ę,��0%�U����=��QБ����&2K/8r(�X���:m���^�i�AK�Ҟے�VD��Y�<ih��L����-����^�4�î�X&��z���`b�I�a���7�@u1YR_���Y����a`��*� D~1�S7)!�U��dsa�ƿ��z����7hR���ҐA���	���kK���ai/_��e9�x�Z��@.!���.�@ϯ���b�Ҡō����6Pv�p2���������vB��i�����HI�T��U��I��'s��/�rgj�|�3�s���e���`�ܑ�p�"��o]�zU�T$���7�J�h�V9�&5:��|�iʐE�pGpL2�5�!ʱQ�rpL��zf�Z�N_4��T��&Q��Ɏ	CX$��fT���%<\��Hno��:���@h�=JJ�D���.`]�W�]џ`�S�HDJ���è��:g��p�Sw!�b�Ib�H��
B�H�tx�.z-�6�CmM����>Z���}��Z�d8� w�Dŕ4<q�~8��^��|��w�ގ(!|��oi�����h��O ����ȿ�E�)0sO��U+!���`�Ы�#�z��^PWWg���n���RƴvRs�������S��>�z��`,�M��d�]#�C�5[����F�5VOX�J~=���t�t0X��h�/c <yVұ�率S�z5D���y��<<���Rt��3-~:��/����{�w��z��FAd�5��E�����^g��IJ�H�-��ۮRddJx,-_Ơ=�Y�p:w�M6���r��Xl,q��,�wѣz��.�4~#�	3\�E���^*�#;O�ST(�PC�r�F��T M�� �l�di�=S�á����y�e�X������%$�������{F=��(">[�q������+�			�uaM�:�7s����$;�a�����Q3�N���?��#������
�ǿ��e���i��_	���wx�J���3��ƿĭ��o�ꑊNWLc[��d۷��w/��[�A!];� v��}Iz�Cnw������w���=´d�Rr-`ӆ$*Q8�*�/�C�u��۶O��˰p3b�&!ƣ��}8:�L�I>�;!���C{]!���~[bPN��_%֔�_
�W�<[��$-j��.��4_����;I⟄�$��b���3@��Yt?�>c�2{�;��4��T(�_�4
�{(���#VEWi
���8������l�/d%T���Բd�տX�*�ǩ�/�wMt�\�$
j��s�v>�'
���9:'.}�9{�7z�NP����P���!�%�?Nl����4�V�G��_����k|KѤ��H"�p�[T/�F��&	<�8V���;J��uu�==@q|&IC�ֳ���������裸���P��?��?b��,���=[u�[�$ӿIX�ʳ�%�7%p�84rZ�cyi���g����̦��~���d�Mx��%���(8�����BJ`���� �Gw��ɨ] ��֜�!q�Rq�#Gl�%Fn�D��Ld�l��J������I���57rVY�t�t��AM�Jѓ*e�����:'ٮK��|c���Eຟ�6f��[T�LIم>���{Ù��ʑf{��L��٣�n���4�*������h�1&W[kg�j0���Ay�lz�EAU��WjްAM�#�=��<Z�j�]��Zs������_m��'�W�?_йa�g^��!�dj�S�g5��v��V��2�[����L(�j�8'*�ش
�	l3�	��ڕ�녵Q�I���g���!�S�Q���h�k'e_/�j����^s=�X��"og	��"L@V.�	]l��bU>�K����c�5?Q�X�e���9h��rt��8]��u?JW�]�9�����zE�e�_pή0*�nQZ�q5�^��&�����T@�eo�7�a*&��)�.�v�\���A7��[�FZἌ�����B�r�D]Z�Z���V���~8s_��6���7Q��	�\?C�s�'E�n�M~�1B��ؒ�_�V��2��E�~Q�?%ǅ������#Mڌ�Ka���0<!��/<GH���;Ұ�P��y鄤ǭ ��{������D�~U#�U����N��}�hAQ�6*
ݞ�
d��� |4��G#��n��hY3U{Y�B͐XG8�
g#�����l j�����#X�P�G*�H�V��eu����A��vO��0,%~\����r�L�������{1WU5�߱�M�,���N^�C-�:k�qmο���aJQ����r�
uo��q*�B�9���p�ψ����E�O	���A���4o���TW4��8Z`=�)Yv��An��J��á�漣mE�d7@n��s�/���u"�}�5G&�Z�,[�����/��Qv�y3vx�s�Kxm����1����ߣ�G=�������HM�D~K�1_�
�ҎxU&u?J2F3䩝B�>apw�u�E^nbV3?����l\�A�O����M�����d�~Mq�R=J�CZȑ��<�䍭�Ŏ���A�a.W��)�4����I�3�PS�4O�~��o��W�>�y��z�z0�OP�F'R?��h�>�:��j��I�|{���ds��JB�
�RX��}�Qڑ�|������a,�3��m��+�w����������"#,d�/&�����=�3���u��/LZ>D�1
L:4g��d]��hBx��m��h����nyjb�l_<+J8�o?2�F�h�����!qZ��08��v� ����q��/�������o;�55�}$i����^Z�b�ъ���[�Æݮ5����/N���)%s���N@��|˄L��:Iƪ�M'��
W�Ogv#���)�3zBw��@7���οpm����w�N�z5�Rچ����G��VT���:0���*�2�����c��/�8�::�4��e*���v��ێFÈ��2�[l�~Q���1�E:���ԌS���Y� Kg7>oܭ�g�q>�3rۖ�40��Ƌ�h�W]�1�{��j\4!�͸��~�H}�3�$���"�լ��W �A�\|�Y�<ٮ��� ��bÿ+���\ܐ���7Ӡ�X޸~+��`9d�-���w^T�y�cA¬��m�w��ܜ���_�cż��aT�/��$�"mB�j�=�	m9�یC�	��c(QC�5;�z�3H���A������y���[� B��SY�"#��c��)�Н&��ٷ�v	��j0���2�<l���ug�=AuMt�)f��{ϙ��^W���3��p{�r��ɸ_��7G���%���ϏiKtV�d9�
S���vy���]���D4*2N��JI&��[���?5c�����B�j�U�� ��넜E�O��B��r���^网И{MM�xS��u�'v�+$eΪZ��(R�v�z.!���<`����t|�W��Q�*��K�q����_�q3��<�V":6�2zuۧ����^�u���*��z���uJU<��'�v'��;~��
��������
�ͪ��Q#�2�#{�cJ��L�^�����"�����u^�����$���K�a1���iY�Sn�IR�[�������\Nw�l����S�p(��9r)t��j
�:p��o<�7GdS���l]���ud�S��G�c� ����ƃ�%b�Qp���?΂2ow'��p8���)y��� ��� ��s,-ȇ��l�@��[EvYΡ����[j�*{�␢~��t�q���m��q�S�v��n�T�1��׮o�" 5�Ef2Տ� �|�z�GF�q��e˻_�d^D�xPƮp�4e1�y	�W!1���o�g�v�ض�)>����r���{��x�.@��g�=+Q�8S�@��H��֕m_�߬U�I��|��*�G)����Vg��͏�R{w��]��q|ٍr��M���	K<�W�~B�	����p���Pq𰁊�ʫ���7�&��_�dZh���	^�)�T��o����1�S��-�N���Lo���4��ZZ?��}�C.Q������Ml�;F �lT�Q.��{�e�L6G��4P뢍{��'��rVk�~�g�u7F�7y�e���9��JZ�R;Lz9�1��wOe>6ջ�?�V5#ZM��w�jAG�����\K�@�����"�n�*���������'�t�o)�8y;(�??�Fm$�u������^�r�s#��U���ә�U������)e��Sg)��N�9z���A����]���S�]S�ِ�Kx���.3$9�`q0���5=�Ҵ܈^��ے�ǟFm�X�Y���8%����#m"�?p�b(��)�<��/��ɖ�FD���3�}��|X*N�%�Ѻ +��hQ���b��h�����!�Q���h���j*�N�,����%�+��{:O�)���4�T�"����FύSQ^,�-��S�mŅ�E�4N��&q,k}.�`F[�)����,���DnS�gE��U��t�a����)�g0\A2EC2:�0�Ы���9�{c�$�7pV�W�yZ��Y4[c�i	�}��YO�5��\��	���|�g]��[�ygy�I�aaH���2�З7Df������!L>w�W7ey�N�Y�u�k}s����5��׈������9S�K�����}GZ�i�T����Em�)�㳫���g�1��J�����3$�yTk����S�,d!4����2�J+�|��KW��6��V;��a ���P���&W�
���ǫf���#�!)M���0#' ���)��߆"���k �`�D ���`���mR�����	��������2c^����]�;��G���^���e�4(����C��m���XZHē�W�_|��;wQ�^�Ԁޘ��rԷF�3���[,��@�CBI�9��$���Z��Er�<��#�1a�ء�ຜ`#��xX#�e\a��˻�u��1�S`���3��b��C�/o�S�G�esY �&�$;դ��Q�{�;,��I������8Iėʋ`ռ��1���&+c"^��!}>F��N��=��X%hx���������!x�;?�[Yo���%.Z�휤�%���G�i�7�6�ؠk����rx��	��Sd�U�9=����RX-o#.��1hA��[�z���VS�(ٱG�aߪ"�~�p�*�U�����8y�9�
}P�҇6ұM��"��x���3��u�g��#m���Þ��
�d�a��6��g�\����f�{��*R�I���nl7�b}=*���c];`o�W��GF�Bc�toZa�PEeiڅ=�S�$Զ$C|e,^	��M-�iɃ��M<�V������Q�W�b���;Uz�e�Ӱ|�r���������t�*��r���5���&�{g��r����m3��Y� ����	v		�(�i�c�k�m�����e�T�$C��KQ�l>�.�l�Z v�M肇����eV(`�M������/��!�2ϔ�9b>2��T�n;�^Ξ�����X���z�c�6w:�ADH�<闟{�qI��A� *�Л���6U
?��M�L�) pʾ$�>�D��I!�1�_�ޖ�-�h�3�v��s��^�qǣ��M��G����,�X��$nW`��9Im�(�R�~���L���q�j�����m���=ыݥ�蠻���l���̛7V(�7��NB��Ch��s�3�= ��M� ��ۈqO�Fp�$,p}��ru�8��4K,S�q�:ka�	N�o��)��w��W�k���'c)�>��i�!ۭ�V=����<��f�}<f1�4���,����� ��sR��j�3[�<��`Eϊh�����XZd�!��Y%8o�z*�C�Cn� B,�G���cF��`N �6���l6����9dɊ��������� 1�ŀ
�EOZ0@L�B#�=@@��t���5 �P�pƯ|�N!ʲ��y,�OӠU���,�rK�R�E�25˯��Zze�HU4<jܭE�=��gX'�0.$����ܤ>�;{+X�ޝK��!M���T�LV]����B�����xȜX�a՛4w~e������&���m���ԋ���+���e5T��&�o<z�^����iG�^�H����<�U�Q���p���p"��cv��v/��YV�[�B *^-�tW]�Uy��5�vR�Y�H�V�@B�5��%�zN��Wt3`���RD�5��HD����.���[ ��M�l�#�n/���"H4)ؾ&��gC�M��6�k:L�M� _YU�4������l��Q������vے��\�������ӎw��A��+���n0Yq*���Is�l�&j*����w��$��O�:�6����ɪ˽"z7o�U�4�aO�?��>{S����r�#%�[Eme���%.C,��`2�G=�W��D����(I�([�Z`L��2g�@d�|��v5��ث{�2=C,ף�ԆGW�Foz�s 9M��HsT����Ve��`�i7�D�#6}�~��~vRy|"��5 ꠦZ�K{��3Bt�%L��3�5n&����"��?۩��1↋s������Iޏ.W�X�< {3d�#�ﳠZ�k2��AF��Tmp��6)hqa�v�vT��X��abi:���ߣrn����R�@б�^G���tV��a��Y)m�:����H��Io;X��:�x���q��N��8�P�p6}��w�+i�O޺[^�ѓ��>�.�~��j�rNt�t2�L�����ߥ�z���n��c��H(�(�W=DrhUiR
}V���ػ�?4�sr��͗�,D|4���3�Z��Զz��z����M�2uӲL%{Yd�:���k�,V�86T�����=cצ�X�/M��+������!5�XW�s yIt�w5f����ޤ#�f��m�B?��d[�������~ztm��Hj!��)���`]e׎�����]�6s;��[o=�+�ACM5�[��+R{�P�d.UL�3}-�V� �+���5%�� c���̆Ӗ��[ �!n�7J$&35�������L�ޏ��	hҊ����<
\壢f����q��'�NJ�#��e�Nk��!n�O��.#:��-��~�iO�0�j>rw�
�M.�.#v��l�����¢��h�85���%�!bR�{|3���ڡ;i�I_�UGO�C���� ����-�j�a"�G�Ku#P?c*����P�G���5�~���1~*���uP���q�x�P�2��N���{��-��\uq��#�헱�~sQp��<��* � f+���#�\��Pi���-pX}������=c;	!E���-��ћ,�C�#��#n�gD��S��c�Y��ԯ��V}���GH}����p�����>�?�t��ҦgY����U�H]�ˆ[~V�B�_c�t�ռ��K��if�N+;l�e�����齢�����AH�$!B�gȭ&v֣�K��#wkX;I���H�]����<4��[8�>݃{�P����v��+�as�g/2��O0����y��&��m+6��f�y���Ue������iy?��MX��RN�\#k%^dۡc���ٚ���{�u��t��:�b4^��
�/m?��S"�E�RQ�%��"{NH,�f����~�u������s�������&����j$�)]�D��(��W��6 A��%�%*!'h�0m��GWI��i:g;��ݐ�Ac�"��2����J:�u"�"����-���4�/����Ռ� ��x5s�D�{��N�E'��6�O������k~��F��k4�0mYXZ�A�N�5u�v��-+/@�I�8f��4�j9�[d�^׳Q��.�G�,y��8
;2����#���C���C`��<�h�\���q2��G�o��aZ���״��,�1����-�V8�&�W�\}����*f� �qDL��8�{ԛ&�<> ��0�#��%F�d� u/��AN�7R�WA	=��svħ���O'c��[����cX(�{�gh:Ԝ~�ǹ�0=�z��?�ּ��pF�bM��*�_�Y*����t-�0�(J�G�4���(c�QI��G1\�\����}q1���#t��X�σ�N�;`_��9)�ꓰcOla q��D<����L�(��$��.�Sb�����4 )�����i>�k?JV7�\�|�&�+�0��/�F�k�}~ͤ���F����H�Dg�m�"�����
�a=��K�����S���v��������5d[ڕ��Uiϭ1nT^NV)�t�c=��K� VXm��=���cȂ����e��x������hE[�q��9�t�5Σz������Z�ߒ?�rp0���������QΆi�,8(�2�9�\R�_�*,�x�i(ԝm٭��On�eo��j\�S�u�)����󺌾��k��s�h�~MZ���4��C�;s��N�Gԯ�ҏD��T�$ܻPƛ.��8��4i��I����o��nq�l2QG��F+�b�u��O��-1��6u��Ptv+l8��P�Hs��}�J���H��)�BφԳf؄n�L'�����ޫRp�V�].�Z���4��G��Dߏ����hs�=�ͽ$�%�-.0�������{�1k�S]����#s*1��֘��GBG)�,���_���9�0��ʠv�q/7g�[��,�@e~)�𙓾zT�f$�\�V�ǌI�-�k�E	�X��X��� �iC���c�lSB[���)E|<~��"�B��@)@k[8��p��KO�I���cƗ�J���m�~O�tq��W`�ײ��2/Z�؄��^!��.<�dm�1��\�Q�G���Lok98���M* +k�E�� Z�[
��dԴ;���;*�H�T.aʲ�4�::԰(Y+c��8���$	U{�U�����FH�4��gjTֹ��>���M��y+�U�֋;�e^�����y�Eq�$�sfrv���������A�6=CL6�;�+�y/Y|$�Cok�t"\i-�1>o.?=�`>G�G�)�q�-��z�sC�m߇��~�;�G �c4EP\�un�薧L��$��*C�3x��K�c�K�CP�߳�^�'۪��[��Z���|��k����N�E����XPHSmڨY�A��s�&j����~睉]�*���Bf[�e��w�nG�[��i��5Y�K��p�r�}��'�H�P������G���O��qx>=	?m�eX��z���a����57�`�=��7�R�	�q'̟����49�*Q8�q�Jw���&~�4y�(3S�C��+z #�e9NО^jQ;:L��	7T�m��̡i����D>J�d��L�o�ߩ������`ϕg�Y5a�6z�G��DWۧr�	z�:�R�-G5��E/!���ٞ-Ê��l'�m+��,��Z����L�T&�c6��[r��K��C����c0����6�Ǻ�.���.p�f�p^>^�X'a���L �L�5~m�ԋ�V@6�O6�xwZ�e؎�͇����>?�>��*�@���*H��0l��-�B�B"�o�7����cA���jk����/��v��7��*���w,�l�A�Pa�A�ϓ�!���I�� �������%j�{����j��`xLsj7��d�gA��|�t�\,��t�}��N'�[AhH�X�N� �X�6Sx��)��О���^�6�š�H��œQ�`�%i�"l^]A���������wj�l~ւ|�����I����ߊ^[{��I��l%j�b�W��K��7��!���!��d"�?� �?����o?�L��&��:wZŗ��{v�s\̨�N&q�@;�t��M"�ӵj���_���|G`d^jWVq voT������<���.��p������;SdԱ�T�^�Q�h�*x*Y^� �͉�5�b���	��������%fs#��l(SO=�3=�D}ϗ�n�o�����qc�g2��e�M�.�[~�
�_���RV��~�ih�2b�����m?��>��}4	�~��w�D��Tz<�H�uP�O��� 
��8T��k�pix&}���J�rK%�>F{~��H�_C��X}��-S���W(�x��Ąn��W:Q﫾�+M�����`OU���k+�rߞR����^�2"y�,����j��G:Ѓ6^���.u���r���x�ڢ,
�����2gw%֡���I�`!��RX����l�y���9-��̎��-�8
4[�K��	E��n�a�U�+O$=�Ͻ!K�'JS�]����<�b�A�nq��ې�C-��d���ġ'c�/5���ŏ��#Ó���S����m<�m�B	�FT`��۞:�"`W��$���߁zS�W=�f��F%̲�;����6|.�砛��.�]%
I�l� 5��d,�}pK4}٩�]�3��s*m"��ؠ���ۈ6��	d�������_Go��˜=y۵!�Nue\�*�!�2_#i���S���W����1F  ɣ#�ج��e���� !���G��� ��Z6Ѯ�>���*�<�r�' ~K*҉Aq�i]�X<��>*uO�
������ӏ�׵޷p'2�d�`\ev�d����l�nk*��2���0�$��M~1��1�U��?D�ΛZ�zKa��)9�\�R��>�6J:J�Q}ݻ�{W�ߟ}��E�D�9���2���v��d���FAU�U����b�j��ڸx�|d����Qq��.�%�*�N	{�Bl$p�\ש:�v'-i��U�y9�B���"�:>8}jp�����< i�#O�Z�5��u�5��STsBOk�/ii�V��~(��*�.~
���ڵ���'�E��K�f� ����Լ��A�(�X�L2��UE�"�<bam�Zv܋ӳ(�'j���M~ԕ�7K�a���`����cOa���W�rs-�-h��L���rAo9��*��i/��m��������Ο��*�`4��B�9!C�PH�%�7���_pY��/x�$�J��\ot~���_�2�ypR�UL�شnޛ7өV�a��<�ٰƎ�w[gec� �Y-����N�t��M���[�/m-f)EmN^��J���~��"ǁD���qi�ril��$yZ�9�~�؝,�/?X�U��♳6SI����;и�����G9�|/���w�DA�)Აj�F��K�K���u(��蓠S����������rY,nv�����ΐ{
�R������3da�Ud�$$�ҝ�r�ժn`K��bc�mv*���ߊ�Ka�eiS���N���k�17��
�W�R��s3�؟N)͏���/���|��Y�p�2[L��lJ]�i�e�p��R=���B�s��^B_i�٤��N������{���'2�m�|̔}n���TK��|��!�^]Y�#� 92�wS��Mfm�=b�o��沸0�M� ���l{���͜$c�茁h\�)���d��f+�ـ�W���'9�R��R�2�0�m�o�=u�H� `I��E��R�v �c�bn��L�l�W{���(Ȁ���~�)��9J+a���@p���R��y��O'����	c:�~��Ol�a)5="䍿h�W�����l���غ갨��� ��J�tw���
H))-�]K.-!",�)��ݱ��tw�K/��<��������3sf�=3��s��D!�m���O�ZW7���E�*�}�;m�т4������.�,�S�F�m/[�P��YmM��\j��yxrZ����5�m4��7E~Z��v�-�92���}uO�k~�)B�O}%�^���^��{��!x�9189��Z$��Z"�{��R��<D�^X�]%@.�=4�Z;��,Q�Z�D�'�ĕ����Dx
�D���p�ʹ�q;��'�a�1ۍ�ӕ�'�[��y�bY��*H��%<	�Z.=��$ΐ/{�ɯ��ܘ���𑆫wC�DO�$�弣o���FK`ȴ=3{�G��킽�^՗�^:������ݙ;T�6��mϷ�tR�E4�/�^;�=�:,^7w��O_�W�5;�����[��T,�T���HLT�Υ?��-~J6����[AL�r��:-�+�zN�
�%G�Y�f����� ?p��Xdc�P��~�a���\�-��ܓMT�M�o���G>6K������%`�;��{��;�P�U�������l�y6Nܜ-���W?E!Y�j�6t�M��ƍ�1��� *J��
^�c�*^���??���PV��,{y��7���;qu�(6�.�@Q9���g�<d�׻G&Z̋�1Fev7����y������b�9-c.��Xya�y;;����̯oiֶ���r<{H�{r�	�Nf�)j��\L�[ �L'�#ƌ�@��g_V� �r-fl-9/�LU��	b!�`qq�K�~��Jdk�h�V��~cc�e���Ԣ�k_!�����Łg���֧a$�l�[��۞�0b-�l���F�e�s����b��蕚�G�u��z~�Y&䵈6ŏ��eXb"�a�Z?��&�RS�.�̞��ü	'm����݅@p�l��V�ڒ����~��5�p8�y�O��)��o�4;P�N�r�%��=�:�Ĩ�Mk-����о&S��2�l���@RzX��Ր�J$����k���ރ��Y�}ө[0%��iO|z�;�N$��E3=&�U��4)ꭏ��&WWZW��n��[�����K�..�;9l���AΔ(�~o���E�_���QCTc�����`X^���z~i��
�(ew��p=��^ȶx<��C�^w���]���Z�5_���ߋ�]�ὒ�~�����ݸi���q���>����W��r|*�t��c�nލ�kQә�HilJv�e�6��`h`W��N8� �V8K������s�j`����@�����@�tK'�.J��Ծ'/(�\�<�w��iyb�#wrΝ���ij��WV{3���)]7~�Mo�:�N�M"_�@��݀ы��۫�d���i6��Tf�Ļ�P�m�&��mE�ĭV���8�i����H11��$����ҋA�Z����gv��g���W�ơ�({��G����ͧt��(�Z���X��X��#5n/GK�����%��غ���掮�CG�[X=(��?[�KNW'E����x��y���.���Ɠ�,t�z~�\�8�+&ى������g��pG^��7&7����J�q���oO�zؠ�]_�V�c��B�$��0n�ٸ9&\y��>����<�4P��؛{�^ �z[��pa��xYz������V00O����/Hd��@t�n)���@A�:}�k�2uq5{��?Ax{M��s�>����floB����^]W�nu]E��&���JS���`��M@b��5^�|�<���g�����2�`x�bS��X8�3��B �3�q���F�U/+�D���.E�9ԍg(��q��
�8�6g���`H���V{]�9�p�j��� ��*P6�:=>2�५)j��4�̓�Y>�7�H��4$p��e���������e]܅M��M�@�T��˦��ů��E�<Ay.�	����W�+K�}�d�<Uz���K�G��n�T�BS:�V�z��fH�n��#��ܐ����=*4����[_{v|}�u���kQ��h{߽�F֥��Y�:ps|Q�^����LP�_Z�6���O�D`�{��Ⱥ����Vh����l�D����J�.<rW�g��ڇ��\#��Yw�b�A�����Z��1Z�l�g��S*��YBkj�wI�|����T���jٶ���^��͜ΰ�u��ċEG�#��$-9��ܫ�����.����o�`}I�[�ZoA��ו���T�x�s=���S������96�D������/%�����6~�6f�خ�_̻*AZ�V)��J�zy3p��%gYX^��mf�����O4,�}3�i�!�yq� �ڍ�P½uN��0,0���"٧�{`��AR]�Y�]�O���
O\�H�y��A�����Bh
���8Y�^����`��S����B�׾��`̀J�D�M��#Ђ<F��ނy^����s����.Qffo�ԍg
���\ΐ�R�������P�)���D���)X;6g��k<��� ��d���eer/o�7ٕ��t�������%�d�Igy��������i�(+�XLκ��1����ucq�2;�xC�Ş천��8q������/�+�?�u��uYvv��λu�OO5�n,�컻0�s����ܔD�^� �"�.Y��I�bt�E�����/Pw�ش�`�;UHD���݄j�� ����t�S�v���-}_v�ؚ9Pt�S��f���e_T=��&�2��I��4wUD�0/�E�j�\�z�0�ۛC���|â��_}�q��ƛ���b����Ƨ�=���F��5�=8���<M�����j����y�	M��Pu�������0��:��D׭)���-#xBA�/���Y�#����\�1�I�A����q�������c*!r9ֈ�-���t+ʍ83�m�̈́�:AJ_r�M���k��oOҔ�'��L��V3Wה=}1zs�A�V/%NzCm��gka���<��A�w� ��ᴹXН����aS���x�������ݶ��YuZl�V`3����=#*|d���p��_N^!~j�{��Ԕ{��|ih�K��c*Z<\�q����-N���Z���@�p���(�xiq���o�@T	`�%��x$*�|�B��J��v�":l':B��U+X~�(���:'����͕���>�,�^����X�MK��`�'{�X��(0\��s��v8�ڒ�8�}h��昼8˱[Y�}lP�=��	$bz
5Y�N8S�6�d��k�_����f��j�s>��U�p���ɰ>Z���E�o��ދ��d}[�-�[�Ѽ���@�'����9v���/�@ݏ^x��A`xj-� U��[��h�*P��^�� �aBV�-P�Խh�֠��Jrz�	U~CU���섁��G�	ۅ ��=0is�_�[22�E��'�}�@�µn�lh�X��Ȳ�*���[h	��Юx~���&�o�$U�;�}�WN���L���{X���E��C{0���،1m
z���d$�%��=�U�%f�E����#��j_�<���5r򥥔[7�K��IOe(QWU��%���?�nk��V�}��;$E���r|�?���~��r�|��z�e<��D��AIh�-CA��xp�*��"��NWC�u�7�*��<�	�v�8'��D��	�=i/��{L^gsS���.k�'[��L���x�&�ʉ��U�?��X����g��]�r\�tx����c6�xOuCp���@��3}m��m���� D�ۡܻ��P>���&�X��;̺�^���x�����ȇ9����S�$K�]ag����u�Ea���q"��JcD��#�/>���s���!���!�f�ê�K�\��9΀�ڄ~�vr�܌o�`���u�S�	r���_G��Ԟ�gN`#K{L�Z����^y��|}�I�j�}
81U��.�:[��%����2o�t2E_�r�?f��{ZN?�;�B��}A�޴����Y�?��e��/�i0S�'��݈��O9�ܵ��%4H���|������+���o'"J�6���L�����>�����gJ��r���	�	l�����P?�,��:q�>�ae�ϧ�b�Q�:0�5Ȯ{�p����|��DS��܃zFfXZ��D}��HQV��V"ӣ��7�̧���\L	��mkO�b%\�*|�T�cp`ꨄCd��额���YH��f�c]��'��iE�D@~�y:a�?�����滼�f[m���U9��'y��t�|Vl���G��a����O�?����F�|�>O���&�9��W
UV?+�l�_��:V7��^����hN��v��
��/CE�:8J��qUw���8o�~�z����"+1�w+��pKz���_���7FC��#�����	^N�ӐNN��B��!��j�|�V�o�?��GuNb�<eg�b�X��4D���A@@�C:��4b]ޫ췇2������헚��s�����TCm��Yr`|�B��؍��kT�I�@}2�=��o>�8�d���Ha�]� �;y����S�;�,t�� R����^��o<����g�G�Q�6��,>,��V�'4�y�B��h�M�r���
�C��Cx?&+u�A(le����^��FJ�viН]3���A�8�h�0�T=�p��X@���K0.@��H7_�*?��?����s�g�U�68i�����a.�y�� M9��L��@���F�&�!���~��[�b���/�O�HZ��>�po�s�a�1����w��=�B�'Ц֣���]��q�E��Qq��:�u'����/�C���6�������ޠ�/��YNn�xgǷ�!�j�	�ѳ
���/4R%�?�'��nn�JGg��<�h`+�Ɨ�߅���}�����KF�']qm�1-ܗ��7t>L!���.|p$g�����L�(�a�4�騥E������~z��$W_���w�nY�켹u�����Y<BR�����l��:���˥/�p=��F?�X�B���}�j�wJ5�w���f�:;�.�3��0O��,��	Z��]�ɠ���u�V%��_�s��X=�		�9 j �/��5*⹍lV�L���5�TX/���3B���l!x��t-.E~���ܒ�	4G�q�6��*@;
q�Z4M�?��jy��߉ rs�b|rD�]��`�guM�GUhX�C��Aa: ��1�_�J��k��W�J�8�k8&�'EQmۣ�	;����V�S�F���/�(�[2��o6��ԋx�2��C<��b������i��lÿ�>ӓ	t��D�7��^$$��^�m'�������g;8Ʉv!�Τ�b9�Q����V��γ���7��ez�$a�8ߗ�2��dj��w,Ӳ��l�]��Yu���c�*���'�Aٞ����ੌ�(���z'*@�N�hu��teZ�>k��hjɪE6��@�]��dĬ��������8��@-�U]��e�0��V�1ѧKo�)�Q=����d�,2���l2�@]���

�߯,�91�������2� 6�lg�:��gPږ��v���e�>_���m��o˭��0�G��N}�s�F����������a����W�LUq�~���4�������>Y���A�m�����ζ���Bw�;Ӯ�@��dm��������c�r�[�ӮIU�A#�=�*O7�cΣ�Ku���+���c�7�<�{�(M��.��7ݷ�_q�^��a}{�<ʓ�n�˰���i������K�*wD��Ϲ'�9�~�lLw��&z�Z�D]��o?F�)谄�"N�������G4_3�@P��>P-@6Rj]���S��EͲr��NK�2te�n oQ�\��%н��ʩiyPJ�����FSs���*�t�owI��&i2L@W�b�X����4��jz`�4���Xj��rҾ��r�hx�1A#򰼡<�.U%M-�O�L���6o����pѐ��M7���\�|�;
�n�C�^(S�RN��`�P��y��Ki��4j^f#A��_O�.;U, �͂��Z�p#<8:b|���
�Aw�ݸ)���G�QF�6��x������ #����P#��Ȓ��R���Z����r�Z�;�1�b
.�����_]�O���j'�JY�W6��|4���q1�ò�
��"ɡ�_|AXXw5U�9����{��)�-��(8�K��9(5�H�	f����d�-c0��\���R7��1��k��*�P��)^��󛾰Ǥ2͔,`_�C� T�f�^ x[m��k+��4��eΤ���Pͻ!��@/@-�]�9*�4C0z�us�A��>���h�40�=�g̴3��2hP���=-n����]J�C���2��͵�.�~��l+3X<����j�2Y������C_e*4K8�WGʹƤG��r_���+�$�	
+O;	��:k�we��	B=�{�(�^��`!ĩ6�D)��[�Hq��lx_�?��.���M�6�28>;�4Ң�ұ�5W�����?R�?��c����p�,�7��G�g������5����u:�z��b �T{%*f��X��9>�X!g�"�@E�B�K����Ҫq-F%���1�L^@<�lz>y>�s����xL��,)�Wڼ֧]�;+v���K�����U�CU��R+�����d<�x�H��w��w�����V��m��kmqS������=��x͂$ˋ7;�ʲ���i��K����:��G�]���T3�l�b�">,u��ǥ!fM��E��(X�itIq��. ��N���C��DΖ�z�X���U�*%��0�M��ۘV�|r�z��a{sԉ�\������n���b���C�����af��3�:�� �^��+2ĚO)""���7<�(���>�+%$%:;�[God�oS���ؗ�%�q��!�sԣ�U3V\��1���\�0��A���1V�4b�*���>O*��ׇcv��ZOE.���ɡ�\���K�mk0�q��s��l�M}��T�߈��Y_�+P����ͭ�+0�8|�CV	ׇ\7dԷW\,��C��^8�ɩ��I
��ݙ�c��\�1��9���)ݢ�*Vđȶ��0ry���w��jN?R>��#)D;��;sXP�I�̈́��?���V@���K�[L�b��Yj��@��:)ȿ
�K� �M�O���~[���榊��g���=a�;�.��wP���}/��@��9E��g]��A��S]?�͑�O_��Ƿ���u�̷~�1�y�h�b~���M}��<�5�$zə[ȯ1�k ���V��>l:�&�nS�8Z.?Zߠ��ku_t�i�L��ۓ�ڠ�ߧ?;y�L��5�`������s#8/�p>q8Tq�J�q_�k�;�>�^�A�{�{k+����Z4y���|�S>��pnLf��i�,�������1� �����o7��*�+yP��!���,K�M�v�4�N�sL���vo�5�و��Η���D���Z^�G�ܽ�:�j���ȱ��t!����~�(=!9;�ߧn3W�!^1+���L���6�0Bح�,������@f� `Ӕ���?1	��K+�!����WRݢE�m{�����^���o�cD3Dh�֎�Gz�����~����P�9�1�j�z:U&1[)h]=�b��H�������!��A�If��4��8E�1U��P���V�J'��?�f��+�%���~���<���fV��s�0�C]5��a��A@q����:O��~�*��H2�R��C�\f1T�>�x`H"�9�qQ7O�j�j��K���yz\l��f��B�����8���~v�TMmB��u����͔f��;�:��Y����N|>�)f�ZJ�_���vx���35;�*+p���'\W��j�����-ؖ�L��b�z���p�$��C|@)�+kq�
�L��Jη)�i���I1�o�E<����8�q����xڜfc#d�ߵ��#,�h��k��R#�L'7����<��7���$���c����FQ�����u�3X�@��ό���*u{%��a0?r����	K��
��b�w$w�X��x\���I�$�)����������Ι�3>��g!�2fs�������(��	Mg�;P�_@�V�ܯ�d�_d�L*��ڹ��|U�o���{��b�P����虹e�����q����~Ɩ�@#&��Ѣ�e���_�;��"��ݓeޡ��Y�x��r6@k��r+؃���ˆ�J!�
R�0��ϓ���oi���G8��7��	�N�7�1�0:�q����w�̉J���|m� @|�_,P�ϗ���B��������`����3m-�4j��j��R���ȓY>���c#F��ȴNYl�Q��$��WV)ǣ�Z�_�B{z�̭���'	��9�h&�4x���.����@��i.��B�3�(u�h6��Sʿ�������@qW,nBy��E�����; ��{����V����3[d/rЧtzc0�,%�k���e���:祾����I�#���P��zr'��3����rX!,�+e��hEw�д��������1�׃��z�K���U��Y@,b�Sr������u�YHA����Qc�dF?1�[������q��hJ�^B6�q�X'�屛��E�rm���{8E눯�����'$c�0A��h��y�7z���P*�k�'��!
���XW	<5j�!'t�t=�i�9�Kv�F%b~s��/|#ھ��a��߲�tU���j+jX*�df���?��)t���)� (�Ťdw�,.���Yz�w��?��_Gp��߯Ь�-�a8����%���X�Uǡ��lz'�3������f\U!V�7a��,qIհq)؜���\��1��r(|�4�x��o��p:������ٚ7�}��������{��x�+��QsD6�L�iZUk��FH+��QW�#��;AU����Æ��������)�`��  2��?.���X�+�����\%Y�@���$I���Z����-�,^Xt��e̿�tg �d�g��>7J�)���c�᎕;% �lA랝�j���n��d飷f��t�^h5�f�a&.�0W*��d�el'��Z�dW�-�靽h��Y!����j8J�Q����Lf�`u��jz�9���ͧ��lt�ɤ�@�ӥ��4��PS���2�oy���J�b�����]����V2~wۨ.�N��Tewh�+�2�d��W��5�q�7�Ȉ���]�K�,:��o��/�G�Rί����q�ϯ�=�z�U�2>�z��;�wo��1�(�`�{/�rG2�;WAcB�>�;W�Jq:cG�&W5X���$�?z�a����P��N�����ӫpC}��LG��*��q�M��7���Zī�>��J��<r��E�p^.������@<���-
�x�覈@+O���Y1�ٶ��9<t^P���k�`=���5G��ͣ=xծ���Y��Ge�!πd6#�7��V���X;�dCG�v��S�H�A�Q׵-h���S���B#�e�q\����WQ׳�^���w 4_Z����I����,�_�5륞�+|�b#��WC�$?ų���_�������L�<�PW{�;b����]������vA�Խ�/J4���K}�?�axdw�g,��y���:ٳY�ܑ	�/�����p���E�^y�D�p�S��ϲj��ߩʛ7E���[|QDwm��!�,?�b����?��'��g9>Hl�H&��~f{A+��΢xY=�&W��im)��'8��m��up�03�g��O	���"��_�`���S1r4����C*VR")#@��*T�?wJ�1;��g���7��A��ʏ.����L�E�C�f�F&����,\���j6��\W��
��h��#��Q�?1[�kF�Rt�%d�\�3��$�R����gt��F���=��O8K�aEE�5"g��ۦX�bh �5K�Y)���5��zx����9Z�0PG��$�ٽv2�>̾�J��ٱJط�N;X�2)���9t� �ϗ����_���8d5C^����(�K�%K�$�F��L�'ۍC+E��	����WA�Nu��5a � �֝�ϗ�o�I�2�(�*Ә� ;ag͐z*6'b�+��Gu[�x�;����BG�u��'\��F���6�dȼTG�����`���w�<��e��8���́|��{t��2:i3-'eI�a���c^G��͏!� k�*r�!B�Y
��P6r���I��H������a��Z[�X�"����JQ�shG��oQ{_�u�1̃\���&���;���8��@O8-��`���QJ!"���ړ�G�8�k+dz�ۉ�Std^x����ïd����c�L[�&L
��{r��^�TQ.	��O�~�&�iֹp��ե䤖����xf��Rku�����Rћ� ����ٓq���`����Y4;��3k;JC�������S>�m�*��N'���0���ʗ��"���&6x8�o�l�@�㹯f�k���nr��؞,���f�2~sÒ��o�İ�?<�!ю ��/7;t��J^��� �[�n�ytY(9~�+���]fA�97�T�ZR�A�6�8�s�������RJ"ӗ�;an�����Xn���������LWl'����9��V��W:�E*������|�<��(�a��T`�}�ْ�|��&&^,~���j.� =z�s5ڍ���PfQ9��/�
��������~���>U�֎G>�6��y�p����ՉR��\��dN{��X�^���I����,Wޤ� �<�����T���MY�VR��4\��A�B苌�)�p72��5+�#��r��VjQ"�Н�γT�cTʸ�x{"��{�h��;(��̜P[��S���HJ����̡��f�ً3t[��5Sgf�~Qj8Cs�/��%��?���.n��p��Z(&t3^?ފ���M�l�<GyH����$�YlΈ�&�K���v:��Y��~�mWyc[�y�1f_GM%��+�T~�7�Ɏ �� �OL:vgg���EJ��L"���^���?+��Q��}Ebh�3̈́*-̄-a�~ʁ��
��/�^\U�U7�*�nK�?c�g��!	H���8N������k�k{�M�=�(I��)?������m���AN�z��K��s�$S�4xZM3�tr��S.
��	`S��{�V�Y*=\���ͽ��;i7K���-�;�,�z�GDU�̖��X��Ab<V�RK<���2�Jw��;�&+dEN�W?�d�^-��ރ.dN�A6"���-o���	��@K/������u�}W��O���4Oĵs���B�?�!k�^��Dp VUQ��b���2%�*n����l��'���*�j� }��U{XLb�7*���&]d�?����]x'�ɨ7P��<�I�,�k��QrK�q�2��)@8n9X���A߹^A����o�򘼐.�cH�jhK���4�o�O�lW9"��y��O�<a�㿥�&zló�ق��D��;�7�yـM^�i��k�p֭h����H��=3��>T"�D��s~^��gUy�C
�T�
Dȁg&��2�r�gu�6E�\�J�Y�eE*�?p02�Y��w�n֑�>�Y	S���r�U����Π:��>�\�d�!�Dڎ���Un��dXe��H~�f��^s��o}ta��o��,.]�['}%441�<$N�qPx��:��Q$.\�\�HJiMC�s���M�ن�eκ��Nt#?t�s8�wD`�g��EF�='V���)��٘��(���Z���Ƹ7jB2P>`�<3�=�Y�{<Ϫ��'�P�R�t�$��>;b�&A�V� ��k+H~R�����&Cͦp��Q ���7�0�$�{V���϶����r'�2�;2� �^���Ȇ��=y�46cw-V2������S4}����
�,W����ϴ� ���G2�
j�YBU~���u'Bf)���GJu#����f��:�ǿ)�1[Y_5���Q����ͷ�����y�p@�@r��\徘�Z%��9-b9G��-�+V3j'�O58W��F����U�k�&��PDH<P��y;Z�\u�n�y|s���˲���^V��~�"Q�9A����QI�)&[�
�:���M�����xqȑ-�� ��N�S0t����`���.E�g�?��I�$L������;d�4c��,g�����1�)sp���d�=N��_�m�r"kXID�����c}X�,���&�0Go�* �Е�$��h�PkFC�u$�W57���D���{��,H��T����:�;,�vg�@��'�j�ܗpcddBl���o��u��b���fŵc�ٜrn��aϜ42��x3Y�b_k�4\˛M+`n��f�_�lj-���O�rd[@?<�:2����m`T�冡�˱����ztt<�3Ml�d�q�v���7ǅ�s�})�3°VK��eH@��{�����ҍ9�\��|�k�@����h:��'%3Ie���cE�� y�ЬYl�+?}���<���:��H���� �3Y|K�4r�����q��"*>R�ٳ���59�Y�њ��M����34����u$�ɦԼ�n����X=�ġ�R˞O��" %�ҭ�l�z���+E�AH���R�P�D�=& ��V��$�s����VE՛9����V�����
 +���-:�p-I��Pp۟>��':	$�C�F^���x�i᧤����X���5���	!P�y�[���#���f�+�H#B?	ػ��/39�~��]%vW�z]>nh8���?�AV���ޛ~x�P�t����pbW2�|��Ǽ��2�_|�#��S�e���~��;젪�������W��c=7�ow=cJIP�tb�n�LL�0JA������!��I�T�כ �>���@�RH���D3�N��Y��a�A�QK�Yw/˗�&^z��.X�4��'׼:�SRE,ƭ�p������R��$��ͺ;nܣ�L�i����U��-^�9q꾕|肥���r�j�M��e���*��Y)o�^�S��3=�}��$�Vzj��$D��4 琞p��w����g�eݩ&�lv�l�����k��K��"lR�̺C�1275YGs&�����3Ot�Tj���1�@�d��k �>��P"~��u�d|�����MG���J/��r��k��n^qZ�a<%�s�k�{Y&�,{���ђ��E��.�j1v^������c����K����FƑ|�1���V~"f6�6���1��tc!V�sۮ	���9����-��Փ0i}lc��鹡ㆼd$-�x��3L (���Z�1�i�}I]�8̟��(L�B��	?��S�k!Ȯd�Κ���>���S�I����w�&�-�Z�� C�נ/�ٲ���B7��wN���V���@��;�c���+�t�;���Ҹ�J�4��)��6W�Z�;l�xan85�p���C����"d�$.t�1{��Q�e�=^v�+IL7 �"���Tn�!��GE@��0s,L�Q��z�8�\;^�؁���������蹗)�t����M��m:�wZ��|���N��V�V�h��P|��;&�ݙ�i����_"��4|4���)%�l�^3k'�`s�Y�Q,����~
�k��ak��U���r9��+�u��8�#�����MuK�
)%-�(����z��Lȼ�ѾM�_�gNi�^�9�rvO�����q/�z22�%b2�ͿRM�.�m1%3�n��T}V*�w����nH\�lF��p��B�RG
tp�U�rސ,�ذRU����EE�����8ku>a~��	3��?3��{I�_��-�UO�[�4^H
8�3��:�bbX��gg$9)�h���'�^�<����_MFh�*pA��Ȼ��p��b<`�]Ǿ����dHD[��O=�)�,���8�7�Pޗf�-�@���+�+���|��F)�r��W��x��z?����+m���h.������Yg�/�W'�`��|��h!ϼ��|� �n�owY4���f
Rτ"��m�7�S$��<���HV��{L1{� V��m���792ŗ���b0��uY�[��aū��x��cV�i��u�����W���m������x�!�~P��1��0"��7Z7n�"�~����P�kj�*HIKgÆ�bZ$�͍=a˗4���厣�Gp|t~=k�����&p�kd���E����;��iB�#�3��|Y�F�w���ƣM��*�ETK��9�I��8�^��Yǹ�)
�66���8e�xy���*3�lk���%����ا�Z������c�}�����@��[&�>�I!T���5����Ȭ�xU�L��;jۄ��ط!�D���CX�zI�����+3�mM����Hw�l��O-�E��o�S�{��^�ez=j��qt�Kw�� �+!�,�H�0$y��<��3�]x9;Y��Ay6D�S�vO�cS��0%��ˣG]Z%��]���_'Ұ���Ԁ ��O�W�H6���gþ(� ����f��9���U�G�/A\{Bo����tց[�T��ܦ�َpV��d�2AU=m։���;���uB�Pi2]� ����%����])HmD=�I���N
�����$�HH�Z����
�g��{����B	��`���{#qO���J���	�䙼�=b�I˭}=ڨ�he@�%��B������݄��9+TF����yE_k���i����5z��E|�K�V����0b��ma��j�BvHHi����6�~~��Z����}7�����k�o��,;�YD�h6�j7\�{� �?�Þs\�[��%hixђ[PdiU*�6l�I\��#I��#�Z�Gy5Y�����x.�ǲ5Ƥ�1��o�U���!���c�x��z?c��%D�$�@��r6�X�" ZU>Q�#�WÍϮ� iH~�V��y����P���0���6��Pͻ��2q<����u��@��q�I�=��\{J��������	���ڽ$r#��H[	�훽��eR���ޣ1�x����I<j�R�C�#y	]:�h�$�<z�t.n�,W>��!�p��}�L�H������!�)�|9v�9_�� ����x�=dIP����G��wC/[�<�%v#�J%�37X�)�I}�^��<�~�$a�S��6�D}�G�Qh�8���� �B��[��ao��U��!RHLOt_tbBB��һ�m���E��^�k�Q_	-vb�;W�7���p�Ss��0���N�Z	�n��+j�����{����P��Ȏ֐���
�0O�<!t(�Jg�X�^�
"����-nT$�V�MM����TS��
 �����zu�x�(���]���V��_��*�»�_�T%�K�ߪ�P����J��a��ǆI�S���177w����uw��
%�����M����J�<���F�H�C6ԝ���<���`)ԍ�ge��Y����1�:Z��:�V�"|�3g�������7�Zd��B�|;R=e88��$��O�������x��Ȕ�({��J�X��0���qZfHc7/���	z�H���Z[`E/	]����`OQc��3�rـM�j�gL���ţxG@줻_"�z�q�j�tr�V�u|�)B������~f��-}��N��_+v.w��F��:���k��HJ\!bU�A������n�q>+�����c��-���l�����!6㥪\�8j�"Z"��UA��R@���g�	�0��Y]-�Zm�2q�����t�ڋc2��/��먠��U'X�W�����X�g�?!}�(����(�&�z��1>��/���{�@0:*$\�[�_|}Ҝ���5G��@J I��6���fЀ�����5�>�:Eg[ɖ{���%��g��jZ]���2�9�k�N�2����$�"!���8c��e`�Ie��H}i|q�]��<��v��X��7�O�qOXD���F��US�GGJ�n�-2�4�x$$�}V��y׳C�~r~l��G
0ڠ�ѡ"`�)U���1׫AV��%%j���H.N?�ڒQO�t�yź=���T,:2��+�H�ʾ�����8*����X(�6����v��j�1B3�^'��)�U���!b�/�)����r���j�$�)Z�yWQ�H��N��7���^9��P=p��8�i�JTΜIz�K%�A����ڬ7�5$Y�?^J�Žr��y���q��ix�k���A�"�0�o��+�L�A��,Vd+ly����_�����M�(c�ￌ�>�d�fi-5k2=�����9ܧm���qӳP(	8�@�m��gRP��I���e���YhLQv_�+k"�γm�X�YZLA�k0�1�&pp�:���(*��1�$��l��j?g����	@����BF=c����^٪yB�G��Uxq�;Co��3B�㯧�]��5��Y*��ʡsNc�f���b񲑳d�#������MZ��I��Ŭ:0�cj+���S������p��k�<g���7�|Ul(�v��r��7�Cs�F��糠�n�}�Y���(��}e�X">���Y���F���YW���}�X�����)t7��|������	�Ne�rd���� ���b&;۸@�L&x�]oZ|��A�\]V6�1��46�D�e�n�����dϠ��I_�,��[�ôw������:�ޅi�FZ@��K鐖)��$$�$���閎���!������^�����kÂ����~���>? d���6-.��P��g�	��x�k+�p���
k�S�]�p�N�U�&��K�I��f��S5���;����"�խ:1+���eI{;<���/W�@l��1Q����Q���S����w���^bGSI�"_ż�����elX��vc�g����8%���1GS+�Զ;����j-�z��b������hJ
�
W�5��K����}	�����EU�=���X}�L��8����R�
��U��e�ɯ��
!�s��nZ�Ƿ����u�F�}J�<���U���\F�v:W<z�ʧB�:/`gW���wmi��f��WW�a=��|3�����]�_XK<���t��p��]d�:���}n!ӽv2�3��Ba�ò�PX�,����zj�=�̡���2L�R�i�)6�����'�\Z����4�w���/֨���~=��m��BC�&�&��ܚ�Ȧ��i0w���Lg�{�:��8�(���tΘ��Q<,)8��̽4���NF�l]�<J]9���I���+�ɥ��������%���1�6�����݊ؤYe�%�CGqOm��g��iFZ�6�K� X����M�O�%�)��g���"�����n,RWp�_�2��t�h��5�&4;$zܿ�W���2�m��	+��f4pܷ������(�p���]܌�5���L<S-�m[qV�Q����V�2�S���h�?Ľ��S�c���"U1Cޢ��֕滖�:k���ũ�$��Bؠ���x3RQ�R";bۉ�X��#����_R�2����B�bJt5�������qcjoE���z���f}_ېښ��F�
��f��N=��m&�z�0&m}�ai��(�I��ͮ�{�/r�2�������	T�Ʊ����\T��U5c^��w[�����ʌ��5�Z�w��}����.dP ��O�f=���0��:If@��pO_��7�7<��)#��5�ƹ�w���djY>%�F��;>^쿒J��m���iɩ�^�ݴ�;=����������J@��D�16lo����:�E��p8���������^��;������)se>�/����
1�0�5Ql&��v }
�<5�i�f=�v�ݬ�>Ϻ��)j�W"���+_����gm�§�n��6 ��>5;u��E�4��g�rgx�6�j9K�l\YFI�}H��p�f⸾�1f�:�w<�۰\�����q>�����������+����O�;��!�b��d<�_i��s�+�9����0�豠�%,�C!��]F�F�Y��-8�}��o���|Ν�>@/�L���ŀ����Q9� ����,N�5}�꼮Z�`W���.�Ko^�ś]�z�~Z��}Q�`���|Gr�x?K���m�J�\(��20a�O���|}d���o:Q����ҹ��c!3�p*�'���)��t�w9�ߧ�50i�^�m��3�H� �_��
�O�LM�1��:��g.Q@�v�p���U�li�n�%�����S���x�7��L�1e�ֱ�ZB��������":s@�5��I~#�Y���f�N.��bO0[6�z|����}���R``۫1M�&qnC��~���U����E8�2�,-_�܁g�|�O�mF�~�r(�K�	��"݅<�̼�V�F�b���̈�������f%��l�J ��*���m�W��z�rC}��X�/��0Fv&z��U���#��݃����+�?"������+q;��&���A���nX��Ĳ�h�x��l&F�|�D�^|j�\�S��C�y�����e,��b<�T v%)�,%��s���-J�Y����_c_t��b1�Xk����0�	���p�*"��%�������2*)v������#���m6��o̭�nG̊)(`H�j-"�|a�����f,�|��V��ETP�xK=F����~6�*g|$������A�F�����#i���IC&f��7�^��9�=�-p'5e2M�J�/���$�AǧkM��]��&�L7�lH�N���s=�v��g:c�R������qD��!blV~�vJ{_J�Lj�S���C�7��2l�=�5>p��xm�̔���7#�����@|��������;�rэq_{�_������uD�J;���[���v���k�e_���	m[�=ᬐp�%�����eD
�e��kw�f�uPV��`�G1��LP��>a�/�y^���Ƹݥn��|���&�M��֋��4�?��~+~���.�����#�ZuHsp���um9����#��/�vI�P�К��<��RH\\-�_�����؞�W��5{0w<��yH��U�jT؜HL�ʏZb%���� Ri����'���Y��mkT��`��(�&U�|�f�7��1��dxd�6���]��J�8mAfB(���N=�?A��5�-�����<����zE�P��Z�\œ_�@�_}7�z�g��+��+�[Sz58����V[��BժRPo
�<u�45[�G4�7Xk�S��c�}	 ��Q}<>����������u���=���6SլűM�ݮ~��犕ЁUG�b+jB�Is�p6�
��X�cKyg�L-B�Xgzϣ�xH�W�����.�;)���2B��G����\^Wե��C�%>���kc���w���F�yKnh�>dg��ٙ��=��߫�C��P��ׯEkR+��;�  �S����M*׮4�Q+�C�{�袜�6i!�sy�W�u{j��X,Y\-@7[���6��iK~s���+󖫵�6�-����'�UȘ��vl�ؒ��?#�/�;�"�~w��ؾy){�Ir�Z�!��4C�{���қ%��~�@@'�a�s����o^RL�\���=�op�����&�;kT�u�w�4��`�c]b�yOOhg�B���vTW���4r5�_!�Hw��ڒ���6����A0���[�^A
��.kK��ұ{�0�:$�V&�ag�����2��kt�po'���gUr���9�w^#p��p�i��R뻳;�Td�D�9�F�c�(��Q<�*m:@����c[pj?o�ro��b3��/���5$J�V�����n��N]�9�E�/�o4���ԐV,��l���U^��kꞻmʭ5��إ�,��1=Z�`X�v((Ѯ��hQ�fU�k��A��s��SPh����O(�{�,��F#���Fy��c��j�����g-e#vK��k���	r�#_/1�c��õ�1�y>�|�(�P����S��I��6�O�T��1>L�#���6�S�{��3��J�V2��f[p�����᫟���j����tFg(�m�/�ˮ����Uu���ގ��2���E�n.��+�DEۯpP��_<�ZbxE��7k_�RJuo�՘X �'��UW?7$BMzpMB�[�rT�fk����������^<�hJ�rY�d�!�q`����a�4hd�I�U�m0��D�@ϫ�-�	y��m�|(�㶔�����0��m-7��u��:NQ �8����FX�lrk�����193�{�V4�|��zS]�w�1!�.������Z@9�
]	�j�A��IQEO�b 秼��|w�^J��@��N��0�"��wv�/���W�`ln��JV9z�ZJ�\��,Y��?�W���#��uR�e�1޵W�:EhQ;EG���~��K��;��
۩�E� �����~)uگ?/�� �;-:�&x)L#���X��?���jr��B���ݹ\��!�s�a%���;xxs�D^��感ԇ�m^��|���ccޔd�4<�61G��v}T�F�u��Xz�
�a?�̑�U[�x�AQD��3l�1I�����	!Y���:]��߀��_K��Z�$�mxjb|nM�7���&፥��k#Čd������"��Z�>���o��4�1Zk��5�ЄN�ۮ�Qv�2!LF�8�C,^*&��W<�5��,�_�f�����ӂ���I6A����Q\_�Vۋ�$!=^�d����1pTo����/u����
_j��.t$�%��zv࣋��|+����X^Y~��2���W*)c7f�Z�c%�F����i�:��;u�1L���oJ�Rf�VJ���^	��wx�6T2&:���|�0xh*xj�u���A�3��@�S�b��f����;�>�0E���uU�Y����!<��W�����)��~X��p	�<4|1�Nݎq���@i��؊4����k����`�s���ZL���6K~���m�.����0�/Eы�F�DJ��; LM��P��=��-�H&��JCJ��o��?���^����aK��QFڼ����[Ip��!��/L����]�wo\qY���^��:zg̰�X�$mmͬ�SK(7p Ӽn
���|���l�o�G	��*qj�<"PK�Z ��T���"��%ʒ΀���9�#a�����8�#�ah[�T�I���=�6,����Ypo��-G/:�+�d������-�Z�hmrɺ/P��^����y���T_��{��N@:�l!�R�����mP/Y���vV	���������@1+5�����uw3$x9S� ���dFF���;�;����lK8x�.3No�Bba<�ϒ�~��������7���E}��;8���y8��{a�.#�K�6�!��}���qń��<�
'�8��%�)����_��ب:]Kp ��oO9����4��&]p��"��A����dv���U�Ҧio�|7^����N�2�
L��݂Rj���?A���Mh���o<��)�ߊᣮ~!�Z���j�]���0N��S��B����j�~��a�;?��[G�/�7��O�Ku�Ih�LT�z� Q�Իc�G�T��{O��J\=L�UP�@�/�f�98�;0��"&��s�����́#�zi�4dһ�N����UhQ���H�~�G�����s\K��
���X�A�.��n�����5�'���ݑv0`^���Կ��(~3�W!h�,���e]�o��8�����Ҭ��ɆJ�1�@@��/���s�c�m��)�7)�OP��toZ採���86�#�UM��/��X��\봚�v�����hH�x��3�ʺ�����^N���GA�w���h=���2���?�$bP �7/+��<�!&���}d��VJ;��'�c���m�F�П*�:+�~n��/@�m9&U���l����H<��Hɲ�o��*��,\?ۂ�����/4^Hu�ĚK�4P�C�3t��C�6z��vVQ����Tb͢��N-��"B�8~��;ܵ�IxL���G�|�C��<��P��ӣ���o%h�/�zD�9�
(��붆'g'3��!�b�?mp��J�ٳ_1��h�3���S��d��%{p�����8f��k��=-�NW0]Wk��b�|�� �{�����\���F�2X:��/s��N m�4b��b\�����h�;m2:��t=*����NM��|z3wZj�������[�ɢ����̹�r����p���h�}�Ϗ��,�g�J�F�'�:�5ml�Q��M���F�4,��#`lX�5�e8�bN3��ᾪ�W��y�:��YW@���*ke�N�|�@�?w$�OiP�SY5�z�H˔�-\č2��6�Z����x���`1?���Fo}*���ֱm3�݈7;��j�0�Ҳ⯷���d�nY>1�J�y��s�8C�'q�ao,�w�6����1^<{��m!��œy_���aYA��Z���
Gkv���+��8p�����C�:Zn_8���~������ �>vd�=<��!2��`�D��ɸs�����߉�5y���?�©���tkЕ�һ���w4A�2��m�m�٨�b�6��
�f�5�b�����Ryk`����J�M�?�拞���`)+B0�h���b p;B�©�����}t�n'�ylkql�(��-PqX�l�m�K���9hsR����/�.��|��	�!o���@�};)T����S[�>fJXlN4tګs3�T��Ϊ�s8"�UDBZ��kj�ß��@��ϛ�ѡ98��Y�R���`bКȹsP���q�6Ӎ�D��G�J?O�#��)+xa׌�@�����ep\�9{��&1Z�������V�gL�2'�rL2I��TRQ���xo��.��F��&�uM�6o��w�#5�E�lJe\q��,�����i�<35 �F{�/%���ծ÷@p�/vj��nf/�C�LO��	 ��Y�/큈pf��L&�+Tu���`�Wzk��ί�vO߃#��/z�f�I�Y��٣����>a5�SO՟KLN�>��=�%B��d��'\nP�c�Eb��n�kT�9� 0�n����h��x����<�\+�(������g]tBc����S���t�K��}S�ˁOq ʴf��>n�1v�9�蒳�TjW%�y}���*-�zFS��g�؍N/��o�㰮�(½�:�<i�9��������y���e�`6��v��x%uʓ��G#�2� �/�jf�Q��T�#.�a.�\2E��f��U����б�A��Jl����eL[bIL;r讲��p��\�-I0uXz��A0z�������ë�l��kF����<��^�=�,yf$�{PO�U�Έ��O֑���i��?,	:�b1��R�U���n��{� .�uG�|�Z>�\XJR�!A��=�dh�tG⹙K<O ������Z���Y�v�`,���c�rY����BQ�&L��2�:��{��1as�/�ݔ��F�Цn�Mj^$L���=���͍<M�@Z�3O@��&Q�Y�����r��^W�q?�������B�2�O(�������p���ɺp�	3KM���y�5�����e-1v1���Mc�,�y� �B����9�jIJ���mt��u
��f�_Z9�[m�Ʀ�Q���ו� ~�ٵ�t�n��g?���	�P���e�Y0!S�J�X-�ڨ�����dg�M�Z�==F���B��e�sI�ҵ�������vq��⍕v�g\+�H�N��ɻ�^4g׆W��R����ۊ��uX�2"���٘�k���=����2�,��F���?�*�ڰ���Ϯ�O��{��[iП���v��[e���-�CA�|��}��&`�"İ�B@>�$��[�V��KM�i�ȁ�����6������'6�q�'�B�kA��l��;��*'#�b�xţ[��[�#�r_�����3�,�+��I�i�гp�y^D�F���{J�l:
���[;���������z�D��y`�
�w�Mv��;����U�V~x(�?�Z��^�������Ϸ�^���ֳV�BFg��O��p�*�����s��Z���r�+��w�30x��Y`��4�¶��H�,�����&1��c�����q`�"$��#��fZ9W�t��z��&��i��ÁS?��fǵ�S�8����_-�{o��@�[�k��oh0�{�ݜ�n&`xPK��1���xei��elJ�X)�|�e��'Ã�؆>w������2��v�s>�;-�tީ-UgT��b�9H�ܱ⩉���+_G�Rm��mJ2,��jz���#[,�4���3K��N��bJ)پԶ��	Lh6Pc:�I/��n����J�53��S��k�?��gСg����ڊ�k�ދa��'�ߌQJǶ�n��=�v@ ��#Y�U9x�~Ӯأ��RA��iSR���M��	���1Ë���b�4kߐ��^)l`��-�	C/�P�-��\r�Шr�$R��o�GEb ��F-�Ջ�a	���Hy���WK7���R�R:L.���h�-[d�^J���N�&��y}���D)^Aѐe*ܵ�*�J�6������J���*G�/��Ƿ���d���z)(���Ѕ'�S��ț����E��g�5	���;<<�g����U�����m\�1�FǦ�.]���R�k���*�l{i���s�>�5��(��fy�T<��^�a�E�g���1��rZ�{�
\�B�L>h�X�B�$�2gp��SGo�ޝ�n�s�@��5g�ԟ�+��w$�`�O���:)
�g|�t��N2�ʵ�ﰟ��[���w'��͆�cJBR�%m���o&�{�u��?���\�v��|��:H�l�F]k��vF������/�m��x�H^=n	 kݓ��ѽ4�k8z20��*�.�a%/U���┣yw%�����?p��������0�����Tm�wwi�����R>�Sj����O���۪�aԐ�5eޝ�o&N톽F4�U1�1�����	�H���Ǜ���wH�*�:���zo/�%���o�FZ�$������%d]�/��_e��;�;k�zg�aU�18�K���7�޾R��V��K�B�qj������Ahv?P.�i�����n`��v&v� �^�����}9=��a<h
�<��S=�>W���[ d�[�t��n�{D�Ǯ�&�Ӄu�M����>�L����%J�V"�Vv�.�T�d_�ʒ�J�BɫOO^��L鞢�,L����?wn�@��Q��?*-�	Q���a2���s��7F�in&f'g.�35UÙ?��lE��^�rTMP������i:�!!/Лf4�N��8}S���rHp�L�픔�W��<��ܼ���uG�0۹{Y6w�_���ޗO�������)��V�}�,E���� ���I����硧 ��ىv��Q?�A9d����=!:�+��� RP���y����c�&�0:6�I]���C�^��v�ʥ��{ҷCZ��:�@&�R�wr��'3}�P�i��P)��gh�� w�jw%��B�����M;2%�{~J����װ��*k���o��)��F9��&�FF.���P�+G�!���W�*9ܹ[bG�|�a���C�0�䮿�	������OZ��F  E���ؠ�{�c1��'޿�(�LV���O����` ��Q|�(�������ehI�!z�N�W`c>_����ar�?Y��W���b�(!7�0|#Z����+��C褷gMk����v����x��W��!ӬQZ$K��2���ԙa���zcR1�R���=/~Q���mg�օ��{���\!i�(��U��𯏙��h��n��ES��5i|l	X9�k���Ki�L܉*�0��ȹ�D�iŨ|�6�������S�zٗQc�4@ɱ�̹�A��2c����0?�/�!�*g���5t=�9��ܓ����̔4�ˣF�hN�Q�7$��k��v��vL�Ȳ8�-
R�r_���xFU����`廽/OT�)��󥦁A�ǖ����:���gL�M�&��I�0}����G�ui�P��`kÑ�3� ���U ־�k����e9�/������y�����=�*�R��|r��V��~�~9T$�����3�����;�0qA�j[ߵ]ur�M�fl�]�5������Cٷ�y��?�/=�	V$���%?��7 �:�̜'T���~,�ڵn9�GȾ�V�Ϭ';�����e9���&���# �=�sf��a�ftɆEBb�>�=t_�1ci&�B�6�
#�\Ú���B@v��"�Q%/�H6��־'�Ɏj��N9J���v��|G�� '�6p>o�!!���޷���\勧�(���L�G?��y�"n��RC�GV�N��n_�ܔ�x��P��OG���>D���Q�,�G�S�*)�/�=��y'Y��Q����B���� s~Un��཮���H� �_.)��9�1%��ڲx�,`yO2=�¥����K\gMD�k�(⅏�Ԟ�V��P���Y�;���r�T������S����!��f���it�b)���v��8���P��iV�+@/r`���¹OJb!��G{yT��+�?[��i+n�m|��l�i�z�4��q��[/
��c��;H���E��%�[|�γ"�����YU�5���	P&a/$d@�������0�6�0�xj?�/��8���G���*_��kEiMԒ3�vp��	�����p4�j�В���YXb��|}K�l�ԝ���@;M�����j��b�p�n'K��	��ߜ�y�Ɗ�-�{����~!؀SX������'����(؛I��-�W��;�'5��ڨ{���Z��[Vp�h*�<b~YW�����3h�f"�1��S�I�.�W�+eKgX��πo?.�HM
�d�����4Jy=�$���r�y}�/%�!�g�u��߲��oZ0�d2���3>���^��4
���O���/�ӥL3��vV��������Q�Z��٘�u��x��7�#/|Y�l�*���yyB�i�~x((��p��Opdds��Tڽ(��k!��I��RO� 4�B=�ΙZ8d�q����p�*�'0{�2@R��ՠ������km1�!e���[��<���}�;x���'͖k���0�6[ZuI 9<MrP^��B>�c���C��Y�@W�/=����P��2�WR�J;�ʀ���j{�e��<K�x'������rh>8�r �ɡ��$	�����������
m�Fh���K4�9���#��Bn��]R)���p�*X�bMv�.�Cw����#S���cs�gG��m��-�=ӛG �>�E 0E�=y�5=���a�ʦ�3��/�����k��Ji2�R��Z{��dM��c��u���	껭�MN��J�8�%�"�&��v]��&��Fie�[�f�_��k|�R
���p� �#D��R��&!1�� j����d�V������F�@������z��ڥ��m�)���67��ߵ/��;),V "��p#��Չ�@��zQbJ	���Iw��U������|�����l�S�9ܘ���o=�L쬴�C�l��W�����	�$���<|kh�9���@�Ep�Ĭ�L�~޸)@r�����S�t�ќI���S�W��Tx�"d
G9�����1[;�J=���@a�<�����r
1���5ĭ�7Z��q�Vom��tn�4���w^2~���X��;��)��΋ٿ�	�M��:�'�\6,��՚/KX�8��C���v:����'v䩷�c��H	d�j��+$Zğ+���g&����<��$�L���~e	N�	 �Ψ�Ȼ�$����ގf�1l�q�A[U����3y0��p�֘[��84+�ZmD�.�?J����"�#�+�-�@�&-��G�0�����uθ6��&����ڑ��C�-��ţ���Qc���TXi��WR�_���G�w���&4�8N?w|i;�)y<^���u��Ħ��䚖Pk��S��L���X\o.Zk����<NJ����ֶw�dN̝� q�-=��q�XHG9O8�J� Z��l��y�۝/@V-���桞\��7�q�n����̷Y��qk>Y�L��6�O./�2�����h~��pX�=��E��wxt��o�"b狨�D�B�U�ފO+[m5)���Q뢼o��U@P(&h-��$ξnPK\�` �.P��>i*��W��ӂ#x	���NC��^km�8�R����,�
(�$
vIP�5\ 8�?�������`��Uۺ�4�ib�?�˸�$���OJ�xq`Sz?�o������%++*>��)&C�M��7�R�r�v����8~��~�<��}F�0`GR[�G�kPK���e@8ֆ����H �bqrk���P6�ϓ��0'��3T3�^~�/��`�A�B�ul��d/�"�E���k8�
���幩9���5�޼�����gJd�Z����xxM�0�3'���*"�������0^����x�tn��sJ~��&;�0����Z�J�ۢ���i���)]yE�ua\�zN;����\\�{kr7��Q��E�0��ݴ����	�n3R���l�S\\�um)�/��N����X�Vj[�Nv3R�A��e�d0A�
�d�إIo��^C�u��_k_M�����UYTM��wX]�q�O���y^2���P�I���w�2�B������ݷh�S�NP��LФ��-�,[yɊT ��+��l�ڪ�?��2>d���t����Q/�!���E�Q��	\��Uq-��E�K����	��#�C���m�G���ш�^��e������F���>�����v�7��#���;:���j|}\N��ݟ��Y��1�����v�Ζ��]%v�M����OA����*_���,Wc�Wo:�)&@�N\����_\�Z\p�|�i���駯���{�4���R����~{7p��lK�P�O(Sr4"����z���)j�v��1�J���oom��޷�=��� NO͛�[|�M��M���:�˜d�lpB��;�������Qh[
{�l4�����Ǫu��?lҸ���,��Ƣ��vL���Fa~s��!�ZU���Y��:XΏ��{�A�+���&ﶙ;e3�]�}��}_p]�l��O��f�א�g9s{��4�1�&�~�Xz����7c��c_�K��r|o�ƌ��@�`ٔ�����L�<��v���3�J�ͮ��� JA�w�о1#�)ݗ'+��2&�N�mb}�W����k�q_�V��g�t$�N�[/5:OؓZLH_J�R��A�f���j��&�{��Q�$T���͖���'uH��/�b{���؟GO�U~�x�s^��!2E��Go�G|e��S><�&�*F���G[�y���v:dIg:��1��Ý��+��T��/�0�����Zbh��k�C���Y[-f�q����B����Q����3"L�J�C�X)t-�A��lO6�`q"(#�Lm�ku�����V�ё8U*8?_&x��^�S��l��WB��.N��I 98�xw�g(l-�c`e��O�t�ْ�j$�ݜ�ħ�L��/����__�g���H���O#%�Ho���}��P$�u�:�A.��P�Qe'4�����zf=���M ��g����Y�@n�M���b��
���M� ����(V�,�mԛ��8ϧ�-6����V���b�����N�d����5m,E]3��{9���a�CHH���s]y���a�B���e:Y���pfP|��Q1Ǒ�`
*���������WD���#���V��xV	��m�ᤔ���<�v%�h��Y���p�.�[�0����_��`ҋ���A�%����b�1c�x��]���qZJ!�Po�[(D5����=�!E��׭����%�sׄ*X>Wny|º���}�&P����7S�)n�0X��)�B[@p�W��I�#zM�\S2v���5��Ul���W�;���7=�� �&���(qj?�+�vT���?#��
��YW��"��ӂˈ��~b���ԝ�IC�J�}��Vv��r��	�̀'�H!9��C[�w֜�S�@�<1�ĘO-������̂~���)���S8G���m%sW��x13�.A��ͥ`�;s/�Gq���3����g��E��U�.P��m��_mB��V�=����c�f1`�YPY%���]����2�>��
^�WI
��[i�����(2�@�N ��>��7bV��ӷ��C�����{K�W���23�����зl�-���(E�C���?<���J������b�*3�͑��,����η�q1�j���@�����-7�|���,�*� �Zuΰ�ѧh����:;;yw��sh�$���r����a�s����?�@�%��4Q��Gg7��ߜ���L����u�:�v�&�����.^������=r�;��q?>�&�_���.nY�"haMۑ��	5�tP��	6���������>�/Y�c�V�^���6�'Gb.����1���AӤ7^'í̶1�N��i-�FeU����X�&�b)U�Y] �l�?a�+���W��r���,ad�CQň|���"�q���� �!���K�U����@��"�H��m���E��s�o�m'���_�� �j�x���4�\�7���;=�[�������Aq�b�N�������4"��"<�����C���O��@L
?j���9\�;a���+���!��aJ���Nrꞽ��OF�eZ�h�;�Ż	~A��{
�^1q�n��W�9�s��콕��#8��:>5�fy����7_HL�Lx����l�]r��m��XkCY:���@�5QtgZ���f�kDxb@�uR������c��*�%��N!+�JЋ}	,wQ� �E��f�ԉ��tl>&1ͭ���$��k[��܅`����C1Y�\6�����;�c?f�h��T�%�D�N}�!��_e|�sMY�βlZ�Iyt���BQ1Э�������X=��p�K����"�I6o3������yJf$�xļ�Q}����x
q̔0�@��ԑPM�m�'�y���+�:�GY�A��!�W�Z���\<y��~��t��D����t%�,~J���I��c�`��Fuq��H氍4Q �i��'�{1\�K�r����� _��'~oϛ`3�᭝+o�KΦ�%-Rp��$�����i��^V��┮y`Ȕ��@���M=��A��F����R�� 2��6�$1���ըi65ER�i���*h�:A�?��ڤya����.���L��/7�D��[����L�@0TX[��t
\˲1����*_��Z��K���^ҕ~a��M�i	�ܹ����z�9˸�z���m>1�x��)�W����ЀE��و;����Y܄Ѳ�}�3I�wy,w�({��{9�$�r���$��o�E���s�kEJJ᭮�\�?��5���!s��"];�l�۷�"yQ����C�i�O���V�ޜ�X4����I�M�Er���1���Ҕ��������s�&�2�b��ο-3��������	��-���A�����C��r~~���p
%��]2�ĥ�>a���%+[�{�pu'��4�	��x��?	��5�_�Զ�KQW�Q7�m�30���i+�;j&Q+��=�H5��rs�x��0�C�z��0�v�$r��W��s���yL&��s�������κ\X���7^t��/�kk;�[�z$b�:�t�[\���o.�	L(07�=ފy�bqj�� x?@&����4�F��ȩnҮ��w-��*!�:�,8�I��UC,��y�?�w?����r��:m�Es{��WCv��t{w�c#�Y�<���l��s��߶�S�A�<ռ�x�t}�Au�X����_��<�Q�3����/p�t�\�%M~�^��"U>҇zQaKE�����s�xSv!�{3�7"���`���������$��3p�zD�g�"���IS"q̱k��4�!Zz�5@��khG�!�L�u̈�-�m��� ��-�,�����"�RP����Q6˨���$w;p.����Y[5�r
�Yޠ�B��.��},Y����}�bh�&��A[[����^-[j�x\�l��eܡ��vlT��$��ʖ�J��J�_2LeA�ek�����R�=|O�-&O~���q�@>�a/������*��1�*B�lu�Qy�6�/��:�ɕ�BK�S�dzF?}��Μ>�M�Qî�Z��V&�ҍ��V��c�h*�_3��>ˮ!�Q5�c7���;}4 +(b��L1o��3CHD�9Β9�4����wpz8]<��U�Z�� ��^w�1�Z�X���T_|�쮳�ou #6A�␠S�{F+�KF��/:?�B���l�J�AF�����Y.�q���m$w��C�bC(�7h3��U�O_��"���f���B�5�/���x=�r���hYᇛUl0ԉ=`Jf���u�`V�B>Pt^�zC���P�N�y��Y��M���<�,�]���CV���_�g���.�x�@�`y�����z$[?Zn?�xq}��w���s8�%��������/���m=I����x*���ҧ\�WI3�O�^X��@ ��ST��>��[�w]��E�����3�7��ĝD�����̴W[s>�9�9h�x�� k�;�����=e��B_��'��Z�g���х��o*^�l��x��r#\�칣l���ES���(�x�βyJJ����j��s�@` #�T_���lw9���D��A���DQ5��������?q>��*��2�Y�SwQv�.���%?�~N�\���x���x�3<wl�����&Y��X����=n������Ł���h�
�_C2��U�9.mE�2�T3CI�ێ�-qs��Ƨ��?�d�q���t�z�t���(�7G��u�HJ
n�)��~򲵿=�I������uM���དྷ7o�`�+�G0����hnS��fg�N%<	�q�áO)�L��<��`f�OVB+�p%/���ˀ����9�&�Zʆ�
�(Tbh���-�%Uk�_KFG<�s��Ё4�IG�h�] tڧ���A�����K��,B���l�Xl�j�=/Zȗ\O� �8P�wl�$�}!���Jy�����,e�ep�'9^���;f_��~|��d�0ۿ�ǟP��;�2�iɏ^��p��/ݠ�s�m�Y�]ݴ�ƒ���J�[��l�Ϡnp̝P�)�1k�4>��^ڏ�
ep���W>B(v���z*+ZȑbPDdz��s�}U[�pR�0����c��i��=<�T��,:*��}r��K�Z3�Ax�A��4lF�0;4� �я������_������ۿ;槸��{������/۱	y��]R�T��_��^�J_\"����뭣�~��qP�n�I�[�A���ҭR�C�i]������=�7޿���|>��칟�����g��A��#[�/u�l񖿢a�<ނ���������������J�n������2ݍrv���k�(�4A���ۜ�w9����[N��R�dp�'6�c��/�D'i�?���o����;d�\Q�R8��7J���g�C��G����զ���E����V6nB�� )zoD�nƵ�r9J�h[�¹n���a,U���gG��=�y>�vّ66�<ƿ?�i��_�&�wdBNP�k������`��󋙑����HG�I1��3�T��Mz�$~<�7�f��F
��ŧ���B��"[&7���:&��OgYH3������k�`�Yn<]�e2�֧x�a�y|��+�kg��U�iey��s|���'�A���3�6<��]�8������%IeU�*�1���I���I��"��{���K��F�݀s����36�h^��
�rS��	Q0 ���IKx�s'��_?���Ў���-���<���G6����l��<��{ qa��c��K�F��K�y	7�s�D?TQ˥;"��ׅ�i�]�ӫ�U�k]��������0�Aq+
���擙��O���#������l3[�)EN�G��!Q_<���\8ze��J/>�GR.X�-�{+� |P����U���4�y���R�]���S��R�yͽ��	�C���X'|^>���A(d����m��ǥ��rt��'LqC�������LwF�*3-�}q�n�r�Cs��V��/N5�
�J�v0t���]��>�T0X8��j{����աF�9Rjq����F�{�ڀ���Df��:-e.���%�ɑX�.�X�n�ت�=��\�k�{�U? �Hd<$�7,z5|z-$��|������)	��;;�	��=?]�!p-��ć�ۂe:^��y�O�G�&��֖fo3�w�(�A��'�V�j�Q�1w��� ӆR���c� �Y ���fuW���rI����C%�ԗ�x�1��v���_A���r)��}��{��C5)}�0�MG3�K�E����CiB���
��,K��{����Rf�:��B��v��}�#	���AC���U����K�{��6O�;�V���8��Y� �B{�Kg /�ˡ�YA�yv��d�rb����j�����C�@����+���8�[GM����*���ww����B?����Y˪e����í�Tc���m��0��#�S}�������3����8?� ��Y2��Lp"t�Qa�8ӊG9��U-;$���VlCV���;�Yc��"�PK�ܖERg�
;:"�+��ܻcJ��U�������n��*��ӆ����a����x���_BH?_#+i��&y��
m7�F&��������8owV_���]�s���h�zd9�c9P�#�M��̽_:/p?o����	ؗ7���Գ����Q���`����,l֍s(W4�^�;�`�'������O�/��ȋ�*{���3��*ݭ������31F5{up�1�|��ͳe.e�d�	M�K�z��Ii\YW'*zם�I�n�]�ɣ��Ěw��n�B�1��Uv��+�?�����>}Jul�z�W繞\�vk�UK�)R�/�g,� ƫ=4��Q��[��?��_fZ[���]�|��%��۳��v�ݟ1��/Ց8�����b_nb��~CD��ɤb���F�a��q ���@�y�I<څB�q��?]o@'&��!�-?��'��i����_0���y����"FI�̶�a�k��߂>h<���MTf����%4cZpL�la ��~����6��>�b�RWWϣ�K��gΩ��*����^?���Xx��?�e[#���ǱF�"�x(�=�������˾��K9����޿��AT>�i|W��A�$v��F���,>W����p��O��?�5���(5L>E!ZQJ]����U*��@��¡n5�.�4�����TY~7N�f�a����=,&�`f;P��84���hky�p�H�ÝX����,��HU���3��ڗ`�KA*f�gz��!U�`55���䴍���ư�	,bH��+]����������Kq��)3�?h�yp|~�D�e�M����ft�
��l������M��E�R���4ÿ&��Hg�q�־
�D�[��y[O���e�n)�T�x�w�-��	�,���1����d��N�C�o���R~V�x����9��	���,��u^����+�am�P���[��R���H��S�N�g`ʛ�;~��<L}�v��dm�O��
q�kO{��=h�uf��+7��7s���O�wָZR�0cf�R.�;,�E�j/�f�s�3sYn>>sAG1[6��ސA�o�H*D�rh�J����WUg�����b���h$�O�T�V��gㄳϜkV o�j�+1Xc��z�~X�-���گ��Z�]�lG��<�8Im�����&�y��!���0$�Vh�����6H�޹��K1U��L`���T�n��+�6��(��U,��]y��I�wq�\XT$#��{G�Ր����P�K�b��M㓖z<ܦ��7�Xo2�ƈ�;����7��(�@G���n����F��&�����ͣ�;��օ4����P��r�-F�gn`E���8���U�WH�A��j)�h��qh��N��\��]��3���89r�O�G�f����ru��V�7oh"-�>x�t&�9�p<@uX�_�_���?tIm��{R~M���?g�!׵=
�,\�oz��U����w�����?$Ы120�u���Ih����]��O��@�q�NJ�CxcT�9������G`(`�+*653��8�Y�&o`)M+�
l�>������ֵ$��D�Q~��Z��d��ĉ韶f~X�V��Sǖ��Ȧ�5�q�lq�P�P����%v����H�w�+
L����K_�+v+0���d����Y���T�d��~���I;�\������u�8:.Dt�K���+�^�u]�g�F�o���� ��|����xu������`c�M���{�T),ɪO�������/F�V���j*��<F=���<��?�Jbό�y���ά]��ak٩m)�/���ջ�b��#���
Lq9�CC*�$V�|v��Y�MIf��[ap��Ds�9yΎ��N�F���ݳo�u|���w�v��]_w	P��7�l���Ji��S�31������w%n�q���GT�����)����J3]Q����gp��k�z:����wn)�9Қ����dr`�/+}#� ������y��ow�H��r��Px�)�����M_�3��
�;T�����R�i���t����b4�Tpm��wT��1��f��,�3���f�'�a]e�c��Fm5;�?�p�=�<�ݍ�����*�k�=(;ﾹ?���1�!b������j6�S��f�f�E2�k%c�[;��7]8�f�z��v��r������xg+[ �`���,���0���.'2C��u�iUm"G���'{+�G,�K|o��'�њƇ;O�B�*���^��.�K�16&�"J�����z`4��I:j�����B����+��ϥ���T��\䧲R���J>�]Kg���jL��c�a T�k���jq���m�!�!k
��`VB�t������}��WSm˧F}wn�W�JE>��D-��琇��C��Q�M��*�{���gN�o����q$��X�Ͷ�}D<	�L�g_up*m�tsٙIk��Ɲ�R ��D�Oj��}y��g���ڍ��rM�}���Ff~*�^M}��f ��͜'��fl��f��/��$ƭ�r3���z�9L�W�7U�IN�S^��6�A�XRv���n�4��[T�VCs�M��P�:�$rM�;�Qa:Y�i���%���s�����Z�hѧMwW�^�{7ؒ��j�����-�R�����?W�+s������5;q����[�{aV���PZpҼs%��[L܅**�Y���9q�y<���/�d"-	�����O.���	����xm�Ot�w�)#�и
�F����W�SK~v<Ý���I����s����~'�4� ׼��ϋ���;����-}�x�"�$u>I<��d,{��C��-��%�ܤ�\l��%?MD�׊Q��B��Q�t����Χ_�#�=Mk�vrC���g��\O�3��#K�������;����U/R�m���=�a�L<���1|_�H����{���)�c���fr5�e������'�=%N�~�_? U^��S�8\� �km&m��,V��x��)Ԕ^H�x)W�����;n����v];�<���L'�M����'h��~%�!��͹�~��Ԫ��y'Z���y�*��M�M�������h���VT�RQ�f$�T�~ˬ��w�����VQ����x��5`3������|H���V5�yhѮ_�>�|O[r���5%M��g����r�M)����IE<$���8-��Q�˘p'��}��-�7�SM,�(���,J��A����4���|	�i6)��5 ��\��+.v7���x`����@����SZ�w�i��.;��%������u�n���[���?��R��#��Ĭ�8cӰ�t����2-�"�.aQ�V��Җ�Ѷ��׽3�T��y/��c�V�y��{�L��f������ZX�/���`�4�и�x0�fKJ(�<'�Pc�A�3���6���/T{���u�����_��*1�r�f�/�?4������S��^��Y|���ֽ�Z3�駍R��������S���~�����t贁����?�'��x�����IQn��$�s˸g똜�`j_�iP�j�������?7Tu��\�y9����4Ī{�x�3�߾F�����[DYf5��ҺŁ~�\����P����t[�����7yTSiq$���(����?zR��Ս-��:��ђ���+��E}�˰�	[+�6k���n�fKg!�y|�U0�z}�����g����=�N��UmsL�w8����<|����܈��Cǖ+�i��W,|Sy?R��!�7�bZMv�|�׏Q^?���b^�D(<�6�a��nFKx��/�H�͵iryX�:*��G wu₍q�a�~����\��3	`���hr��Z������ƺ��[{c�z���V�0�W.���p��fRi�4~�#R?��zhĳ3��n#�6����[���Q��U��n�$���JK��@BY���0i�2ZX�.Iq�L��� Fw'ݯA�I��xZa����S��yvEE��=���K�	����%/-�Ss���R�;BTC	d��l�+�U�7���C�cuӜ_�Ϙ��c}���r��+���k���a=PxT�|��a	O���Փr�:��cs0u�&�Bס��~䄟������k���T�̫�n�̇r��ڒX,w~���yj������H�
�No���M2�����{s聅�#`�Jsx$ߚ��{��Я��/[����]��;s*��p�[�v@���ǎ05%֦�q�i%]<~x���߳E)�2�L�O�TMW���D�J��^0��J�����l�+�M�]:�,(*Z�§� CM��qo,���E_%8��N��֦w�U�M�g��s��4u��K+�����wo������f�$4A�94l�����N}�
��fn6ƅ�\�2:QV0�}���Xb�6�}�ɪ�9S�3�?b���^��JS���k���ORs�?Z~�[�s��1�C��*+I_7�	wn�Z7�	�bMZM��y�z�����!�z�,�v��|1��45�Ā��P�ˆ��9�n�Kq���񝥼ü���55/3s��f	�~����X$��?�Z��c0tZ$܇�(�'�UUF�%�I���v�\��9�H������I���Ҩ?�W=�8���r3���2� vq�!.^|yCFޭ]x=n9h>8�5���#dk�\�&wfKڮH�j
�ZzW�#�.&�=$Q��m�����cѪ5�^�:S�Ʒ���ݛ�]��[_1^�n,z���_�L�w�	�D�����~�LMI�Y��2�N�sn1�92WY���h�̔�
���S�
����p���UUcqQ�҂���&���ɪ���9l�����P�s� ��_�j>�����8D͉X-���c�f>��Z-�Ч����G�١�)����Zy��E�f��!��>A\q��4Yp!����r{z°�-��[�P�q=�N�d��i�$��^��p�B��Q��D'XY��8G&|9���{��n��f�M�P��;���k,�\��j(G����<n��G�;m���ld��`�lzo,�Z������$��a���j�qu�������l��}ޑށ��Cφ�~~��x�:U�^�=���C> fO�p��@?\H�/��K�;���T���5��,��V�V_���s��ijv	��ı�y�˷2�V�9���ē�4YR��r�& qd�U-�X񼑠��b�Fi胧�|%��@�������s-���y`�v��}��,��.��݁*`�$�Ph��~2�դ`H�'I���!Y�Z�/B��?���$�P����>��\ʽ̸O@��O���[UX�q��@x�1r�Ou�Wc���4:z��l�ăK�[�9Fq�&([���������֫*��|�7��~� �U�8�դE��\���i%_2^3�(�m��߷�8K�XI�O�����ݤ�z�N(`_�e}c"b�o��7�o���,�
?߫��1�+�^`��b�	9�M��F7��M�'v�^6A�=ʿ.�b%����>j�5�>�蚆gx:$5t�$���U���(@��?�n�~�t�\;Q4HK�lev��E��i��f��87�->)Gz�J�M\��������mO�@��mSk��`4���յ��l��/D��8��p`����z. �7�ʫ(p���}��݈���W���޻����&-�r .�q?$�;Z�>	�~9�jF�.s��[ӕё�޿:���//r�=	��pO��`8{�r|�ZnΧ�xc����'��ػ��1ڪ���n\	��
W����	��Gtp��`�o�",,[�����Bm�5W#�N��HNӓ�F���K@��F<�N��x뮒lK��]��0��OQ�����a4e�2�� Yc�/�;�{�?J����pY���3)C�����9��S�Knf���<@U���Z]t������;J2^'qR���*b	U�|���A���d����ӭ�쳵D!�!{iN��G��Ib�.V�r{� ɳ�S(j�=p���s��י����+�}�(�C�ʨ��Q��9�Mϋ�s�����&�]��f�F����n�8y�s���;���9���[�y#_����˦w�83���Y�Hj�����HU9���Q�)�����(��X�u?���5��1N�>�y������I����9�T��9�j�[q�n�iI�'X���aS��I�@ف�*ǕW�2Z���JΠ���ݲn�t7����M�O�%�w���U���5f^;V��3>2��!���A�9,�u�v�\�q��F��Q�V�ҷ����6�Q�5|F�Pv@��3�i�Ⲏ%z�2Y]2��F�͒?%hB[�1��	�̟�/(���oɺ��+<w(.)�|��|��V�����G\+&d�p
qh+����������a�s�b��.8�m7����aX�<�r}9$�j��ŴE��b��G�|�b���e�=�H�C�3������%|z7�so����� �d�Sޗck�g��S���%�Jn̴`6{㘏dD��+��^m�g�����Q\��x�Dў�oK5����]-���jX��	->�y�Z��2��ƹ��\!��P �'�*��]�����*��f�_��)}�~���ߙO��&U'd5ELązO$f\�	��ʭt�³��]����o��#�z�n6N'������o�H(P����.�wUqm�4Y
����#�־O�p)�������L�sGl� �&���$w~�;�Ζ��gE3��I����.�=����q�0���4��%��UE��6�j��Rh%�q���2�c���D��P�(��Q�n�K�g�D��S�B�z&���Q��/5Q���ۋ[J�v=;9Wa�9�����Xn�*&+�֯�O�٫��b�ۤ�ȕJ�Q��X���;�LxQd�7Ђhs5��my��r4�C��̳�pwDS���ì�)����I�s��u�d.�ܰ�͟�{!W�A�U���^����e1�	/���#F�֨�)Q�i��G�6�8�1�9Vcj�]u���>{QTl{^'������J�9/��d�I� %#�Vw�܍���JU�V�B�ew�Z��c��<�+f��p%dLz���j��ar{�-�]��ofK-o��Sl�lܢt�d�45���/�O�W�O~�G~�}}��	���jx�R�q�]���|�
���ei!����N�߭M����d��@c����v���>r���b��~\��-��A]_���F� ���o�euA�i�J���
T0>ُ�D�~�ևO��_/g,�~!�V�0=iL"�iG�>��F�	�L��g�#4k�biDb�xn�g�!.ӡ]&�5Qa����2��K+�WSm?Gl�����&@�3a�� 嘶:ljwTZfqf�bJ��ܱՒڿ��5G�\�ٱbp�H��G���ˎ����K����MJMU��b�0+n�Ԡ��wM�4t�5����Ծ��X�7a��aLt;������>9���V�#,�!�A��8a�rqJT^�|49.ͅkeaw�X0.$-��-W�m]�X||�ւ!I���?p)��j�_}��}��M�Ms����K1o����n,�Ed�j�}`T[�Yg��\��Q|����NL�N�o����[6�gʫq���Gu"��U��(.��ʜ!L�zC��u��vx�uڲ��X��u¦�����6rӬ��� ��}�?���D�V!!)\�/�I���Q�zZ�K��I
��_�9���&ǟL@�x~�O�����T"�W�]I�c�zW�Z��P��������їT����-h]+���T/L?|+LM��AW�GسW�o�����Hc�Y�ʞ����a�|�</��ۧ�50²�(o�����u�dk,�#[C!������ `�S�Q�g1�U�&�6­;��O�k�C_&����Do���"���-��a�ːx.��v���o���hhwq�d妾�g��T���7.��Aܥ�<���k��k�㩨��puRӘ4��Y�#ɸz��ʃ.�Rr�R���������d���$��'U>;j[|9��J����dP5����i/|�OF���)�=� ���K��X��[���2H�;}0���W �>��4�G�Y��Wf.Qذ���M�r��٭�8^1(����;�Q>�֑~z�] ��v�qW�}�`�Z_-���Z7c�����P?��mFP�Y���xΒ����]s8b���3S�E�s�x�F�Bt[Hu�nF�W���q���"�1�ހ.��	�׮I�6�wn{��8�ޱ9�(�;�
�g���B|n�H��x�3T�,RWk�v�	�i�����?;��N:����*���	B-^�&j����<3@œ����'�<ͧ��}j��!M�7�r�:��D��j�2�n�?[ĝ'_��8��h9Wdr6�lj�-ݺg�L����F��)턲R����
7����?�m݇Bk��05�1rԡ}�	C�
���t��È�k��L��(���Ro4��&!&�8V+�:N��a��#$]��9�v��>��/�����(���c��u�?�Ӷ�ڤ�|�jb�>tE��'G���}1ۚ�i=A���2����MM�{Q"���M��b�˥�kDO�tʣQ�Ζޡ���Q��䍍r²�z�ګSӸ]�j�����CA0��
����x���S�?j�=k7��<��V�	��Liu�*�V��*
�]�g��O$)%%��.�s(��ݓAH��]0�$�>PR�$�������=:��������"�޶�[s8�G���Z�RU�IS�8��7�F��8�2�̬U�;K�9x�L����`�18�Ly���~ΐfr܊�[oݿ\����I���1Ae�����?�<���}�ё[�q���>��E���wkZ�9{�������S��P�L�B�y���Qֲ�=�FG�犅c9Q.�i���d����κ�MI����%j}8)��q�C��6֕?g)�G6�O�zg�ȗ�XN�MC<����b��L�d5���Ё�+��_�#�YokV�w��[\2���U(�fKcJ���G�n�Oo�P�6��
�QS�\0��Q��Ŗ8Z'f)�̡���>w��@'����S:�՝���C�l_�C�u[�8�sj,<뼲t��@���"�jio	��$Lv����uX_�X܉��<w`�X�򿏃�o�(jhP��M_u�����?�s4�f�`����\�$�P���W�[��֮�T���((�`+�e��r�3H��,�6�6iZ���ěU#cb�s��,[`Q���k�Hk^�8���ͥ"Jٟ,D�r�՚'@�Pl��8io.z�ѵ!%���$4��/�/��]���������,��`�s�.��L�[[��	�o���=0���dƻ��S�1�1�r(*z�J����qJ�B��ʷUD	��Yӟ��G�d�� רy{pv�r%I_߰�DaQQ�4����
Ԑ171˦�y����>'��CQ�T?����P?��[-���ݞ�J׉�n3�N?ޚ���X���ܸ$_�Q��61v���k,�ݚ�ӂ��x����k�#��o`S����g� xG�����b5���O5�Ʒ4��9N�rRb���nJ�\M�O���늑��5ϲ�ػ����� $M~b�*QN-�����\x��64,��Z����ݥ	�#�y�]��v�>�k� ���ΰ��3�v4/�L�g�=CƵ�h���D�H����N�x+F�-�2&��%O�c�ʅ���s��c��ZQ�{_
����z�e��}�ݗ8r�=9�:��4���ϧ�ͳ���m��t���5?��)�Hk���|N�>r|���!��,�]A���<Ә���ᚤB;OP��>����m���'�.���m�8�EY�$ޫ�^f�y�#[��u��\��S������&Q����f}��U�\��&��ʭI3]�f��(�j@�L�I�U��WP���)�C��P%J���QI��\] �ã�"��N	��m�G�dX���׎6tJ���PpUC3�?E��Wf�����7?��i?U�i�|�z^~���(���n<_���>J��5�w�.i� ���d����G1G3�!FK�H�a�6�>7���pA�DvY'wb�G���_�Wc���##,
�?�D��7 �H�'��i�p7@y�K���"{�`R�ؕ[@o�Ժ�̦��+�8�!��R&ܞ��~k,XZ=ן�F�+������z9���n��T��/ۙ��ԙ�!a�ݵ��)|��a��hAv�����Y��N�;|�;�A�!����0%��sё�Gh�/�����R�7�Ҍ��ԉy~��v6u*���X�^��8������M�y��`d�p�;��&Y2�&�S�z���%�[�~w��x����ܩSuL��7��*�����!�@�wX���Ӳ�!#�~�Dʻ��ɀCTxJ�VS�3���pa��c9�2����n�l� TUQ�RE�o�.��(Y���G.}�?�<?�ɜw�����%��q0�8��ѯ��G�ڷ؃�$�r�=ޚ)X1��?��ϭ`�gX�}�V��D�����yf��-3�\�e),��c�|��~��;���J3�yMS���4�@��&�*���"}��辟�+���2	3D���p:{!o}�-TT�p��$�45���iş|�qذ�3�.s���V���[2��tzj�T���S�v�)2���A�mPc���@�չ�\Uޮ3�ey ��� eŕ�L�yJ;���Ӽʃ=w��7�s�+�¯�R�T#��&����b�n��4��,x�H�w<�n0a҈q��ֹ��(+��w���u'�T��o?�V�9K*� �r I"��(�F��4?��m����9��׮A �U]=g���$�3��H2���뤢4���#�[����`X��}t���B���\�H�#��m'>��ǭ� �B��/������#��Z��MU�e�D��_��^�,妋�X��n�H3G��<��H+�]�oU��DQ,24K��� 3�}E
��R�������L��uxز��,�:�c_��&��u�`f�;�w>�TH��4�	������:�d�~f�,<U�Y.���A�l�k�[��m�����+�9�#z^F`�OJ�:E�nf+}�G�����Pe=;��|��6�Ճ�.jf�A�XSf��'ce�Y�Nе�.�龱��$��\:)&i��Ӽ ��#�ӧ������Yr;l@�kzz�+�σ\�W�x�j�� �V�S�vs�8�z��y�d�#;����54����Q#�.�Q�)����߷L�L��m��!�(��\'S�Z;��5Q�y�4 �3e�H��u9����"�2v.���4⃟��zaʔ.�O\!��0�֫]�rL�6(�~i�Q���\�P���20̰����J�|��즺jc֕۞�{�AR��G�ϖ��9���s�wU���ۃ���-"�턀���"��m����'�JӋ�C�s*��{�^�<�f �����6:|��Fl���k���Q�!��K�]q�7�ub�a֬��4��|0b3>�fb]xd�l���fP���d}�H��T��`�!1��h�0%~lp�)�F��m���G�̮qE�����\�h�tbK&��ZP-������zǞp�r�?����5~��I�$���r[�[ǘ���Y���GV&儢:d��XV*��Ǵ�����D����Kf���4Z�z�	*$�?�<Q��uh��d���rЪ��KYy�D��7K���6����ؼ^�{C��}�c0�xY�io=,:X��X�һv��iK�7F4l�]���z�lrf��TG	�뮭������g����8����Ô�ӧ\p����$hms$�I����R�t�]�СI�d�ҽ�� HH������e��b�KQ�Ј[W;��U�ܥ�S��b?���t�j֔�&o��#{�j"�%"h��A�_lR�ΑF�{&{چ<�����1�z��Yw��X�Wex)�X������ov���|�UK#��!�4�:��Q}��L�% Ŝ�.���s�Ŗ|�-)z&�7a&+����X|����怬�G�%β�/��.ƍ$���NI:t�*־:Ww6K��}��\t�X����?�����3�ڿ�����{U�����e���!�,;��T �x���e�]ͬں����s���B�wΌ�צ{��c�t�/'3!�<�E��� и��z�����$c�C�(�D�1�K��~���T�q�jb�0���D�[s��V˙އ���[��8�`���B����j����Vu��:O����t��c5G47�H�f�pp���;�&�>����V��i�բ�@ا��ޕt��" ���K4���V�Gޓמ�?��z�`��k��~��7���]���^�
<���|�_L%)��/���Ε�	w��ps���Pߖ͐�W]���{���<Z�k�16�����\I�A��Ղ�b���G6BN,������K�{#;;���ǰel����j�fA�xi���\�qN5D��������H���L��_N?x8��}�3~����0�>�&���	�}��� ~[o/�����Wm��������
S��T<A��̫ip�U���J2^�V{AfKm�} ԗ�B��'���7�B]R�������L�w-<o�1������I{��+ħ,1�&j�.���pA��a����Z2އ�,�_-'�5W�F5;���U�)g�eNI�Z��՟��|�k
�*P��c��hxO��Bpm"g�����>�jSPS`�W�O2h���|%&��\�Bw��]26�_{w�!�q�B� �0���!E_oΕ}.�9�˝���Ț|ay?Tr�6Ny�_i�R��=[�t�(�Ec�il¶�>��u��� C����B��� ��ϝu|�/�}�c ��X��y�
��U�������+���$'�H�g�7�g��C�&�a׮��*�2�py~ �QM���q��GC��nU�F.�Gg������Kt��/k|mA��4��FDTG�oX����4�3��M��+n2����k�̏?�Ȟ*`������^d}�i���1�v��+��G��8���m�6�CL�)���y|��Ȳ��5���2&^j7ם��)07a"�+˒<l�����`���w�PK'ٱLÖ+eO��)[���US�+�c���b+zA�&��m-]��9��"~�ӗ������vv��"��
�� ��2�1��J?JC��'��(�-�oDC:E�D*$���ʠ�*�r3@��?��Q�>��;�A$]�>�v�mRy��/�`h6z	�_�|Zv}x}�,z6���Y�)�E�lJ��'M���x#��e��,r�|���eg8�v���n�X�����K��5C���{��E�v2�G^#&�_�<�)-�oX���1�+1H��po��(���ti��+Rߡ�D�u$J~��z�P�7��O�Vp��%�M��c\t��>�m���Ԝ6d�Z��ˌy�����_�7γ�c�'D�_QJ�,� M0K5$0��,�L�U��.�z�$�N��3�Ù_�G����^|p�џ�|��;T�C��Y9D�<$qa���h-���{��\-e��)�i��_ݣ�"��N�^^>	��."��4��^�$�-��٣�EE/Y��~V�X�G��1�H=�L���m��9nؼ��F�d�t���X���c!�#A�W�~��xy�������HŶ�u���<�D/7�Z�ф��T4��ę&i϶�~T�
;�4:?���:e��+`�<�WC�!L]o����!!6�m����`Ǆ~
��|��X��]��y�7LBm0E���)@#H��v����Ԙ��S�=k�Ұ�Y�J��j*�E�[�Ó)�+��MkZV^a�-�=��n�����_D�t-���ߑ�ٍ�$;
�`�7���d�/�?��||�4Y?��&$c[I���vwcJ�*挿�}U?c�gF0�<��J)dNC�Zr��_��$�o��R�<���y����[���I69C'_r�M�np8����MDUk�[��d�E���GOܭ��?�6�-��t[��[_?:��� q���,��c�]/���Y�_�:�ƫ������[���6J\�k:x��ᣔ�R�~������"�廚���ڽM��F��A��q�*�����R����6L�B�A���Ɏ����Y��@�3�{�e�:�Ĥ������w��ϵ�&b���CvS�J	�h�f�(F����syy����4y��2�i��'5�
�Eϛ����:������h���ʨ�Q��ԤC$VS�瘾����
[F8C	��"ϻG:��[҈�������^Ɖ�N�V_I8��5_�(:��n������Ě�l�DW[�.�~��m�z����S;4O��t(�(��)��E��e�7���ؽ�ٝWjߢ�$&���:�\�?TTU����ɳ,取p���<;T߽d������3W9i!���8�t>�h���h�Z�����|�� bK�x3�u.��qл��[-x�]JT����AA^�G������A�����!͔
"ª���rO���g�;]���Tۖ��|�x^�k��o��v� �?~��[ڡQ�q+�.T8��8\;��_�P���A<C�a@N�x��0�ĚhUwz(bW?�҉"���i`�񃚎4�`����o'�K,�٘�L��ᒸ��+��@�y���]��7Gz�1��'[S�L`�{���:�G��P�u�҄vt.g-����ʘ��	�����zPdC ��~�0�-�k;z�,�IH�xoٳ��E�Ƞ��ez����b�������G�K���H�*c�ɒ�tk݈A��:�����G�Y�
i�95*Vp�n"@�K-���!�۶�Eڏ\m��ݚ>�v8ZA���<��<�Ѧ�]a��Wӑ\�.��I�m�����n��'W��xH�
�v�<Ү�@PM�S����T��`ʻu$�}�C?^�Ry�b�`�]�;���@�FS��dSn����#�{�).͕���.�p8t�~�[�K�@�������7����ʻv���^�yA j`��W��65��;S��$�1�Kp���2��"����n����a�v�^U��ȱLث<-���y�c���e�V�xΨ;>�h�����șp�uA�w"�&�dJڂ0�S�xi����j��O8.r������]�`��ҁ��G�������v*������>�s�m��,��n���`��8�Ӫ�;!,(�Sd��@�
�F����<W�s&R�1d�`+��n��� ;�����q�QQ_�(�%݈JHw%� )�]1Hw�����-5t	��9t*͐��s��������ݼ��=��O���Ve8�HH)�7s/s��ܨq���{,�]�*�����&'kh�V���3�&RY�6�]|ݣ)�Vh�GXٕ!���6����)I��c-3	��a�,�e!n�!��M�y%8��&����'���)	����7���a��b�������\�/k] �WA�n���O����ក^K��߲�����'�)=��)RfD$���޴��̛�9��u�]cX9sS8�},��;�R��7��Ơuh��Z{0�H���!2{c���z5�����t ei�M�K����mC���0I�=tq���.T�p�H��L�a�B��ke�[���W=4��2�:���70H�pg��bP��ecL�)�l�e&��ܭ�8��8�Ȳ:Z����WT��K�=;�� G������i$�3��W�wu�9=�I��3���=�*U������ ���>TU��3��li��#�+1����?����u�"ת���r��(e�*�{6Ș���d�[��W�WH$��=:i�U0w�İrh���8�ޱ-x�oK��+$'�����E8�֌����P]iXظ>�WjF�>&ænq�ye���U��W�g�|�*ݣ-���� �^�����_yu��6X��Ѻ-������	X��Ǐ������+2x�F�������aYz�滍N\:��/ �眈��J�m�c@^���>� �z�E\�����R�K�A)*2��"j��y]�W�(�����/��K�+�X��3��J�����~�EҚ�7ؽ���g�\���=V�!\�	|�NP��I��CN��_�Í6k�G�ƾdc~4n�ֵ����b�����Ї��`�o�(5�q��ׯ��*�+F_����=V���=>Q�e�Ɋ��Q�Q��6]��Β���y��w���_y��N�(�U�ɔ��m�;p\��1�!��a�b��4��1	g�^Ƅ���������9ù�(��S�Jx&c��"d�G��8_���o�B.�c0Z��,K������t�D]*�K�?���{���P�M;�eİY���5SaM���%M����F��?��~���ށ�8�on(a�M��\��v1�N�CGUe��}�H��Qs�� �NP7�RId h�l~N3vO��Y����q	���M��#x;u�0�
R��:��2ӟS���:ϓʹ��������e$l��t���;b���z�x��;!��pA�7��d����WcE7޿���������"�XO�8��D4c����RW�٤�y�E7��J��!F�u�=�!öQ�n��⚂�. �h�C��H9���G��=?ʇU�.Zl����E�U�N=�Ŕ�z'wy� ���jGR�F!�h�D�etF{�י��Đa�(Ϣ�@��}z��@�:LǦh~X�\�xy;�be�o��觏���80�0�V��J���ڣ�������;�+����h�t��G�h��P8g�|Hhu8�����)?�L�\��9١�;�(���IM�oK��͵�n�lɲ,n�;h�w��� tޒ],����LHh�>m#��u�.ueJ�;���l�A�������@A��C�z��IZ���V�9��
�GkF1)�,,�"3>>�1@�?2�4�f�k1k�2_���u7עҫ����,nX�����[fpsN���S���3u��8\"s����_I�����c��O������5��c.: (���V�&z���C�Q���R�WIj�(�k�����I.�ޮى	u�8��d�><a����<T��g�Ϯ\��;��%�k�ʶ��=D�i��2J�����eK1udB1�`)�n��4U�2�ۗ�G�$3�Y]A��Ÿ�^l=y�i��E��UtȲ�� Th���V*����8��Q����1F���kC\�G�5o$�oQ�W�m���S<��~B�85�|e�B>��?D��N̬u $|�v�G萇�^��l��gc��J���d��ҡ��W������ٕ�E���n���[����ã�R��b��o"oB������WZZ��Ŧz����}�]=���[���j�Ƥ��� ��<����]%-~�ܥ#�G�u.*��q�uT�:#�_���cc1�Y|���4e�g������Sa���43�R�/��Rn�c0�K����˝�lwPkc"J\{p��uFx��Y��]���e+Z͸-�ؔ 	�4�	ƭD�b������[	a+�wd�n�]�$hX��e��f�SS�_u}?J'�@���u��v�h��T���<a0mеĵ]f�H��V���'����\ߙ��4U�_i�sCG{�B��w��N/kT؞u#\Qd�?9��UJE�W�_&x��:����zYm���P�'��n��	u������09��E�5��铎��[}�������V��Y�����8�]�_�0wv�R�v��@��EE{��z��k��x+�sg|jZ�*6����ᘇ/l�11���G���
yfr����R+�j_�.�|I��g]�3�2<8����g��[,��d��*�uV3!����h���A
L��*�X��u���څ�Ra��=�n|rGQ��(߱ٔ�j��0RC)q�����r(ݏX韫��wT���.�1>GG�9�AxIW/�[�D���� /�z%&BJ�����;�`��_��
0��l�]�s�N�(Y,U��4�,�ι�t��[{a�д��[�����!���)�C����\S�~��@:�i� q��vk��}����di��y�5)��X��k��:Wmċ�Ӟ����������-[Phi��+�eb�7h|����t�L]����N��T�$�۪�-����Б!�2��Di�O��I�Sl�ޢ�W�������ՊӬC�ɂ�L�Y
k"�/�DA���_�L�p��#���&��|�Z&/���q�1D
t/�d4�A<]ƣ_��+ܧ��J��m,���ђ�-}(B��"��\#�z�~���3�������ڮ��륍ol7���'u����1���ֺ�J�Su���, ���>�� ���dĘ�7=��a�޸���5ʮl���*�G���.�6�ő�fҰ�{�����>���qK�� o��@zko�~�v(wCh�v�f�u
l ��Z�k9s�6���3*}�s!�X�� ����Tݕ%t�LTUO�lpc�#���mZ^�,[�k�����vQ/E�8�o�� h1�1�O�g��[�}]Y|'�&��_���D���u�PT��y�0�)�c�2Ԋj��m�^��!sGi�Ǚ�^�Q�k��Q�Q�����(��rI�o���>'�?n��=���-z���gn�% �&����K�	���	�7(|�`<�GcRȝ����#(~�hFS�ʇbj�x�Bd�k=p=�ʩ�=k�i�ca��Gi���_�����jM�[m��b�)y��F:͎�����﯉KwM\y�i�L��h�;<cs���F����t���,daV!�<k�jC�_��n!��0Ӗ/I���ݘC��W�\
M���]e)��cY��-0,O�xw��X"�m��Ξtk��9�}8�k�u�B2>��y�s2e��e����К�p�?�(�.) �[�"��V(�r�C�;с���+Gw�b�f��o�@I�����P�H!�B��Lst�o:�,O�=�mk���jx#����U�����]=�V�u�g�WF��[vN�{^ɊL'�W��.�H/�]|r&���3����AK[�o!Ww}m|گ5�t�T�`��PT�0gU�H'�S��~VM���J6� 3gl�սP��ז�_[��گ�:%��mG�pP�5,0	Iȧ���f���$���>1�m-�a��)	��4�;���'	��.f�Ɔܞ����Z�#���V��i\�;zyy��o)ڳC�T��p�6�>ǐ��d���L�Ѣ�J��*�$�Mٛ�MY)�]����r{a�B��}���P�V≔�1c�c�{��;���n�ˣ���s�^���j�<�T�������Q}��4 ��*�m_�ǹ�5_�����M� �4٭�'/Kt�.�3�X	�r�U�{�z�w�R�z_S4]E�=hn�����f�i��h��ʈ������������}�ٸ)�C��F9ҴD;�F}|s�c3���g�������ق:gz�v����fQ�7 +s��~���{(���xX�+d4�v����cH�&6����1�1O�f$�$Ԛ:�����˜�D�u��o���z���m��5o}�f�C:�^�a�� �=���XTN�~	�Whe>XS8� �7��,N�юۚ;��|֏IJ�2N�b��,8�~Mֳ�+��Z��b3��Y�Qg�E�w���G���?��<���.�n�6[�R*��`٫�dV�8�H�//�T!�"t5�>^��8�Ԁ���m���
�����7�+���w����͚���S�p�E��Ҵ�@#XYI�b0�ã͢���}����jw
ٙ��?���2�3z!(-�q�t�Z)��M	DB(#���܁�ԃu�c��[�{��tB]��wAނ3s^2j4#^S�qB~W?`���9�5��� �3G��������;,�-UK�9�����Z�ͅ�%!� ��E����~���Ͳ.V-;��ҩ�X���۞U�K�KҘ�_:xZ;u֎Na�c��0��'A��VW�@�0AF1��q�{�h��
�������׶�[��s�g>F�?r�8l>p�Fr�	�r!�n��/k�bw|_k����*�QV�P�
]��0��$�K�t�� ��w��-�Ks���ɪa~�g�u�P���:Af�7��f��'����������uQNV��_
G7��$4��%n���y&,�ܚ'�ICNrP���+<��'���=tH	z��j9)�{�O����e)�u�j��Nz+mxLҹ���@���ر�C�W���I��%��|��g���l�Wz������+zN�[�a%�J~��č�a�D�,��<B���������)^\���RC>�K���%c��S�z�Q��c@H����� t��� ���M���# ���������DW��Ѵַ���:wt��E��m����3Z�.����G6�^��~�<��e����r�6�<o+'%G�<5t.E5Y�������g���Ȅ׾x�j�@����]�����Ł>�=i�ũ�ܼ~�=V�(R����UM�B��2������&��N�ß�Ph�����V�&�>�>��W��gt'҅��C|���
���1���&/�P��Z���НI����l2B�N��{��b����@�Yr9~�]>�)������?�^��l�/.]�*���e;�e8���ke��|Y��nf�3���i�T�K�m5����&���Uʶ��W�1:��E��-u�FM������]��~�
��fO{_��S��t;ܞic-��T�G�$F�%�i�54�JWY9:��~u>�+�	����h���aBE8����0	�ġ��.��4*{��I�3)�:���\mc�8�$�T\��S��SY�Ni����Y������=�|�ڞ�	�D)+���ߙ/�9v�O�Df���j�Wv�4§̷c�d�,^S1ݤ�~�`m�W��iWg:k���S����b�.��$E_��;U���Mc@O9��
�*3�\�s�gL����R�mPI��
.�'�VP㹘������j�m����;t��������ʶ*�7��3S�쿝̽��4<��������00�z�uw��Ĭ|�/�,�o�(���:+)�&�νH�u��Xb�W�ok���r@�t�����!-�`/�o��()�wq;̕D���z:����?�h9�+T����j�3�!���RY*�_��m��J�2]2!���}�L�X��Jߟ�9�g	�Jvեb#Z�-6��P�DL; j���[W��Υ�����G��ȵ��Z7�{�O+��e�M�������YVאw�L <z�/^�� �pe@bs�x3�_���xR���}��ܛ�;�Ҷ��vh�$�xg䇭�@0�^��y���>셈�y?�k������s��z=�r�����*.��5�kuZ�gY>0����b,3�h2��,nywW��x�e
TrK���S��8ͱ�:jO��3����ԩ�H��Yq�$�E�vCF^ұ%0�eS ߦ@%����5.2���2ED�{?��#Kh�5���t�oj2-OU"���{aQ�,�cB�+ӹ�7�'�C�Ye��[������}�����&���-g��݋u�'���_�.�z"��T�+�n[�ҧ�Tɣ�#�Um{`���[�� Yه}�P_�e�K�M�e��q���4WZ�ii��b�ɖ��C~���]�9r<��:e�+��
3����R�F� R4�ߙx"jHf��ETi�.kD��E�:��`-7��.���}�rbl�F�yN=��{)ۻ(TL6U�l���j�[�ļ~�)ߕ�8��F�gw�1�=	ΜB �պ���q�G�%��C8{��q�^�G��V�A�%�ϭb����S�f�^�E9)�UKևɇ���Q�����8V���-3ƫ�A�����r��y{��-��S��W�p�MT}lW;�	��һ�"��xOI$:���tq��!����w��X�i4��-o�zef`�:Y�mT�V�kev�jk�\d��O�d�eј�	��Z�5ze���^,�^A\ev,͸w=yL���X��CƠ߇,k�H�(e
K������=̲�d� I�<��#ϸ��?�	,Ӏ�͌n�\c[����H�Ds�ڨf��^�b����F���Z�����r�� ���zK�W���,��	��8�hTT}�Y���I�z;���
	��k�&u����Ĩ��Ʊ{շ��]���*|˥���!֘q��&�����MӋ�.���~2������ĩ��

��̥H�*i�ш����ܐ�e�go���>De�T��|j>:n��$�����E��M
�����9���(��P�w�$�#��jF9r`[|�f)�"���H������nGd���AZd���X���m؇�Y~.m17ܬ�k>�.�PB�sU}.:(�[��s�3@��.;�i��b�W�#�$rh������P-�BW.N�'�4_��C ��Z��U{�Y�ؤ�M(�\ �l&��%��V��Y��	4�сޱY΋���ʧ��3�ɐ����%a�w�ɓXr��q�Ԙ2;�t#���;�d�{�f<L)��@���"`ve���5xk	&E[>Qh)+vHs飭�gYږ#�qg��i�WH�&KC�<�����Z�vN����ߜȌj��9��M�4p;&�W9g��n�����\5�۱f%���`�!i��G����
�L�����I��̤\��lM��Y��H9��z[!߰�o���K0H2P+M{��A���Q��\ߘ��($���r�!�+0Z�;ʭpw�S!�Oq:��2pSe��#��j_��.�odF��x���X�ZD���t���W�(HeD�|ޛ��̉1���&�l��L��ʸ���	\;�X�d��ĵ�_=ު�c7)1�.�?t0��.V�P�X�O��n/,(�����n]p�K�Z1a���V���ǭ�����Yp���T����b����}[��C��!�p����m�ml�za���׸���Ix�|�+8HvZ�{�q͘�
C�w�h.�t�[���f\�9`���.˶���r�D'��9�5�Yn�8�{���;"w^���-�O��='�?a��;\ڥ�Jo����#Z�>���p5�����jG��53��P�գ�"�6�po�N�h���6_��]Ƃ]����!2֜N}m�ﱜJ����zy4��g�\�;�����Le���/�����M<K��L�:4���>��o,?3۪�/��5��4߇�U a��'X5e�g޹�"���IET�ÛdQ'����J_����ir� ?�fX�wE)��cc�7H�f�CI�7sXZ��c���)����Ne������$��#�l.��f�趫�!��?���7�H�� ��F����>.�^���TI�"����3nh�M� +5Qu=��o�7v��b��n�\�N�8��>��^�$������:8<���yZ0�U`��P���[�`~/²�{��&춅�q��][�\ ���42�u2�=����)�>������J팗ĵ�٫�¿�B!w KL/��*������i/�{��l��K�~Ԅݹt���K�v�6ag��}B��Uݣ1!u`���/G>������!��⠡��2� �&�	8�;8�gf-?��!2�G��A���)��yk�-1�5��pR+Wg=ic��;D/�ܑ������1>ӍG�
$0��oU���5�E��6�Ƃҽ�k���x�g�����I@�3t$�K^�����F`��/]�6YҕQ��,��*�+Q��Z�\;/?���ޓ�%��V��$�7E��f�U�w�~�eM�(!���f)����h��v3k��;�"���VI9:ֈz'��'�ft�L=X�� �G��G1j�KH��k�'�"�\L�QEyw��YӍ�h��'h���e��o����?��N�4~�|�F}2��v�kGl��hs�	���d:�&ŮfA!|�%F�S�� 	m�x����z��ɑʠ9���_ȼ�[�:���/��{CL��z-�M`��QE����k{�E��o��X�:L�O�9vYz�7?��h�yř*e�W��G&�7b�QN;;�ؘ��)��}�������� V�-�����F�G��R���n���Mf�0D��6�K�����(�}��'gm�&�[�6Uѳ���&����q=��{!�QR{>d���y��PT�}#�T�����oZvJ>�+����݃�9���Od���'�f�w1��L|/�Ȝ�:�ùFO���J։yYa^��o�3�_i[[�E��ڽE�/�J��G�Ji�+xmKu��GC�z�9�H�Zy>��"N�N�mQ�fmm�6N�V�i�I�u�zi�Ǉ��3��(��/&v0^��gŎU8=�����>�B�م�	'�x>�_���?���}-;���N����hQ��yެW�3�ֹF zX��h��M�?�ħ�%l��ڡ��-#b��^%��U��Ws|�=�)�^���S�����8�85�\��O�Usj*#9o}��H����kX7Eo�}GW�x�l�˝)������h��������l��}xg��z���9���QyAĥ��	~�7���߭�O��N�W���5q%��|��u�n"�/K�
�ok�:��|�u�m���2���� D��Ϥ��6M��jh��/�<P%����^9�+��t�����e��۝oz� o�R�TI;����a-9j�6SƽX� YpЮ`���5����-HQ�5��
���Ta�n����b�mLwky�UR7(o�V��;�����r���j��ܘ��{���\��mGR
t� y9����~�p���ۄ����vU��w��蕮B�ݼ�ձ�7�W���,��.��.���Rq������]dĮ�A0\n�Z^v�/��#�sÿ���[+�p�U��܁�\^�AIy�E �!D�W/C����k�:h��vI2,�W�S�f��7[֠�i)�5]p����j���H���$2��z�)*6�;��}�^q�Y�5�;200U����7v������w�������X�����h�%���\3>�V���j��{}MOvu�d�2�/M1�[T�/e���L�NO�������Բ�8���Fvc�s*�Ɗ�y;���[}�j��:��6>�U�I^!� �C��m<�r��YP���>Te��3|$A�U;�~Cx����
����Á��KA"��1j�0 -�{މ�����mϤ��O�=�1�Y�������eb~�f��#�B� ?�w���'���*TF�r~I�-�s.�+��z�A�3����u,/W�����'�k�-z�"�;ԡi�e ���)�ѡ�US�t��-H2�B�r� �*��?��4U�x�h�i���bΜO��&X��m	�� v���H�yTq���^_t�'���5)�M�6��۝�B"MU�	�[�z�O#�?�@�{�`6W9������o��涊��|$�����)Yl�r�W:lu���u��Ŧ��nG6�:ӎw�-�d{[V�n�#Y"�40��ȸ�.��c��^"(��<=j_�d��=�).����a,ޫ��n�@���.T�\���&�ˠ�B�*�yTV̓�Tl�D�����wY��4�kb㋞o|��?ā~�	9�f�E��BR�&Ŕ���4z�,�26���7�����Dff'BG�صg;�BF�7dY5���A;�?����#�'���6�}��o��%�Us��i}ңɌ�v�"�\�yĊ�x.��YN n����2�U6M�d������9I�.Zf�>ri!�4��uD�3C���L�F���fL2q"t^�{��1��+��Y�&�+�;���I�wv��4T{e�F�Fb-��L;�~D;�y���-��񂊿`˺z�E���q��2뛶��ǖ�3��WD?���[l�{��v�B��+��1�ʒO��_\
պ�a�1�7x���T���^}��x�̂:��)�����'�&*�M�Ҍ_�Z�I�ʦM�Vlz0г��� jC���@��OP �4@��j&>!7�R3�ݭ��	�jd���Fy�Hh	�]�
$���E�)���$����(�_ǝf��a�
r-;������2ݚ�.��)�0�ޮ~+�i�j����&�����v��PhgVY��{�љۍ`�Mx�'dD�.1�����$(0���k���#��J�L��u��:�Mu{(i�3�b�/q!B1l!�bpF��u*/�1i��p����FT�|�+3�z���0����.����萴�aK��\���ʹ�f����$���
�w����b��+G_E9�⒠*�C1sϜFF�odۛ�������*��ʾ4~�<+%?�5��l/B��͍�*��sd�X٤F�����*�R^���$��~Kj@��qQLB�Qa���P��6y[�b�ܒf*�c�+^L���oh��ô�k����02�tdB�$ љa^ �rz�ge�~h{X���A���� ��9wM�Wʣ�`�}+��wѩ5�E�L�_���X�V#J(7t����>,��E�3k�DE��y�\+�]�y@Wd^��]Q�"|�4R�^S��D??��_=H�#A�,����i�95L���<5߬/JG�H굿�K����́Bj�`���R�h�V�X�t�kd�'�u�L*seqg�I�r#X8+]���B��&�t�ʋ��.4���& ���=�9��L�sά���a}5���H��mӴz��N,p����[���WA5ۃvYQz)��3a���C�l����f�j��ERtp��*���b�g3�w�m�4�U�OTş�rt���,}R$�?�ՍjP��4"s��j�(FWJ��7�q����~3q��(&��ɬ��J=�0Qd��;��@�F�֋����G������F�e�^_? &܇��[.����Ƭjd^b;��yֲyAQQ�m�t��i�3TE��99�s�
�v�޽x�6��ghѺ��l����ر�,�D��!91��؛��K|��jRH���N��.*��uċ�8�������z���ͮ՞�|y��� 8]	����O�Qv3��V�3���Wh����0x�3�7;;��(Ӌ�ӛ�§��b�$w�[����O���\6���=o���_�=��?Fj��j�f5\5X-9k��Y� s����{��ٚ�����k�i�w�+[�s(�Z5��T�:�W��sc{
4t�6V�bp:Ҿ�U�f2���Zs��z�G��4te����6[�w����=��-��&�)��_���-L�_iR�(0wM��s��;2���o��垿y+#�g�eU���~�I�����zF�.V��~"�㫠��WnK�`�s���n��a"��'Q]�-��Y�Ih����W�$�b�N!����<�B�����$E?�)����,E��(:��xGW�G-��@�]?�%�S�FУ+=�Cb�aBts�! ۤث5?c���*���ڊ׹��`j���҈2��QU��̣�3����26��u�z4��`���ǩ�	]�����d��и�~������SF ����������F)X��/��[qc>H8�WYO�Vh�� ��pB�;,	>af)����춀�+��Ә�p�< _���� ��NVp\t�J��*-jV�+Ԉ����]E�Fql��[���+ؠ��[[��Qm����1�p4�pU��5-_b<��	��/p��s�pu��drF�Y�z
݉�<8�4����,=��l�i8�����#����_�y�Y�B�>�?�&B�V�\�)
]���6z@��ԐeaBD� R"��M�E�����_*�q��!V�U�F��{�%��@9��m����v%#loS�6��)�<��z�Z��8N�W5�����~F������K�M�Y�"��,��]��*�8�_
�]~���=�l���Y��t�Y_�����~��5_�:�sD�� ����I%�YC���);o;�͋��UF���.�Yu�y^�݀�0My������rr�ټҿ�&���e����WX���8������̗���0�H��,���8�Y�eyB��?&&ַ���Q��;��g:��i1"=�¹�U�6��4�s�0�O�1��9ܝ^(5SoE 2�w#��5��aG�Jx�O�Y�s���<ke�&���X(�!c8�f�~����v�����~���%����V`'�ju�����E��"M�[�:��qy
o�`��x�z?/\Շ�T�\.�;[�10*ܰ���;��q�g�A���>��5\��[��H#�1l�Ntڒ��-čb�K�D��g�0�\�O���
���>5�G��Пr��j���b����@0����w׽v׭��,�K;X��`�]�tۭai��	���,����_{l�D?�)ԥ�7Z��E��s\��׬),9Z-��c$�}s��8XS�3\��"}�^ "q��Ҏ��^��m3�k�CoJ��«]L}6�Es�8�J1�X��o�a����-i�N�W֊�#`��j������^�D�z$`n��oc����K��`?�'w��p]T�2Njz��m�~��o������i����F�1���ps Ioںx;VA��7o��)��X{G�ht�t8�B���A�St����[��s�����d���$Dv��D}�_m�#]�.�Go����!�6@�k�Cر���ƥ�}�8Z=��^*� %��z�[���N�M<N�/�DN!m�1��ld�.���W5���=o�4�$�w�u{���$pV<��g뵄_�����<"�ߠ{$t~�!'�2�2���wJ�k$ ����T�#�����h����
�U9$Ι��X����W�塇J�˹��H�p��ۙ�J�[D�����[��H��#��F�w&?oC��%�L=�D�Յ�]�Y�W�=�>:\Ҁ7s�8�,}R��0��pC�m3_J���f����/_�t��,����~s�~ ?lS������:2w$��熪���Ms��r���=�t�L,ٳ��;�������'��SĔjO.|���h#ɶ���4ŐKY��~������_kn����+fv�|^�죩:V��7L�UA�ͣ(>�zČo��*4j�U�ϩ2�;�Ox�����+�UF��G~�"9�7�g����J.������He������N�~��ђ×��=���0
ar{)��s��� �H��}��J|��/��Z��W6я�[�-Rg�A��q~U�}Ɛ�֦��C͸��2f��:VR�];�����W��|�-Bn�PWy>f����)qq��B]��0w�I�G����@���_���|�f��o��s*|B��*Y"����DL�)�}�Uo�NPGO7������́����P>���v���+ٻq=[p|k���$�f��f�F4Q�m~�7�ˏ�$�Q�����6ѕ�]�$)`5�C���$tBާq^/�)�E��6�.5�{��h?T8V�c*��'�`��i�a	�U�oF��fɍ��I�!��}�/֐2�Ȅ�Th4E� �[X�,'���������.ݏ���~���Μ��(>g���惵�����y���nңE��2��0��x�!ݸ��ʧ�wG�9o����۝pl.�ڷ��z3�y~g���<-N���g������"�T��]r�h/��ۛ��@D�Y����R~Z*J�g�'����|h;�ԭ����[����V�?��?+�Y��Mc����~z4��X��w����c5?/ɹ�O�� ���g������`�]�R_.�g,$��֦�]����y�Gw���[�I�T��ɱ�{`�	��[���
�e�,{3����^_�����p:]���a��8�Rm�z*2�L�ZjP�l!�VU�˵��{�NBKS�E��1��u�>����{�ޕ�[A4Z^��/�#��{���ڠ@��fg�$q1C��S���ΦpBZ�;�;�"�iS}�����lg�[R��;} �WÎPY���_���o�:ZHܫ�����޻׌�h���&�2n����������������%}�8(�g$밿Ix<�c��� P�k�7������k@���X�R߾�W1���`[(�o��S��4u�.,IT��G9>�9��ze�8�.�@__z�y����z,wx�����0߹�б�//�-]!_v2�7T\���<��H�u9����/DG{?t��Qi����Xuѷ;L��"^��>�3��c�[k�7�@�������yqwI�.?4Ÿ�R�tu� iщ>�9�Ë�x��ym��o�|zf�d[�~r�����R����J�~sc�3�[�����H�����ް�1&��0��Q��V?p�L�g�/�Ӣ)��}��{�A�	G/j:�d� J��t�r�@��V)���eRe�ik�BtT�W��Vo��ܳ��)��(ǻ����^��t�Ӟ%JF?���!ם���Pϟ��[4I�(�w���u�o�B����}�T���납�#8yf<e��ۃ��?�n䎄n�I?�u���/Wp���&=�M�����u3���WY�;�Ye�2��l�������vS���`�ީ�E �
Z�_(_Mem��`nD�_�������%s���o(��v�\ܹ�Nu�T�9�6#ל�7��4.�ϑ5�NW��?᩽9��Zr���s(*��8D2��]x� ���� J!�^���rK��Kz/�S�� 7���A��D��e��@3TP���e�j뫥p�-�f�D��G�{�.��*�"���/_0jF�T�ֻj	2��m׌��k��a����᳞a;��*c��dg�V���$���b���ة>���d�j�2\�4����(�O�?�<k\á���
Ņ����r���#g/?�dO�1����鴍�1��E_�uɎ��*�n��<���?����%��x�&��	~A��QK�-9~��Kƌ�r��Td�/S��´��ߔ�ON���*�
�ɏY��l���I�B�& ��t��y�)�M�ۃ�;YM�����.�+�WO	��~���Ѽe1�W�(��f�,D7������=P���Yؒe���s$���/���&���O�>ı�����S��#���v��o�����~w�{����W��<�	�,?��OS�oH'\V�4aI=l�Ϩz��T���-\�&�$'�c1�y��	�]����-����۳����0av/��5w�����%�̝�>���񡴂}L�p�b��l���?��� )_��i�>��~0g8(���	��+!��}�@��^�,c��� ��l����� 	
Ɵh�T3�m���'NB�6B��z�ŀ���};���K�.[9��_�6�{}Ntncȴ��P��y�.�.K1�K�|�1� \�/Җ^��c��dt$Z��λ�381Hu��]d�<4?2c׏E� �"t�� �Q�"Yf�1i���<��6pӦWW�H"<h��o<f��ok�"����?�)Q�6��������ÿs��EC����N����f�'�s�Y\m�5o���w���WE}�۠/ /��Ms���	vÌ	�����դ
B�m����>U�o4*ȶ���fUΜ}&`2,��Cy<�[�$��}��s�J���o��6@G|гs�H�?q��&"T���Ю`�k�X�q^a���m�h�o��7�tww7J���0���%%��4�J7JwIÐ.	�FHw7�������z�m��v�'����)�q������jD7+�/3��G����g��S��;�v�����c]S-%��z�d��J��޻J�<^��n�+�:CUpph�/-���ŉ��)�?T ��$���D?T��}Y|��V���"eAh���ҽ6:^J`�ND�iӔ5��T��@T|���.�p��6�2�I�]���ʚInSfߞ��,�Lo��p/�GAk����+
��fM�� I^��̸:�K�b�e��~{A�	�'�/�*�EW��p�u�$zbg��1j����`%��4t<�`N^�.����Zd�t;Ć�ʹ��C�����!�M��e5��_���B��[�G�$�[C^	V_?�Ͱ���n}����X���[]���4��8����.��ĉ2O�K�+�=�FW.��4m�_�B�{#"����M���J�ة0θp*�����+���:ԻRFM}E��ѽ���c�4`ųK�����x�:�H!p���]����b����ƥ^$ʮjg�a75����>��{<�����cU/]y��~�������wKJpt�����̂ٹ�`X�������%r���7�&43��������1�k�"�V���&ު��}����m�s-���8?�x@���f�^�[��n�H���퐬U��~�k��u奍HǼ�thh@ǆ8�E�XԊ�%8��K8�����
"��+���J��l=1Uҏ1x?o�'�`^���z4|ƣ��P�+Xk��N��1҇=7���:��<CB��XE�!2䎕���X�4�	۲[߆v�W�_�~�ak��:H!!y�lѿ���!t"��U$��*�p���ŏ���eY��-5��HU�Z�J	ޢ�;E��1�"Aju�R��;�J������?������X��&-�F]))sƧ��X&�/U���!��& &�.����o�'ﭴ<tǊX##�#�,4�/�R�c�b	�Pp�����і��G��v�t��|)<�l�*�������:gV!��<`�@�E���)2}�_Q�Z��I'���ѱ�镋�yi���1!�PH���6J]�5a(��6:~0>�y�ʂW�wV<@Z��m�ڹ�R�SM���|���q���,]�[��Ь�ܝ����|���gdTԋ��b4j_������մ{P
㾏D!�9~���<��|:12�+���JMy�į��ط��@<��I/	Z�OͽGkh�=�Я��}P`���x���ɒ�\�/F�ҽA|����kk��i6����5
�$�'�E���W-Ȝ��L�Φ;x��D �wnn�z���_�0�:����o�W�r���\N
�w?�`8��6.�P=��>�S�Џ;q�`%�bCvp�2���Kb��
m��>:
�{�cUn�!"�dl9��,�':�v��:%�����.�	���y���W��VS�$�.����O*��d��2�&PA<��+=|;��k�tU�@���8!�����L�sN��V��g.\��;fae̜�z{Y-�C��)|�,g��鬠�kJKa�|7�Ӷ�s.M��`q�׎�|-]PA�0)�&��kb�	y�̂v� $)�ax��^�A�������䀅��a�*�GS�^u�(�匲��>�1�49�h6t���s�l(o��u��/��i�����h4L]dw����^�Q��J�~R�P̦�0<�g
>�M��hv+x�0[�ڙ��"���>܎V:���B��C����6�g��q��Ȕȵ)#���ߕ��|v2�X8;|�ߘ9O�l;���%^\*��[S��kH�&�8�T)��P7������-�o�g��~�&����.����8�"���{I�"w�Y�f��Ɔ��D�>�ϱF�a�@�\�c.a�j����8 O5z�xX�ŕ��9��3��ՠ]��Nz�R����Gg;��G�ydU��ؐC��6ېq�h��&n�pScsl����9l�웩դV��J��Y_s�5�I�E��Ĭ� $.��X� P�J~G���6���2�P�!�{%��@H��N�Zp���{��a��5S���xU�ͱ�U��F����
����j��k�q��ӵ�-3M��{��s�_Գ*�M�`^������a~�p_WcJV��gN�p9�����ǃ��a��@QW@�E}�D�����m�6��O>r���Pa���T�!��(긺Ɓm$�I�Uir�ZO�Xp�qY�ڈ��[�Q���m<� +,�����9,{t*~��lk~��T�~/��H��=!�҉�,5n��I��+1��1+�H�3�O�I���Q��a����
�c�ϯ��X �u��?_@�@��Ə�t��덙u~�Q��g-{r*���zփ�'���R�ی�pﭘ1�(�&�^���o8ae2F�����z�[R�fN��x����!�i��ڛ*���9hLTF����@i7��,���ٶ�zB���
�T�m��&��Z�F�īh��T��2R�=Ssu}��q�� ��U���D�3���S��Q/�ߜOߗ�..mxD���#_�5�^,���� ����o�c�ax!��`t�3tj��^,�nz���\(� v�`b^iLB�"�x��j`��?�I4;	�:q�|ʢ=�{��9bF5xv�>�;���9����"�����V��}}�f���F���Ԁ?.6�����=�E��c~u����O��m.4t-�l

M�b�E�G���a�`5qˣ.~���no@2����X�~8�D[OD)E�稟<O-Md���A�ހH������4�5U� �x�)��Oi��7�b��З�=	f�� �x�d\����O̥��jL��Wk��b ����Q��A9�D��+}��rX��Nz��7���4|����z�R�2�~J�a��Q�^;1V ��o�K`�.��*;'ܔ�IP���M�K�"|K}����I��н��l;��X����L/|��Wy0S��79�<y��aRR#g^��>"�w����g]d�
6����>}��x(�{�� �RF����Dq/�)ךޑ�v�Fk������9%i6���t�5���@����QPք���ߗR 8���� �ŏZ�۷��v�� �	�7�<B�m��hj�M��*׻cn ��T#K��/�1<B �f�
( i\�?C0�}dU�H�W=JV=Fš�� %:4�f�U������~6�yRR6�D�ɷ�j�(7��^F(��}�4�> :��?ʩR��?�:�ቬ`��r�\&�gB��
�	Z18�
O�)=�i�$�هj�W_�6��*�N���-��[���?���msÖ4Ҧ��F���T_�km��>Z_>D���3��F��=~��Ր�
�f��1�Ac��Y�-1�-o��;��u��2_���A�ޏ9���>�M3ræ�\�=�-��$�*U2
���i�ٴ͌�;So���$+��h��}r���e'���6�pl�¾�~�Zg�*W)-4��R(���=|�hOwV�5��/�з���P��)�������YNL>�+��Ih?/�Mz������,�]L�57r��=_ß	'��&<7��\�k��/yx=ӽम�֣Ƃ����Ӊ��,�����,��/W`��s׿|ɽt�qd��5�\0�E��q �[�?�^@�}Xyx��K�W�MM��z���y�N�ޒ�!s:K#�BH��m�}��u��j6���A�jk
)k�2J�Ko7�qE�v�Ǧ����z���w�9L�ı�]/���QZ�h�������P� ;�{���bmU�36�'����Pʂ��`0¶	��l2�CR<'���a\�@HWP��ù�40�)�| �cp�a�ҬoF�3e�/�$
W��������H�Q |���2����*�#q@�����c$)�_�̢P�gUM�uт�Z5�'��ai�>��q�}σ`�����6A���&oDG�M��#J�iF��o��m2�y�;�2��h��y�;98���{!�Ƶ�5죊���ݘ���r\��G ^��'�����d�jQ�,�WvpO�N!9�i�_:�0�r�Vn}d<�=`��'s�*���d��R'�%2e��ݺ�a9V<\�ϰ�/\����T^	+�?���l��ܦI�L٪���!��>J���(B<�A�R�S��c�+������ea������HG,�) �1e�ˁ�1TN 
���G����>y0pQF���a:B��g�1�ǳ�7�;U�]��t����rS���K�W� ]�3�}�����A��<A�ū���c):Q���A�
��o��W��\."�I,:%��/�"�C�\�tq��_t�c�	:v�:�9��R��{�}���D.�:$�
3>�_�af}TT�Ú>�>I������1z�>��;�`����[�>`���.����[���h�Y%��اM�a�U��\KF�t纙,M�k�j_)C��Z��_���F�R%moH��Ό��}YL �����F�9&�9�����q&̞��-:�)�\Rʭ�ux����*m����Sq\�pYnF����¶`�%�R�v|�C#���C�\R9ь/�Y���y�#m�[j��5�/ٱ$���e�ק`�ld[J@.P5G��M�����R4�oX�J!:��%��)(#FH�Z2t~йf<�'1S<]D�s�OQx� [Hì|[��IMP�M�Yn��Gv�"jv%��j�
,\(_9L��\������G� ^��y�x�=�r�}�<��y���j2�|�ag[�m��w>�k��g��V�!Wۇ�rXe�\�{������b�������i���oqj�
��}�1tI[ը/&K5N�G[a�𔵙��9�hFvs��ї8YQ-f����B�o��{`�z�ٍ��Q������Y�ڰUe���k�Ⱦ�|��~�n�v���N9_�GF)�O���o�~��խ�W���wBN��^[R�� �{��ԉ�zYUׂ�Ą�U	la9Z���`P�~�:�do�y���C'<~^��c~�
�� ��l�wCm-��֫@>d�*�A0�w�(���^/�$���͆�nm6p�[^�� <u��������B��|�6a���!��Vf�@?$���Rk�Bs��T���T��ZN�cO$�B�M$�������`��Ji&~��U5����&U[tu?�zb���w�ޕ�W�����5�?dO�h��sT��z��CmM`q��Pi
�%Ҧ���yaC��r�RrsA���37���CK�H:�2*|,n|��Tu6o����_��/y΁4��U�=Mh��B�b�S��ؒ�v�G�2��h�'���55
M{D��M�k� nD��?�?��^K볠[쪷�k�����Ww�C~��0=����B&���
���g��W��A�r`�i=��L-K��J�S��@��h'Y�M#P�_/�Ձ��@d=�<E2.R�
|o���{Ҽ,�`��Wn�K�Q�Ö�q}�����s�ys����c��� ������
	L�\��م[�h@�.��~ƌ�	�/	U7�%+���>���V~�DL�D�92i�Fz��4��y��U�~[��P��x�����C�+�QjC�
q������w.��/�%�{�}�K������;3b�Aƛ0�������LU�A������㭻7�sFIìK��81Whaٯ��Y�ݯ8މm9@1���0��I��ϟw�'M�cJ�I��Ǔ#��ɿF���(b�L��P{D6���?��!q�#���ѱy�g
�*)��A�~g��!-�Wv�
�*�Ty�Q[^�x%_B�4�3ή�/���-����rf32��I^L53s['���W��&�*A޽��U�&����ZK�蔘���qvd�ځ*u0|y	��f�e���z~���i��T)�,~�UK���������̿�?Q�G˃z�9K]���^�11(�d�(P
�ry�W���_!�����P�#7�����x>���ѳȱ�!^��1�9Α?'��H �vNq�{FI���}p6]}�/U�Uh��B�d��L����B��m�8��P����"1�) t�N�1�qC��BY�Ub��Z��t
�:����[�dFD�rLZ ����B�%ϥ�u|^��QT��Xl��T(�����	:�m�ݚ �J�֨�I�6���U�n��\e3X�kqu��TB�fY����*���`�.���뇇��J�)�
)[ Uqzn��S�x+�@I�=��|O1 }x��y�j�S̭�'S͟��~�u��.9y���h�6������25��FY�� �8�3c���eCS��y3sl��.|���g_]��}���`M����ᒖ��q���&#�rJ�ww���`�Q�M��~�_L<��6���;���m���ժ1}�h<O�C�YDO�G�+��������L?��j�W�鉩3��b�y���|��r�x-7�ynM�Y�1[*p^-�iл�N�� ��pٱ�t��R@mL=�d|^2ٞ�j4����s}Q\ć��@&^�+׭��h*B��'�[#��`}�l�o�7�XM�*��2���	����F�R�e�'[��CT���Gv�<���O�Mq_��x�5�ǳ�Lw�Ϙ�<s%��(��V���j5-��|>4���'$;�-ͭ��V���-R��l>���9w�,�;:����I0�PL��[�xݱQ��j�\ �������/�a���V���م#�o,m7�Y3���e�j��������hEF�<1$��%�������e��5����1u0i(Q o{�\x�}��%�E4Mj:��OJ	.��?n�=���
���R��N�z���T6��H��T~;f���l?|��a�y%�EnG��^�x|4.K+�E3p�@����"�U��)ݱ�EjgWNX)��x�ݘh�%o֗0$蛻̄�ǩ�Ə.q�[Gֻ�^���nM�%iuR/�#�ڤ��}�\qNx;$5�B�Xd��H���˥�3�(��ş.��/]-�����Tl�S����}�K�����ݭ-+�*z�5]?z8�+�0S��s�5<{r�8:U;���;,M���6�A�$�1�����후Ê�W�C$O�LZ͎��\�~��	'Ǌ���+o����]��>?@�� ʶe�Z���3���-A(2���2���ǇI��?�/-��^Ω����}���|/g�ps�SH�_-���Kr�t#��V��Z7��(H<���CL���؇��Z^��h�b6ED `����L�>���\߆��6�� 5
�+��3���4��<Nd4s��	�_���w~Ɇ�g��>Q���y�d{���DC�1_�3Q��:�mU`�s��׋�R[�������-D�������/	M)ͪO���SZ��M�֨Ԁ}5۸S��B�ן���� \q93�q1���&o48h��j�Z��"���r}��i �"�5>�VC3ꏹ4�f:N�@Zծh�O�<��)�Ȧ���M�
����������zn��+?;Oœ+�-����p�U���`G�{A��$;��E���x�J�_n+(t���*Sa��4���ڀ��|��`� oYlg�kR���z�%�����;�Q2*)(|�*!��^��">��;�}4�Վ/�=��67c|��ħ�ui���j�yd-�<Km���p���T�֖�+�kǔk�/B_�U��|v�9))X��"�~r�Dor�s�`z��o7)( _>� ��>�h��������WJ��B��r��=N"��aCMf��J���ި��Mjՙ�������vfiri��.i�oI�LE��XX6���Ԓ������馝���f��9���F��׽l+�����4=Z�<��X� �N�X�+Z[xϫ�NQ��˜�4Uf\gl���+��´ìfF�5�6��W
:�h�׍]�|]��0ÿI�e��ֽ������k^Ŕ�">ޣi�|�,��j��v��uz�2�n�?j����o��Χd^�n))p�Z���ft��!��bk��Q�݇lT�A��e����q�>ι_��*؜g}�x�1*���J�"{���;���T��H���^Iv��e���[o�̢��Y{w��f�<� �'N�r��{��1E)�rb <Ԡ����ʫ�=5�y�^&aZ�*�.��������g�&�m�1q���X�G�i��c,I�)ۗ�Fk�`��Q���q�U��ߔ�`� (3�?��Y�׶�f��nz��Oe�L���!��oݮ�;O�LQa�3�(�Z*j�U��8�����1�[��`����̾�z7m�����w���aU�C�����jOG��}1ŕ�����;�q*�5mD�$0��P��j�3�$�=c=�~o|w.�[˾�d�C!P�p��]�#^q��؀��I�VZ�4�<8�S�E�M�,gm��A���%����q\ِ��;U�}@���xk�A@{��6BN_�l)r���F�ז-4$;�o�X�3����.&��~pz��F=R�<1�>�h ��%U�jY��2;
�Έ�\�N/Q�|�����]�hH��X�43��q�Ib���*���QT���U�$]7�f����X� �(� ��?�R� t�G�'aI�T31�n�P�z�5�v��t\.�4�o�9�Y��&^�M�p}w?��ІIwUwD���8�9,'%���k�\wFk@s∜��yt���'�cc�2�W���%;�R��u��E�o�����N�z���t3�:D���ԩ�)�r]�6�/�,b��iÌ��#�HA}tZ\��m��і�1��\�X7�V��K��y�� z�Yh��\T����P����?�Y�0�+L�:����7�u&��#��yt�DUh����qqJY2���&���A\k~��q�	�РBfWA냗��K=� ���)l��/iԷ�$�-(4���<LHݪ�WҶ8&�mƔ�q%�t�m�9��6x�-X��2����z�c_:y��_]%�IP�H^� ����;[���Q���i�%Z�����e!T��S'z�be8i�k����u��A�oR�O��V5�;����1���TŢ��U�M@Sb`����
�أ��Y���8Oh)���M��oo!�d�tS��F{H�*��r�����w<6y�`��b�o���+�"�h��y��:�1CZ���m4Ҏ9���B��$A�#`1�W����I+(5���r��sO�
72�Ƴ�C#<Ӥ�7���h����֢=H���x�pU�3'�[�f������y@B(�"4x.����y3�=���q���ԄP~����0-��TZv9Y3p����}�RbcM���]�''�~L\X;��Թ1YA�H�wDP��/��P*(�Z��1t�U�u)�E�N���ai�E���`�"	��sbj]�{#��s�▗��g���"����?�3w���K������v���Y`^Q��|����4 �i�ǚ1u�%�y�����^J+���T����u�IP�ިd.�����ȫ,�Z�F�.�O�4�W��tu��7
�*���MU���_k����?(�&�g��;��H��ѽ9$�AԽ>��ݪ�8�c6S�*�A�w��2����L(��Ft�̼[��CԺ`�cNY�vo���!�3�ݕǻM��.W�;_Rhp�х�د��Z���^�(7�[B��(���9���q��R�m͹����J,j�)JP �Y헌d�8�>}	�V�m�h��ۿ�wGY>-"�~���	�`�k&�JA��{�Y���tRa�n'�f��[�����ȣ�6ck��@_��?�\��j�^C�4�&����d�9����1b�6���r�2�딶�o3�3��3�.\��/�^mH�9�5��y	#�m��ץe�6R��Q42�q<�y(;1�R�������b��	ZJ�[h�4�:�GJ-�F�Z*j<^8�N+f��tMb[��o�sX	�9p�Rǚ7繝}8���{��n1q�ǁ�iڀ�8�%S�6B1�⋆�tP������,�%�w�
�70,D-�A��x�飄\_N-�.Ւ����t�y٤ɳ�L.�/��4L�^��L��O�<����2H[�*G�%r�W���;�}�d�3��զ��)b�;���}������PBq��'�},T�/HM��~��%�<�W��e�3���	,Im��Ʊ�������~}K�������J�A'�V�Ui���#�.�i�5�f{!rʱ���5
˰���*5-�	B��r66�C�H����#�c]��n�>��+.�ih��l��s�
�Ly�?"���oq~aD8��t��x9 �Ej�C��
�eI�ߠ�>���V��uE����#-n�4��i���nB9 ��ι;<TӍ,���2���B��6Ek;nu��dg�i�5Aw�٤��N�!��l��j���0��Y�\o���k O!��Z��B�湓8��Dg�������8����Jd�\K��I����a�z@�����U���	�d��1x�P��;����zUԖ�H��S�Zvz�l{sg{��Q��x�E-HC#�o-d*�fI���e��������x#����)L�bbuE�P՚[�����&���Q�ӷh����6����d\ew��[����E� �W�,ʭv5��G��'\��W�����:w����t��D���8�ΩUUH;�m�΋D����|����[�m&:�!��C��K�.�p��l,4�s������9e��Y=�%�p0��^ňˎsp�5륬�S����b&@���+G�J�d����Z�)e;� ���J�T�����-�_*3��W= �=����
ȾJ�0d�7�+��E8��w�l�w�\�)(c�0}��\�ڋt�C�:�w�zGD�ԓ���Z�0��e/���4�bI����-�� �/h=q�<�	e>���^T�E�3�����Ne�������}AK\(ݔ������������G=5�*a?���`�g,�_��i(�~	��m6�����~�[��u�>�:U�W\�����8q?W���f3� _SCıّ�������+M`�B[��2���E�hU;�Q�.9i*��A�_fo��\8�hw-���_)&�]L�?r�K�D�&�4�P��n�m4�hC�ŉ�o%��O��c���dݧX��k�V��_H��s�����'�r�C���� P}Bp4�a�Aq����}��"NA��?��!�l�zd�;}�Bn)].�g}�iQ߹,Y�[C������0��i[�D��
�a)fM��q��P�\+q�%��-?v�RD�Ϻ��dLl��ߨ�0�-�`}B������Y��a� ��$?)aK�h<'�Wם����.^3�$Z���1C5��?�pJ��;rV����ɭ~��)���xI��1(
��8C_Y�@���A[�B�Ev�m*����-��R�MЯ�k�-/��c&�`��2�/K�9>fb	Aā�M���<��q<
?z6U�0��u�V]�NxS�k��Ų��?D95�O� ~� ��?A��7��n���O�nqrP���S�ԕ��V�<��M,O��D���G�9�#�S�R��o�G����,,#M�p#����j^6��1�V��j���f��G��`���/�0���L�)�@/m��{�.Y�B{��T����ea��N͡ٳ���[�~;�U�7H��9��Sb�lix*�ĉ��8��{�+(��6{�L ۤԁl��0j������J:����#�'H�|݂-��*�q����d#�7mv�f����sR;`Y���tTHс�+]�AG�G:MV�F�cmw�O��i[gj���.�?7�����p�!��c�D�oX�;sA�z�_�̚��粑�������	��@B�^�^؇�3v�$��š��4إ��s�sB@�<K�uB�nCW�7hOG���#���;�[y��6ņ���EfNlsw4���e�
��=F���љ��]%����V^c�� �G=!�m�-X�[,X�`W+�j������o`J���s�?(�_$��ex�ޤ�ݸ6z�)���F	l�c���4��v�q����B�����gӗ����>Q���-ԇb"1�n�t4�I����5q�h1�c?D�o����2�����w��I�u�^��tPQ��KV޲p��:�]����)(�À���j���x !Mޠ���I�E�l�Y������'���m���	���'>@�@�w���\34+pzY"�C� �җP �lqAg_�o�)p��X؟��ى�cB�;�%�_��d��ށ-�����mGY�tK�����gYx�I75�p�+��F���.��s�Ѥ���,!��|�y6�~;&Q�>(n�RXO\�|8���7C�~���ѝ�j����M<J���F���R�0<<�����y��Mۄ�2���l�t�h���<�[!�R�Жv>����I�z�%�F�˖�#�VU���U���N����f5��v�5���)��E+������V�L�ܛL�Y�у��8��7y/,N�m��YLz[��X�����y��34�'郆�J?dl�?s��6��;�w~D�}:5At<�ǙV��ӪMq짯�NE����	0�)��F	$�lȯ7�t:+ƀ��F��^ŋ4��`4�g
粎�M���1f�?@ܚW��L�����O}��#nL�D�	�KkK�і=D�|X���߰�����sհ>�w��Gy���=؋@�7�u;�.7��!)�(e��Cu�$��P0��K�j�]�
���տ]��).�ڻ��=␹ٱ��EH�=�3�7ŚLԠz�=�䀌�'��W�hF���{O��u�� ���Ã�y�-)p$z������D���v ;�ǧ�C��n�STH�_�wm|c��L����D��iy�&ـ���}/w���\�Z��5���\�[�����$�
+�J��q�j>!ҡ�Z���2k��Ҁ�>�ɧb���o?�	�RgS���AY2���� N*��,�5D�ygüN�w�bk9ɷ.�$> ���A���^�ᡠ�Z,�!��`�jh���[��B�7�SxB�J�><� E�'t�;/���6*�����`ٌ��_���ooc3��|�AU��v{x2v���
���!y���ۛ���w�~��6����x����VdTu�}�Khl�y��{��v>@���Yِ����h�:d�r�R����[�a��lY�[I���E��������u��ʹ��.� <`��a�%��!Ye���y vܲ?�`sC������_��r�QR��Ń��Y��:WI�	���yL���u�'��C��cJ&�qQ��0�ʇѲpx~p�ly !:���_7(=/�t��.p/R�r_
I^-V�N�w�����8Q>���'b>m�<��]�~�$i:É�����{mK��� �2��t�7tH��(��gq#B�"��j*ͅ汘^�N���{�<RQ߫싋��W�߭�ض��J-s�q��g��v����*O n~w�zv������Y���U�K�g��ر�~��GU��V簌@�v ��D{9�U@�X�]�`��;�e����
9?S#ߔ���sq�PR���U�@M�N���/��N��ڈ]D���f� �n��1�R�OSB6v�J�,�Y  (@�D��YQQZ	�>�CV���u#���w�n����c��B����T ԡ$�������/��&�*[��"�T�`��'�$��g'Pĵ�O��*��vN��'hjJ�ehfF�m�dMM�<tE-�T���m�z�F}-zS˛e�)n8�p��$dL鞖�T�B�DA��Z
�b�����j��5lc܅w�~:���e��8���9@៮���sLP�6Z�RZܭO��	�Y����}�s�옭M�p#1<���JT���e��q�=�qQ���^+�O����xj�ឪ?�w�rؑ}4I�z�I���U�(��͡K���\��wϛ�Z��d1M�A�A���/�s���ý �!��e2�.Ą�@�mn��2��ҷ���1l;�f��!0+��E�K��ɪ��肵z�^v/�,f�ӕ����a��S_�ૹ��hX���XR�QӶ��=Q�����4��V�ݘ��;"Э	*��Ł������S h����D��'�4NqN��ś���"��?e��H��X�B�DO?�n�r���#t~0�~|�&׍��k�u�M�=/��vz����\@�h�*U�.е��H1V�,����Ee� ��b=�"�Z��Gr�T�Χ�Y
ukukǁ�G���\� շ]�� ���w%�͕�ǫ����1�|�+�F�j`�
q�-�x�6�c�g��Fr�e���6�i}q2�Y]R}�
����U#xsM�9㻆�I��m��Wݹ��w����uœ������M��D�J�7O���U�%�H,b܀��d����kĶz��imZ�GIwO�1КC���������g{���&r�@�s����«!<H+s8J����FΗ����%\9��X$л�`*�k�� �E�G �!��T0(����o46��	�^U ����saE��$�w�g��aJ*�YA۳�������&�^;�ϫz��WFGFƮ#������1�t6\%�*�A:���$ʥ�6o���Xa]K=%/r?!; �ϗCx�H���������f��/i��i�Gƣ�W�Q_��I��͙���4��"��e�:[���"��"7��I�� �$�����wP�`���_T��"�6"fo/њ�|����}(�N5�Y�Y�%��"�w��L��~����Ħ���S3���u�h��n��x�
:87���<�|��:�b��v���oD�_����$����[g������B��Rg�&��և ��&F;kh��DZ����(5(�_f��������dZ��'�����u�WVִ�,����h	�l�?�ex��n�g��@v����+���
g� ��ED����^\0yC۪���6�aB����uFi��ޒt��B�k�4+j[����ZRTq1w���'�XK�i����i��+.�=��qW�r�BU��ы~[��U����'��iVi-SSGd-*�[g4��H����7���z�o����IW/�UO���=��[/,�Tƿ#E���l��%�/�Ԋ�O���?�~2S�/U���z�i�)\g�w��=3��&�ɰL����{l�܃�яƕ��CO9#ÍL�j�#�<�E1�t���-���+mI>.���\�dT�>�:�4#��"�;�߰���Ӽh�QQ��r��t���q��k�c�W]�����3��Q�^���t�{Y�]Аf(y|KH7���k)$2��W<�.���V>*���3�d��<��P�Ȕ�c\�ǀrQ��S�����w����.#LѦ�}˰�)��D�o�&�ٔ���S\�%����{:��D�s�Y^Xo��C|09��ZP�<l�z���^�Q��	V���F��'�PxT�����n�m{X;�]�4e����+(K� �R:�}(Iz�\���U�-8�Y��X�&�r��[�P* K��iN�+�[pT?E׸��5��DЭ���y�e�MH:��x-�l�49������0�X1.�e��#�ܶM� ���a��O��h}��~cd��	M�����.+��0����ۀ��.�7�&�4�e�"�� � �����DC�F*}��z�>�]��NNW�Վ�-1}�����v+�_m���-�5��a�b��C�34��?�.�{�C����6[T�8���:#�)�-˯��:������sM���ڈ�5o)���(o�R;m�	���s{x�7ۈ��zM�[�^��zW�����(�b/V6�%�V�r�AW/�9ɑ�}�<���7��T�cƊ���^���	2���-����x*r�yW��U����ϯEU�	�c����n�-�b��Fg8����'	�	]������p$ƴ=NxKo!��E/0贤�)_�B�߆�������x%���<�T�u3���ls�/PQP�3��@$}k(F3���"��v֬��<����;��*���@K�|�տ��B�Hb���5z��:~#c���KY()Î���oTs,I30����r�z�������A�Y�5��02��$ޅ!�ش��Fd�����P���a'�5d��H�����w_��DnxȖ�3 \�����{}}�[ru5۷�u?�؈�M(���39�2=M��#_7��r �����b�w�ɘ<RV���Q�35j_�����S|��s	.��eIڼ�����k��E������}�̈i�пn���Vc��e�����ޜ�wޒ"��l[<j@�L~�W"ZT��F����2��l����
c�C���x$㪟؏Q���f��+Yȍm��/Rpv�%5�7�����n��!k}���o�[�U���3��m�N�J�]@A��������Х�=� UDDz��Z�" R��H��Cޜ{���;�sތ����מk�_Ys����{3�������Yn�hF�?�m	$+�O�
X5t�)�q�|�#3sf�^�ǩVxl�~�-�����Pk��+�Ǻ��^q�O��:�U�I���2���.�ܙ�����?#��p��5%�؝�{��Qg/�h��s'��<��ʊ���ҒO0y���n��$��)��AF��3��S��9X^�%o�	78Ow���3��5�W���&�!޴��iki^�]�YJn۪������]AD$@N��|7c�.Ѧ�_/dӐvV
Y_�Q����M����W������C��T]M�-��0��y.G	!˜Qj�v!3��o�N/}VUş�ȏ��I������PK+vO�Ⱦ��De-�~?�~}���L@V�����f���=?�J>���Œ"�}tՖ�'�áR7��kᇢ�R(;b��7�3܄���?~������t�8l��R5�Z��Z=m8�F�O�OS�E���ѮC�?Yˮ��އZ��b�"o��%�_�W��Ҿ~��U�}[�������sss��4���*�)�3��nO��Rj�cz7��b�b��F@Qs�?���v��Q	
�m�l^�����ؾ^ˌ����	Ȳ���Ѩ��v0-À'R���1��Ϛgy�ZX�T#H:�1`��y�jL��Sc��M,ֈ�?k�4�C=�OZ��wI���lO��DBw"�mM!{���/rj��%�!^��p��YK��	r��?�@@����x"�P�M폨ɯ�g)@��R�������A��@|y�~�L����+y+ÜK�ڍnw���Y�;���\����C�R}���=]���u��w�mHo�g�\:<���H(B
�#Lݍ�Q�x�^��<�w��ف����I�!e�����%��������.�%B��H%�8�$?��-$��u��z]DH绿~�16�uB\��#Dzc�|0>�*��+�_*Eӽ�??����c����V�z׹�����cNy���Q��o�c$���/�
�9^���^M���&\2��%��z6.��4D����a����^
���z���*����W��	II���|�z�	���|˟�&�g��a5@r6HS��e��O�=!��i���[�d��c�l�1��\jwv}�S=<U�zV��]�HE���ߡ)��rJ~{q����Qȁ���Y�"�ܧ�ew��a/�f��Z�LZ M�ԡv�����D#(*:�S��׎'l\
G�R-}]�#�C�Ici�"vn���ٜ��KzzQW
�1�qY}��0���Rp>A��c`uſp'�ܫE�]%�dS�to�@��CyQٴ!��w��C˴��]Ln,b�zͱ�Ed�R����m-�6BP����5* �h_�j�Y��݀���R�?��+*Z����%l�(3�b�0��g�4��'f�Q��?^�\���
��K�~����@^�׋:���,�����/6hH������O~?<mV+z���_�\�O>|k��>���O��&�HV=�-������Z����2ܹ@n��A���_1���_ۮ"|��5�Z�ٍ��Tl?�ݚK��<Zy��=ە�y��O��ӷ���ΰ6*i���T�8�Fc��rW�9��ޝ}(��,�{lS�k��g`�����ْα�}�~�Z�ia�w�5���@<%W|�1{v&&��`Q�&ꥅH�F�h|��B�(�O�����p ���y��WԹ
��d��K�$�3��	|��L{�)����ک�k_Y�)�Mɓ�TfiJ`A��� e�T��o!w%�JARRz�FAo���c`�!�d�N�S �4��3��<^
f8��E�0���X���Knßʠu+���p���)/�w�x0�W��m�~q����T��6���a�L��46��Q��V��/�`~Я�	��ʶL�~H<h����[���m�NN?�밓�D�P]lp��
�+�B��K��$~���~�%A=�S���L���DP�*��� SF�<6c�����/�Ӝ�I����Z�%ͱ_�A� �K�����A�5(4��p��;*�g�������V�S�Ve�淮ݐ��?<A�<S��� f�7\t�v,��?���� ��l\�%/�$��fFhk/`W�*�@�!
a�i(��+��=N�[�]��#k��t�F���}�&S<�������*���_N��fP�z5E�Q�z=�S.M!���s��(����O,X���H�kk�������O�0�xPr0�d�"�zCf)�6�����	v.�&�z����`���yST��d�y�I?��g*#��9��3�nC�Ⓚ�9t3U!^觵NC��v��ݽ5Ͽh�f�-����0��/<��W��D�>s���3��<M��d���33����k<f�-��^��4���P4�z:rc{��2uc*h�)�B<0���U�EjZ�oUF�?�`���6�`�����:�=����n�_$������
ѽ��^X~0��BA7q���sj7�ž�9���u�J>0�V���G ��a���F�⽚�U���ԣnv,J�r>�GQ��E!n�.��x�:6�<���	����'o[���<X���Z�m�z�8����J�]�tOGW>��)L�Tos��޿E��h��*�xЪ��>��jՆl�ȣ�	�D���>6�ևq��|>S�Yۍ_STAG?�U��|j!v�P6]�Jf�u�K^���hڡ��D�?�rzB�,���Yj��!��d���ں��wӹ@�Q��}���D�{nk�D�c2�4a�U���,T��ۅ����9��B��S�gZ�)��b�X�߈^WAw܅�HI0 Z5�cܯ��&9�%���%�ވɑ�j���{JTUss�ۋm��ȿ-�w�ޅ�m�f��O2��J�3��i`	u�;�[�$�(W��U�^}Y����A���[��v��fdh�hE3zO)! hl��	��Ⱥjj�z�5���ϮM�q�e���Ҹmq0`�j@_�����N������^�/g�Ǘw`�ӯH]��Ynu7��mu��P�սMD&ǞO���2�h��ӗ�&3������#��5��-��C��Q�8y�j���z��4�t�q7%E���aTT7�����5�L7�l1����,4���XU�
t�~�e
����mS�to����U�U R(p�]V�.�\��}j���k�@)X�����	+��GH��Z��ж��%m�Gu���j���-`9���.z0:ؤ�V�t�C�٪klIG�����, �ti�T���&�U�=$a��Y��"~n[y�2V;�6�@�_�Bb�e�;��ĺ|#��A��'�[>(nl���$f�ϊ�ZjK^~�R��wK^�#���Y�7��R�>��|�����[<*%b{����2���e̝*�#� c�xo)Y�z�y�3��#���U��Y��g�{R9ԧg���U�$�#\�П0}����Y��L]݉s$�s�Ϗy�w�/.g��m�^Py[m�W�G�I�c��)��Ծ�[֗��Q��,`hOL��t�rh��؛�R.}^@@���h�q�!]#�:Ҙ8�Y3�欺 q~��ALs�t�d�%��G���`�ب�]���r�yD��($�.�P����V�!��*��3 ��a�<��w�\
�i���ȯ�'�݄�ת_�v,q����ݟ��/����?�	y����ǐ!H�N
��&é��In�yD<쾖��U���p����E����C�B�H(2���45�)6ӏgބ�Ù�	����(K��^���HC|��{�zV�L|�=��u���С�:���l�����֥�blf%�]����y�>�;z-HGM��I�����bq�i�`�l���͒��*�Uh�n��ړ�wX�p��zW;�H`/�h��Rt{H´-���z�GTOc�t^�Zhp���;��S1\������b��,��t�>x��-q%�RX��͚�X�q��t�Ÿ"�0�j|M����_�`r�x�EӉ���C=����^G0O�,ȧz��/��)H��fT�<u��7�{]GŤQq�|�'��e����\�&(�A�(����?�A�Bw�L�4w���Z4p�Q6�������^�@��;j���p��/�6���t����j��,{�����n�Uy/ȫ,�����_��h=g�P�ElW�"1����?7592R�,a˒�?fP��`�ՆG0��o*=��X���j�({�Jv^����+t�\��~��S�sn�]���Z���������dI09�5j�:l��y�x��/���7<��r|�Z�[���Н+�Jv�b�Q������>�Hr�x�o�G�Ϟ,�=���/a G�M�v��9o�D�;X�(i��|<alP��Iqt[E�<fk���DtJEGo�6𐔇��P�Z&�C�m��e�2�]��a�T\�E�j�S3�������;��N�����2�,a�S��9�'��4�����u�S��;"I��MM�!;�!�V�N�dҵ���$w��B�*�U׌�c�'���4�l��2�)��_V����}K��M�����i,�]=g�F)`ttc�i�5$z���'/�����L�\˔'���c�V\��KjO
���B�$W>�M�9��pY���=tR���k]�g�_YH&�ˠ'�Z���)t%O�u>��tƓ�-��eծ;�	��qo�\~��)�����S��}
 )��
�]\�k]�=��`�g
�qe�������B�Z��Rps��~�ƻ�����,�K�;�M��#�M�(P�#t�h�	�:�ۡ����3�M,�팂�$�� \ct2��+�'�t�Jj}��݄�|S�>��^e�+=�rJZ[��ZG��3����9�$	9���a$��4M�iF�������<��{�?EM��ۈ����������uA�"�D�#�t����Q��*TS8��@�$sjr��d�*��Lx`o7�����1;N.��L4eN���ͣy!D�n�+�jH���6/Z*}��w��}˦&�I,vH�����_�h�*3�;	��S���M���,��z/7�5jM��(;2��d?�"ٟq�t;B����j}ADN�-��X�ɎY�����v5Zg���͓��"2�5�Պ���u>*���'�U��Ø#`���n��������
F쉛HrS�!I�%I���ҽ��C�`Te���K��(F0$�*�5��>q�,v8�h�:������2]DZ���!U��$o�΂p�qV]4���=E�.E	��&��3l��
:o�Ǉ8�l��pO�$9��} �ǀ%�Ɏ]�&8�j�ɐ���i���O�o�S����mc��)h�
)�UX��`�7�<7)-Kr�㜰��lqM�o��غ�䠲�̋�^���{���;����U��:�}��,K<�F��:���K����n^E]<i�v�L�S|�0��^�Q��Q�k��k����K���~~�o~����xv�ѷ�4}�[��M�$HWaSQ?����쵇��8ƹlGV8�Ծ�u�K�v��sY��%$|{s�Z@w�4=� vvx��>��}<�
Q�F[9�����?<��ڲ૮u���:��s[�y�*B9h��3�#Iv%��\C><)r����?ug�aу(�g0��O���8���Jz]���@����c%�&pj������p�<��&��U���z����� �;Ln�<��T�#��
HFKF�
en�����@ۉ[�^59O��]��q����_^�4�@)Bza��<��VR�^~��K���7���Lc�vf����Nl%x�qvX�90 Mdo%���r������1:l_o�m�*\Tu�ͫk��8*A�l�C��I[K���{I�j��"A1��%���Z��P�����O򙡼�l����+�X���p�	��CO�,(��"4H��q�=��!d��1K^bT�Q݀�U�Ȯ��eN�Ý��B���7�7W�t)�$Y��4���s���G����s����f�=��k?���=��M���q�n%X`8�<���F�Eh`.���P!6���8��"��2��^_�I��9z�,M��0,�t���� �9�	(m]��[7�)�� {a�̨.�dʽ"��hu�	=��`��#��?�����,�^��C_�O�V��?1�-CNڀ����J!���;+�ɷu)��������#��D�/�ﴦ\7�n1�G�q�H}��s����>���*�(�ŰpK�#��ؽ��F�pur��e�G]A���)��~�]�Ŝ���R?T\U���a����9a���
U���%.���m��:��#�^�'f
`yϘ(��>p�?�'k�H���t���	���A��pz�9LA�!S�[��+)_\^=+2iQ�d�.u��p�T�&�Ö��"��Sr^U�huU��%J��n�*�~f�F�=�1�>,ݗ����|nP|%�����t���g�H��PX	z�X=�	�B
�|R� iYq��q��խ�!r\���*Á�bpf���DF�������2MXtx��B������Zo�/<��e�|�(���kS��D�;��z�O�����s��c�����t[�g\#�����=��� =b�
��0g�u6�(���"��v���9�'���f�='���@s�-��b7�W�샍7�əcW�UT�m�^�����K�8�Z@�$�i��yԅ����7J&��0;�	k�������pݭɪl;�~z����2�W�m��hbR�L�a5�2ﭖ��d�̼:�P]�mQW>I�}�c�C�A��p�L�+�v��W$#*l/0���"%q�	R�y���3b��������z����_��A-��[�A͈����K�yq��)墳9Q_V����i��P�)&Ś��:��Ŋ���ߟ�N�[u���t���-;!u�
2f@��	j�sbW���wp��=ǆǺ#�qŰ�i]�hdH��l��t5�ˏsܰ�N���\�cq@nǐw�Q���hS��1���-�(��(�s����lʇ��5�r�/�ʦD���R�2R?Ej�(�P��s�VM�B�{��E�ߍ�d��)[��l� ��{� c���žϞ1Q˓���7���h�>n\�,�QOzF��VW=d�o�Eo�M�5�Np�D�Տ�;��5�S����j�6��l} x��E������=�B���j@M��҇�C��n�<j��l4��]���k�#C�<��m��h�ŜWX'
[TU���J"af^W�W0�ڬQTȏ4̱fyQ�c�HH4�e�O��A��F� ��4O� ��q�1���s���_X":I��0�ȳ:Ǖ���L����wV��Co$+Oi^��۬>_Κ��@��B�&v\qij��׹���΂ۚ=�1��ˎ��xY�c�ZL�el�z�!=H#�SA9��ƌ��#0+g�{^������@�����aU����Gf+���%��R�ed�
)r]��R2�2խ1ЁEKZ1�ց����t':�Қ|#�nf�c#�O!(5�`X��R���6�1b�rU[ǧ��]�V�:���ѫ3�Z>����!���x	��=]�R�l.�%���]�I?��V����
�\=j�1�}� 4���g�*�{j%��C��D0�<�ôػڣx��WQv����0�`�[W��
�C�Q)XL8n��HLe#~��� ��v`�U�����&ސ��bn2EJ�B������,Ѳ�b�~�x�)o-
�ɖ��&�c�W�PI:�f��O�V�����+1���A&$��;L4����,Vl�����Т��l� i��&�_���l[����zV�����|d�o,���/n��c�"�[�Cp���l�de͜�2�ǆt���~�朓�횄rGԂŁ��F�j���ٺΉ�n������_�YY�r�뼨 ���.��o�G<�R>����d����1�L�?w8f�PF·yr��q��B�����up�B^�aB���P��7�1��2�55�G�ᘋ���e�,�Z�Y�--���bM�ˉ0�U
@Ep�tF!�s���ĩ�r��_;*�ӂ{?Q ILyEĸ�nZ�K@�] I����ϛ��!����i��R�B.Q��k�w�l�k�V�O��`�����,�/��N�db� �������t����I/���s����K"b��6E����u6�D�yR�
�C����˺��7u�&]����퍃=z��uEt,���kG-c],� 9yG ��}V����FԈ�oR����b�+o�`�i4�����Q�:+�4�E��7d=���Am{�{!������rAý�*�sl�5����w�d�j�ݪ�<A�i���RK[�t�p4��N��*Z�Dy�Ib#Co���p�ą�o��Z����hl6�-�F��s~��{��>e�ķ����OF,Q������~�$C�u {Et������*�ăV���y/u�|~�ǋ��,�m��!)"��jiÃ��([�������0YDA���垅f䛎�Ob=��5��ا��qy5-����y��p/�e�7�n	S�9ֹw�)X7
d���ޣlz��{9��w���=MJ��5_f�������0{��_���O�pp���"�F=mlMa/�
�<i�9��g��)O�n��Ǿf�H�xd���&@���qۤG��~+�q�u���"���rQG�(��5�E!�Q��`?~�~��
1Q�H�n��Rm�s����$�$���i�\��Y'i��4�(����z����p���X�bN@Vp��v/�f镌C�.3�"�T�um��$�p0��~�o�7,�K���9Ώ=�VL�|t6�8K$+���/f{���fuX�ך���J��͈�<a�u�� ��]�B���ƻ&dx#	��߇�JI��s��W�)f�H";e����Ŋ�{�5�m������.$ Ğ$,r&�(�g�J���]�߭���7"�O?Q�O�R�"��=NS���0��+ p�J{��Jd��m�X�>��=zߨ�����[ ���*ח[ oE�l������rK������W׀F�\�A�3����f�"��^]��VT�vП���t���N>�5��rFZ����Z�M�[�~�>����:�h6���'�D�ß��?)R �h�|]��G��}eîHW�����f�N&�VC}���M~��s/[>9Z�G�a?��2oÇ=�&ں5�gX�F�Sg�i��[�R� ���mҮ�e���]4"�Y,I�%������
⊩��Qt�>�����$������(Ģ����R�z�Յg�q0n�Z�ĊE|�K�DN�,�M�O�U��]^����&�V�}�6A��Vu_Z����7�`�u�������p`MƯ]�M�K�wr"�7��χ�^�W���A
s=ͧn�r�W� �OY�%������ٌ��|�jْ�W�˾ �J:�����z��f_���hG;^?S��9P�����su�TI/��n����^��tu��{�)Ư��躻�$��Q����+M}�ƨ���|��M�o�;J��E�On���Djd\��I�$��s1�Y3_����Ǿ��t���H�=J�ܚ�7�#��C�Qb#X����b� �y����)�ˀtr� Aj��[��
E�/P��ruf `��K.�74��CX�T���'�[f��ז>?r�TC%�u]��ub��zJa�Z:	�X�ӑ����� �v��+��h��u۬|�>~�f�E[���ӿN��jIƺ���s|��n�t�X��hxJ!2R�$�M��5܋�*e��Rms������jf�K4-����`"���\�A�Y+|�����#a�/?"�X�n���ƅS���[�Tw�H�	;Y�i���1$��V���g^Ȭ���@��2��1zRv�����@�Zq�]m�6P7g���,.���",rMlr�D�s%��!D�2�P>��ûT$���P���p[(u�v(�m �l�Xy�����	��_<���N��f@��,�eE�޶4}��Ud��o��V�ȅѻV (~
5γ-`��a��,��d�˸�eZ��NAR>{6(]m69�je���n�e&�$�FU�w��)	;7X!^Zz����Ic��y��dͨy�^���|�?�6ٜʢh�F�0�ԆEf&nm^Y!mx�#��Yo��~^�#����7�E���$RBfFP��;Kri��(�l�^�G/��Ӆw�������F�f�38H�atA�p"����|��3�}49�E�$�R"0D�S��c���(�?sZLdT����ٛ<���0g��k��p� �����ry�'�{�ʷc0����y=�h������0����l�.��.w�����Xc�yK�O��~�_����Q�� ��+?���.8�voJ/�eR4����qP���gYTt�,��4,ޏ�7B�Ks��|���ih5�G��M�ƻU)��

��"�x���k:8��m�!�H؉eH��'�oW"h�!�s����d���,�q����%���2z�0�g�m]Z�v'.��H*0�IR���aV?��IE��xo��'!�0&�U�ߨ�<��#�u^os��M�=�ߣdr���il%:����>c��|
i��n���_r�|���@�.JJ��?��_k�N���KH�>j� ُS"��צ��im����ib��tR�.z��F,Ȉ�\�G�]4�ai�3��<Rڠ��%�X���\�_���3�&��A҃!���<��rB��z0�I�J�;��E���8�)�ƺ�0����	C���7����E�a��n�C;�"B��#������$7˓ͧ�~Y��_?7����ҧ�MîV�p��,�q���Ʈ�)������0�N����[���yO�N�q�=0+*��I�T2F~�!i}��&)G��_�$�G'�j�Ξ�v_]�H�b��������(��I�Jt��b�@S�bj�Ow����:D�Rz���C�;H.�+�K��ۄ�
��3��e�� QL'0��o��H�cc{q��o�^����xI����{|�vvE�q|>�B�m=_]:���GN�������!L�0Y�βmt��oT{�Z���m=F���w5?d:y�j�Vۆ_�B��aK���
�s{�R�d�-��΍��3`PXiR�(�^^୔2*W�YD�彛Y7Z�0�Zߪ<W^��6��C����Nn�W��\IWo��#-5p\�_ڥ7Ɇ�H%����pϤ	��k:�k ڌ��凍Ig�*�E�b�Ut'\���<}w�NڐN�H���O��̼�4���t ����g�<�����nr�c�c*c+E~�<���#PժgA���TC�Ũ,�h��&}%=�������B��K=zws��8�q&��#�L�pU��q��	d��]�-�ѹ�9YXvp�㒣k�R�M�;��4�fsT�h���4��N�v��OVgA��&$=c�Zh�����'i�����WD��b�h�"�'��i-���"7_a������,\�����t3�
�u,�O���ki��ɥ�}`���5e6�~3!��OI����u�uѪYWo�3���H��:r]].�40J�bn�Y��������;���`f̱������0�����J�}�]�l��Q�������$�)�cA�8��(��y��M�[�_A����#E�*�ϛb�GWd��m$������"�Vy%6O�9OB��$�w�Pe�G��ܧ�	7�d�>�ݼi���z���%����d��2JA2ǩ'��P��K�(���9�xb�j��=�WUk�V��2&Y|+�C&�煵�ƈk{�)]��"��M"cdiUS([�z;z$��P�������r4�`��QXK�W�_4�p�WV|�p�)���0��#�<���>��\
����h�#I1&t�C��-�k�0�mi̚��q�M>8�V��f���[D�����o;'�����Z�[ANh3���{}X���҃��{y)ӽ��gW�,�DɎ� �EES�{�tz����	����2.��F�B���A��z�=
�]J�Ei;	:Eْ��˙�pn�U����|�k�T06���'ߓ2��L�8	��[鲋��sQ =�%Rڡx6��r����zQ�|����uԺ�W���Ò��ϙ\�P��S���"�M�=�{�d�$���m��R�$l����H�ۓF��n��BN�E�,y/�N����Õdb�9�Gfh��g		��,#q��HL5T�r��T%mF)�j��Y�.����]խW�gՕ&���8�����*#c�Z1��ϮKG�zC��B��������>���˸��j������,�5r|c�]ep�5�;�+���Օ�V����F ��X�/����'����wV�����K��*��V�5�ļ�˪�8�G<u�/$):�8b�ܑ^x����֫heѮE��恔Z�_�
 �����p��A�>�C����/������PX��S�,�1k��LW�:�����pK���R���ΟƅJ�@��W�ϾPb䥨�H�TD��[A!Tf��$�H�W���()��ou!����ܿ�b����������|t�3Y�[��S���^�0�W��J��g�F�����D��T��x�,lt7��l^]s�͊�^�^��ݞ�u+���4����I"�d`�Ԧ�5��w<INQE�(���߀�H�� ]W����$���6kC����S���ֹ_��B~CE%+��h&�y�Q�p�Y�Ӭ��&ܦ)'��[���q[�/R80A��Lp�j���'uϙ�f�ݞT(k��r?
�
W�~y�*w:�������}�����Ãդ�g'E�++���HH�}���(1ZZ�)�3>��Ƣ������旬`Ӹ.�YY�cmM���ڮ`�n��0I�C�����Ďh�^j��E�BM��:Пn�J{�`�Y°��\��:� #��1�w���>��-��5oR�6�Q�|��wx�!����$$4uS��U�:���8{�@⪙>�%kֹ8�m����[����,�G�X㺐II�TCX�KVhT�E��#*SM;�\�������CAz��ɌR�[��L�H3��qS�:��Mr]Ӱ��^{���mys�6ӕ�^߶(y%�i5���~��~b�]�����G�c#�Ý�4}��ՠ
��5'��(����(�[!��PCyϘ}3X��~���N��{o����P����џ�.��v���I��z!��9(]y%9+�'{�*���[�'[�����1��f�-`uz"�?�
��^-J1���t��z���E�����bl�h�k�s�^v�5��.^�,'4��ӢK�֥�	lp���0��7��+����Iӎ���H9c0!�u��&W�0p�=:����s���0���+s���L�U�l��ɌV�4lz<������-HBH���
Vm�S�q��O��˶j^������.?>��%�i\��Q���m���7�m�#\%Q��S(�q�;���J�D�����A?$A��U�^�(�T)�{��蠼aa"���)�A!@3ըY�z�I�������J�\:�󣴷������~#��}�-�\�7��A�M��	����-����ϰoQ�φN"	�������=z� 6T.��ē�v���Lz�j��v�x����MyS !��K+�>�Z.u_�C&�'L������K�$�g(��_�Ԁ�!4���J�YV#m�M"��A\b��D��_nS�l��пJz	��2��\���ؕ�;�������p�Q�c;i$�� ����b���b��#�q�`�Ja�:�'�|�[�r�WN�,	f?��b��Pf\�t�l?����%��Λ��Y[&N�|��_ԕfOD+q6�-��c��_�3�:�3�>�l)7��;@��2�E��~�В��s������x�wp�2�w�Sl�BK�e6�^y����޻��h�/E�!�	�_ N�x�g�R��(��	Fȉ/��n�^�6E7
���/���T��e���������|Q�d~��PCC���aC������uΒξ	�����@"����}�{}=�`��ͽ��|��w꡷p�O�6M�r��-'w�ՍH�c�@	�O�
��Ƚ�5��������M�7�v�>n���V{͌l���9�,�}!	�u��
Z��6Bu��6��35���h�fx�<���:����7��
�&��
4Ƒ�?�nߏ^� Vd��{6>ķh6�l��o�5����>f��2!P�5V�>p�H�U���؏kBEQ�x���\TsQR�����Jla�/7�/%�����¢��OU�n/_�������|{�T�iA&R�$����{C�Ԭ;8 &���s�e�u��x$1�ʺL��!V�3\8�B)$���~�����R�GvO_"�^�ӆh�	��P�>+��F=�y��';!a���o�	����8�"�u��ߔ���(�2�Z5�PK+�X���b�X���7A���.�T���u��gԭ���~���˜2#��q'��zD2��#޹�N-�0^ �]U����o�/����B0J<�e�V�Zqm�^TC�G��բ��o)�9�@L}�|9����J5�^�V%�!3�����5�c�\��2����P�^r��}|��	p^����(}vD�bkYV�B؊@�'PQ��y�
>�[D��ӵ���ܔ/:��^)�|pc��S�q��Di�s�f�$����.�3�o06z�e�cm�<���_�a�;�i�Uɱ@�qK��P�Zl��5�=���ĻEny�;�N�OvA�Gvk�S�ѥ�d�/L�P�Q9q��$� ->������N�~)����?�P�AFl��f��M,/��{��8E+�L�K����#��zKSy}��jQ�l��hj�[�e_�kJ-K?�|��e���}.e�����B��J#�G����(ͽ����D�B7���M�����/��l���eR���9����Q)lk�B`E���n�%@�%���|�(���{�/��� M�()�Qw�3���315��
c����b,�'n�e�eJ���[��������?K��`�4���v
	01k}ы��@ؘ��F������Gc&�w��Om����<8�U���ɇ�䤤6ǏjMġ�:�����+P�Ȉ�;�$46l��~�+{�%MA�,�rA-�vV~%_�����.%s��іMk���{��6]�B���_>��]5�w�u�"%�S�GQGk�Df�s�-��<���H�u��ʇ��7� ����ե��I�I��?n�i�',�'�ay���V�d<���%���L���
t�$#!�]Z����[�b�Ԙ)Aq�/�/��-���~��[�c癯�~H���XK�֫��߬&IQf����,P��ߴ��τ2Q
S'��=�|�ä���=�(Y��]�Y��/��.���(�����*ϫkMS��B4�3٦ق����D]�Z��B�T�oNM�N�;��W�����/�'��i��,�g��.	�0!���>b�|:o^������D7���8ZbW�_l��;�D\:wN݉�URG��yxYT�Ļ�$�#$b�G�OZ7��Q/���٦�&���E���?<�;��ļ/�^�^�����N��'�/Yvh���g���<�&AYwo�ji�<�O���K�E��K�NH[пz�1��3�����Q��z���F4/n�V?)!B8
���6�+���N `]��|��f���p]�c�(Fv�T~��~�+|���#ׅ��R�U���
�U�_�{�r��r���)1`����&o\)�Lbv_�F�k>,��eD���L��q^�U ԩzz�1sk�7���������Y�!"ځ�_j��i�r𫞘�ʼ9���׿�bB뇵�Z A1&[t>���x����j�T%W������R��-�z�Y~��m��%��Z �/y�����˅����;r����]����u�Jv_�㖎![mf��Yh�A9u�Ph"�ٸ�ƽy?ɓ�\>$`M�a�:(�\(3�	;&ro�.�!z�'��ޖz�+3k�����r�|`X�U�]�l1SJ|J�7]��r��,J����r��f����A�O�@�/t*�o�:x�pM��G�v�S yrQ��%]�x����J�r����_��kwLh�� ,ֳәm%��s�&@�0Lp��-��}�iNx]|8�ۨ�$1�?��3�w��������/��W>�<$�X0I�20�ǃ���>͋.������,P���A�Q%�s9����vq�UKe;��J�`7��-��f(��I1#Oxj�M�s՞����
����E7{ '�@,s�/��ǂw0]Q�B�^�f�m;$�Vno\[#-Œ��gڠ* U��}">��6�����nf����M����&��9���K���55V6qEq ~����F�_Z@X�Q����m_��%��52��ʧ��ޛ�wh����s� Fb	��3��8T�>LU���ĀQ���B��� �n���:�������V�{����fۿ[��m��ԪU��^�֦���v��&�U]F�-�fQb�إj6�$B��4b�q?w��s?��^���:�����<?�X0���Hc���]�;�D���6�7��R�Ne�^X(�܍L�J �?>9��$�\��B�$US��M�&�
��@�f���g���].��:)n�Ǒ�."�i�?6�t#��v������
"�S��[y^��\x$Df���u�-O�	i�=���G����0;��k\EÑk���/��*��8H	��T��[��@Ff��-衫
M:��+���wض�/�z��_yH_&R�b��+N����P���n�R�_�[!7���d�:�";+]k�'9�^Q\�l[�}WA�ڟ��u�K��$j��WMCг������I,����|�*��`"��Bnk�����7��Ui7Ēnf���o�p�k��I��H�H��2�l�MI��n�^b��������r�,�.���ĢY�ϐ�k���Բ��G��7ן=��o ����5nm��i�t�QU���[�F&ۼ�}��駷]�l�݁�]h�3�DכeS�VE8��\0�&7���gYE��	�,�Q+�~��_�����L��#3_|e4�f��`h&���_�D�K��m�Hw�=�#}}y�ddO�ֺ�t�_4
����.��N�zB�!H��s9��Om$�6�j�Ch��&|�\��c?�b�3`o	�6;��O{�#"�^ڠ���ң��fV����(��)�v��]�Hh@�7��]�\��H�;�D�0��6�up�J{G�Sו��j78�\�B~dvGL�.82��]�(eHuA�H�lyF%�V'�o���%��;�<�����͒�}���#�1�o�f]� g{�@n� (���T_���}�alg
)��"ªLD�/�l��iM��xa�o�-�����"�yŗ2�� V�%A�\�T�~S�������������Σ;>k#����*�喡��褿����Oz2K��z��qj^t�&{Q����dp�i�G�)�
87��������=8�N���!3[��%� �����x��|�<o��E�m�e�~w��M�,��T2�	up����]��CxTl*	r�y�C2�kŽ$K&=��-}C�}�*��0�D&�[T�Q*:;��sk ��]YbW��+2�{�<Mu��^n��(I��R�	�禦���:�x��Ϛ�6��)����>��Iw�AN"�����Г��;�G�i�j�00�˥��q�R�6#SC�ǅFf�<�4,I��8�_@4mf�pNDTq}E=�~�n�[Ƽ��cb��1%<��ς���XB6Ǆz;EɃ����B���G�����>�z2��H�өL�Z���/˕�4��<�2���#�4͢l��
�T47�Ec������w�������W��V;�O�?��L�=��`1�'�.�t2�63��=��>ցf. g��x��,*���va>��ޣ�kY�O���_,^�M�z�c���e�#�����F!d�$�n ^"��ڶ��\hC���I\Y�m�'�r��5iv�` ܳ�=�8�#��2��A�G����J����	�}���EH�,_��6㨍�6�2s����W���Ҳ_˟\s��/�Đ��q�5b����h�y��[C=���uF�$�{��{���4t �x��A7n�"�����rڊ��b�mTXΤ��{Pއ�GK��+���w��e�w&�D�1�\�ή��	x��qRO�#
<�c5�o�z��I%P��i���Rc�%�8zտ%
N��� w�h?e��t��!z�nI���Aެ�����_O�gB� -UZoRT�?�����H����_��x��_�lH�_W�LZr�F�8ޏRi�Wr=�G��Gc{*^)��O=]+]�:���#2�/p���Ne~ؠkc����w/�ōVI �^|[�Z��z��8�#J����$"�a�h�C����yl�߇~fҌ��z{��{܏	�h�-_TDM�/��͹��M��?jh���+]/���u�>
[x��UH=%�$�U7q��@+5i.ru�迾��/�۝9���E}�w�3P�~cǲ���W�t�Տ�瓺\��u�4�\��jO���A.�6x���ٖx/���>�[�P���=塦`)���/�v:#�)?���y��k�95,�/�`Q�3�Uw��%O�����D�8�*��t8�3@�3#�ds�d���S��;�eZU�˼q�W�k�v�2��,R��Zo=9#Ra����`B��e���w�Oצ�7������:��f�)���d
��Sw��DH���y��F͋�-��t�W-s~�]�!�s�z1�yN����OLX�9IvPi+���#����:�>*���˨�D��)	�g��Rk`j�l��-)����joo�W�8_#ٿN���hr.�>_r\��u�͔�[:��5����.�<�!�r��dy"H�]��[V�C�Z�r~����e��[JGN�J��6	��)g�4�q���4�>4=��mmOӎ�Ϝ>x��#��z)7ӑ�LM>�w��]��A���:ڿh:M	Y�A	�u�%�C	sn��:���r���<���f��^:eQ���)4z/�@�9^�@=R��=�<��%���K4WF%Ϊ�P~��������˷���C��z/��˼�Jœx�jWV+&E
F��ZRKB%򑤾J�qǵEI,4躍WP$������`E```��й,��Ӛ+��C˯N?�o����6��+wY���g|<̊��	;S��&��9����n�0���{CX[B!�	'��X��U� ���'ÔMo��ɊZ31�цHN쓯I;t�/�!4r�6��º+c�"�����$-VJ�H���_j$p>[�g/|�Hҡhҡ|󳚉ڏ�E�e[��h*�jT�4�M#4�������'�brOO"F�(S����s�����]^|L�I-|��SH�����Ix�2E��2E{ �*N�[����2W]0�caR��媓޸�|��I���͹^�h�0���#�[S�tJ���$�6#N���?-�ǝ�����ؼ[�zi���c��2�&4[��ue�'�	�^��(���@��Ni�}����j���3�k7+�읰�D�P�r�Ι��T���Ċ8��!'��c�W�����I�פ��1���	 �����b���Y��a}إg{�mk����M]Q�g�A`E���������<C.��E):A]6��`�)��H|LޯnDc��ϋ�vg���OTdM�l��cJޅ	�_����q8��f}�3�H�+抴-�Oc�"��ər���o��,�?��J�D
���U���
}�{bf٪wW���Q���yo��\���U����"�����^h��|gdW�$|�~�/���Ʀ��a%�T���Ʉ��ir-~q�$�e�m�t
V�\����V�>kFP!2�{a�@�B�C�5�K����K��`Y��>�����S�w�wo�a%	�b��Ä&k2��2�����5���o�H�P ".S7�<��&�R���O�`#[���y��&*(�K��6	̹���.��L��d]�o��e�z�X�@�/�,�3HE�ʍP���$v\�CR]>~�)_��mBW�Kn���aA�E�qZ���w����L�G�3�{�C�A�o\+R�����q`&�'�%>6�Kؕr��IN�ZR<�J+���4�窀� ����9N&R�{��}]��06�d2�{�V�X��nA��T���zf��$�y��҆�UAO��G1 �c�S�$Ӟp]K�ߣ�����q5�!�<}��'� �&5�k�2�/�R�{��������N�D��R��'�c'cz4g�A�i���Ex�ű_lt��5�3p�g��T�u���mj�W��Ƅq��▽��o3�gR�q���
��m�N����{�ڽ�7�5�P24s���~�<�rw��E\_�1�Y\�W(���xM�Y�U1S5�"��N����Ǝ=�`�'S=�$����%C�>���*A޵X�@IaG
��ҽ.��H�3�.��M7��J���!��V�d��*$�j6�v��Pڕ<��S`�6� 4G�j�rK�E��%8A+xz�p���c`�:��� �/���x��UW���+w���4fżS�#gQ�ks��i����-��%�+�����?�2���+�	�q�H��W�'�cc^�+T�<s,��,�V�%�z?I�1X���a[��ABB1��"d�v�����^�c��IZ%cl���0,6	=��3�e�w��A*Q�O�
~�����S���� 0lͷZL͑;���lZ|���2�&�uh����dύ��A�����O�T�q�'KϺ�0M�AԯƠb��f+iҷcV�"6�f��IS����em����6��:�����^q�n�Q���`�y_��ڸ̖�h�� č���������O�5�"T���G�w���_a��0�Ҟ�k�D�j?��qt�(�O�A�-� &YsB�c�O�
,k�t�h�H9����آ��2�wc��ѥk�ИյhA��JcE�c�%�K����ح����;|�'^s��[�nЊs�խj0�X�%A>�u�$�=��NX2���cØ �g���l�tK� �^�cd_,�>f`�X'&���UR��^!Uݣ)g,�wlU�[k�zD��`���L�C`�d���vƊ}_��4��� ����=�M�ɪ�R�Br+��`�ɷ����U��4"{�ٻNr�V7�A�"��-JO:�������`���9pH ���W���_[����1V>�"��8����"�Av���;E���kAڋ��#7�:تJ$���Ӿ�O�ߌ�!Ѻ7E����N*s��r�yQm׽@�� F��\�,r:�����!�-���1֘�Ťr�SW��j�=rn��Z7����  �(R�ڣ ʲtn�������N�C!5Y�Y�'T�����0ְVs���ifk)3�"�538���/��-g��J+�^��`��Dz@�!�Ï�D�e�G�$��&sʏ7�	��@��j7���J���{��5��_~{��q���O�E���g6T��\Z"��65�����Ba�B��#c _D�n���yb�#aSi���ƿ,�6�Wv�V�)�m�Mg/gE-p]9����@������

+) �e����ΜleK4>�d4��V,����8��Zuc���)�6���T�?v\���h��:^\NH/�����q\��f̩\E�k���-߀r�$t+�i�ϸh���N�U	�"��K�`yQJ�[񬁰�bqA�1iw_ŵ����G��u`p[]�!�P��^��ZN��I�o�Zޓ��֓��ˉ_�n��Ġd/�)�n3ە�����E�8\����)�e���G��]3��m�P��>�*�H�瞧F���j���H��_����}_Hlx��'�ro@���ֺ�ag�[Q�-�C�X�J�Y��S�wȨǊL���v���h�f �!#d,O��ob!�?k�CM�Vu��Px@	d�h6r� ���K8�60f�����>q7�P��k�j�ݥ<�OL{�"i�Gq��Ñ=��Z�Y�῏H/����0E��B�l�	�]�m+'����������Ϥ��/��g7ω�5��*X'��2Nr� ���2�DǓV��;Z.-Ua/����<����J�
�Ŧ�j������ ]�=�(����k�M�vϩ �a�V��+(ۋ�K���U�A���� S��Fxa,�e���˔�	-1u�GRC(sl �m�TCQI���97�����10�rk�ɞ1����&!�Z�X�ɓ�RU6{�:U�F�ݽ	�rV%�!"<�K�W����@���j���H��	o}���tq����7��l�(9��H8e��98&��{&`�"�&}���/9E<tGBLC����r�l��.':�ǆ!O.�ߝ��� ��u�X�bDٴ,6R�Cm�^���n��/A��Xļ>x�yF�򺓾�� .��\lm��]�0�5D����n�t5��@
���)�s�*��v�bN'��[�����I��ծ��6QA69,jO�e:{��V���e����4��lP��F���6&�|ǡ{ "h�ćF�X&(�&��H���䲓qX2�!HI�읒⽖(k�[�ox�}i}Ӆ[�4��Ɓ���$.(���	�y��=S]�Tz��ҟh���n7#B��MsLdx�����{��E�u�uD̈bru��}�<�.��?��So�Jj�{����2��U�ᣊ��<����J�"~]�e�<ۙ�M`�̣�-���E���ڧ���z���)�� ��%Wm��ɰ��� ��E�j�π籠Wfm���.�"���gՊ��Wʒ�<y#��C5���hw��l�A�#���0�c���!$�V6#`����M
9���{��"�|W�*��zߓz	�}�`�X�'�̜e�dk�����I��Z�|y��+��WZ����ld�����bR��!@��~�n�c�3|�� ;=Yv��u�@������K�!A;�q��I��[��'�e�N��[|v4���}�5
W�/���|�7����F2�u>�T軕r*&<�SA��뻾�n�~9}�+�jq+�$�ˠm<�zZ�yҦ�s��s;=2��=�"���a��x�x�8f�b^��q����C��X�~��L�nC@���&�m�raZ*�]�Ö�o���_�œ��W�]��p�}�˫x�eM-�[��m����6�9_\�5�#In"?�\��ՙu\�R��c�k�(V-�v+�̰��Vaw��w�XL�G-���hK���-;;aB�bm�z�GR%qZx���ފ�ot����Qgm���=*�%�T��!6�vg�A0h�<2f��4�~n��;2��cPa[Lz;���a�����Z̙AW�<��|��iq���v���"���/U���+0˵�������yʦ�����e`J�u�O'Xd1{E͙bf�m���j�#�+������r�]OW�ٹ��I^w�d!Fv�j��GBV�C$��#9�8T4݊�$!�F��e���<���mP�-Щ�_g�&���.t{v����v�7�{j�i���6�~��]h ,5�5��+V6�$���)G���<�M�}�;ςk�9)�U�^xj��m�uE�q?ui��ލ�|���g��i5�]����ݮ85#ұT6��[do�g~��Ƨ�>�f0��nsU����v�/f0y�\CA���c`X�~ �T��#ŝ=lK'�.����;,�'���]�%[��{{�~s�#��� ��]/�aU����$QL�/��b_�<�"#/�Szf��gh%�ha�W�&�ϬO�C��#'��k��!�$�f5��-�E�����h��.�ZQ�b�6�v��ťqr�l��G���n���љ�]᭴U.�>�_c1�ٜ�e���@kAgy��|V�,�̖�B�E��z�>OVչ�r���~y&⟓�mh�%�r�`���
��]=_ �<4D�_Q��o�%�	�`�g�oR��^8�*@�n�������P�@`��`?�y�@}����":�|��p�MʾbN|U�n6�9�Щ��F�;��e��]�K�ΔE��_��\����==v[y����	S�h�1�*��ռ�kP�'\c�
`���D��L�g�~{� ��Չ�Ld�٤Td��s@��0���|���u�t�UZ
��;=�J��o���qd)��1�S[�T�ӳQ"��5+7`o�Qt9~V$՚b������{d�J?���}�+.->G�	HRh�6L�G$����W��raJ�ޠ3Ow��]���⾅N��b����Ƃ�j�X��7�i�vΖ�;����z���h8`�7�sqW�7��L�TT�	��57T�!���-]x|fߞ��c��ȦI�,�YA�&cC0���:H����=�wS�O��b�+zD�U|3- zI?�JR�����2xv<�~��^3�1��S/"�=za�����"g$ǭ�s�/��安j�2m|�w�i���/U�?���7�\��=��L�׸Yy�Ze-z��̪��������,4Ϙ�=�]��fL@g?��S��c8��Զ*�4|K��5�}/7D|%ʲ����"���ژ`U�[�[|hC-��vv��~����d;�+S���\_��@���	��-�6�D<y�r��,�o�:���v���۠���1�g���!���:�M�9���zl�A�]�L�.4�ѸK8>��GK��*F�n��	��z��D�:��k���_!V�ø�G�i��0����Bf_0�L�m���� ���P�VfB��ǈ���E&]�OO�����e��zsH�Zy�g؏�Ŕ6����g��0@Oè�M@��iJ�t��4	'�F~�1ԑgo�ko�
����Mn���h����@��� h\�� ���V����t��iqE�!����#��*q?M%��Ƌ�h/����J;���Hk�&o�xz2�3򁺆1h�3tsz�#��nl���xWO�/r�Ϧu&	m�q�?q{�Gu�������!�]6�A��b�0x??��'����SPZ�$�"�xN���0�e
c��d���� �|7��wKɻb�i�>�;����Z��	���L��#�5W��8��_��]h�J�֜xX��z%�Ɋ���c��� d��7�����BQ��z��ٓv,�sPI��ٲ�ݱ���mz�ic������
�]1`�=�k�/U���7G����xAkA<w������{~���5��� /N,�f�����EH��-�l�3��m����ޡ��a��X����Mt���ɱS�˱�*�l���;���0���F���YUb�pk�~�r�8��_��EսV�����K�m���&��`bG&&f�ݡs}�:־q�0?�1�-�^\z�-�@�?6��?���E�\*��#;��e{Ϛ��{�3HCs{�k��Q�j��>f�P@6�&ps��j��v(atc{A�lZ��l�5��`��H�����v\uA�h�5�'���]�؋��\��h��Xe���D��,f��r��K1��ZY��4L¿Ѽ+	{%���O��n�Ӯ
ԁ�*W7n��C7b�Li����+�-8a��m��ŏX2�[�Q��6,p�� fEEɥ���A�s��
e	!;��m�ڱ�Z>R	N�L�#��	!ʮ})�Aۍl%���'�\��a��t�.;$��!�La�����po�YF���߻hƵtA��m
y�V�b��4����Cto�@��T"C}��Ѕe�R\}��J���8p����AL&����e�4��q���1n-�}ƀ��L:1	J�
k��^�/9k'���I ����" IR-9!�]ר��a�{����N�� �b��Ԇ��63��{����)�i��Id�(���x3[D��l�h7�
K�rdw�\`�q��Vl|��U6HڟV0U�����O�Iq3+֔=�l����8��LsX$nR<����� 2�G�W�6w�c(����	�q)���ݩe�%DaE�!{����Ȟ	REX���H*��EbI��3�#�'�08�,��z��o�Z�w����^���s{�s�ȷ��ұL�4�7�u�8��
������R,�sP���8��x��6�����>�L�D�~�΁�0��d���,�b'�����@���jP���'%?F۹p`)���	�(A�=�#�vמ���9��6�����{�8d�_�,*>5��x�jM�-�����;����C��F�0�!�:�z�Vv�_������%�]/4�X+��gSu�YDW~9��}0T��4���pQ��<��.V{S�&��1���a����&!�&3�qxX�̟�q���-"��1"�����Q��#����wzx�g�q�����O_���&X*��M�0�T�,�lի�_��=C-�
?�����1�[٘�j���*��Lߋ8���g����e�9.�6]�� �_�pX����J�Ƨ����d�g�'p]�'��w���E�ܯ��R�����y�D?Mo���X��>�Il�P�O�����}�/�oK�bIV��i�_۠}�?t	Th�i�5�|m��P+�P煩%{-�����haM��ݸA9�"C6h/}G�$=" ɪ��=�Uy"�>����!�a(1�HJ�Ɵ6Ъ��lDa�]��w�P�tx�`G��x�f�y�X��#êT
�������+�����&�B�SO���f���8��#~m�T|f+X�TdK���o�Ƿu+��Q#��"�������[[f#��֪l��X���@ N)c�Lr4"��ƄaLo��� 2�E%����(�e���q�'�s-p��7�ci��,��n��sd�q�g�풭�����7�����VЀr/w>�O�6�tn|w�P�#e�]kN��')� iZR�ZG�9�g�~�`̻� 9������juI�+Rrʃ3ҼecEij
cŀ���H�1��J�*g���uͰu%��x]U�6��-r�a���6��zex���ï�жdXq��v�q�v��:q�Ͽ�~jC�|�X��Q��|��,U� ��>����2�Wz�O����.�\�F��QA[��!�vR�J��v������j���Y̊�Ӄ��в���u�`��9?]("�GN*��P\���rrIᰅ��Y;�˂�k��m�G�Z�L�x��Z�� ���=�陡%v��un��>��Mk;��E�q[�"� �2ѵ�˂�Dں��Q�VP�q��.��E�&�ȠSML�	y��n��s���"U�&f�8
���}�:�^\c
��\�+9UL7����cn�^^7���}K�k(��*���zl]6��8�]y�7��~ݥ/p���A��@W���y��:�0ΟC���T��=�dk�**�Q�~�L1����n(��ƃqK��tެ�Y��T��e�0�JU��Jy����H�ɷkL4Hk��o�1����к���Xm���-�8�0��	L�?S���2��8�ק"Q�B���#�$��n]��)$R;��{}l�8N�FbR�!렓D�\��%ȆK��`#a��6oy!��"M�.�h_�f��� ��\r�&�t���;�`K8u����x$q/��<�}J����L�1lJ�����ԱP]�Ť�5�Ϊ�h��Yn�Eo�=\�Í�F��1�*凿e�ч6��ƜY�v��W�U�Ϭ�z�i/ٰ6%��f�9un��>�s�nm�����p&�%�tڶ�Zg��b|�N�|���.p��������HJ.J�����ob9�����
�jb�#K�rKҿ��ab�m�>�=��e˩��,j"/ ���3G�dUx����0����ۼ�9�7�><�v�_v����*י-� W�����X=�/+������fh��O��3�tr��ޏ���j��E����A�S{W����a��ن�^�9��om���^4�Pj%@Ӳ3a�U���ߋ�ƨ@�Ywr�><Ue�qwvɮF����E�ѳ����S>�쨾p���p/3��v[���ib={�˜�W���?�c2�8Ы�˗��qo?��:������I����v�
� _�s�`X��3����Q���"iG:���0b�w�`&F�ρ^������w,�V7큸��%|�"�Ƶ ޒ�"D���X���`:��V�4�ﱫ�=8:�9�pW0I��8(w��:�vNh�caRk+%�b����H��~��/}��,hb�e
�)�Ng��H=���7�;���`��"!�U
��G�~L=��O3�Ԭ+>b^o"��o�%�ù�1�@U�O��(M��H�U�cW8���Gɂw	 ��q����S�����]��/~e��
��Hc����-����!i���'���-�v~��+�˔+zlGi��xU�r��ػ�K�$$��l~}aK�0p��N�R-�����Z�A/D�1����6�K\�<�ţ�'��w�Jg��K�Ev��:X"��9�9�z�.R���Z�V���o�눹�������nh'��2r~���]����Cb��q|do��1���$˖�\y�dHצ���ػ(d�u�t*��~zcCt��d�С�LP?��̙G�e1�(�A�}��ga�h�oðk
�x.nQ+���L�����C���&��0�
�N����V��������S;��r�	c�u�쩡�P���"Q����lm24g��gsv_��,���?�Ô��<�o%�����ť��6���{xr�ѵD�X�����%F#�Zepx�#2���$�NZ�IX�e5�lIn.8���=b*���M*o/���0]�lY)�rG�d���*�4�-�G��o��\�4l�ګ�y���T���.��+<�A���K?��r��'� к��/ �W�^~�@����^��Ew�ZG0J�;����"Uh=���4��;�!?0�8ҴO��4M����i��7фG���ڲ�˭����Z�D�m�b��څ'0�*��ÍrЇpк�hR���_vg@�4�WA�x-Ƴ�Ѕ�~*evf��?��k�0�(�<͒�8�"*��~�S x �zil����,�=���!x�:��;��,r`�s�AD6g��@���{gT�}�ʪ�;�w4��4����|=��]�ƵW�����i�͇ͨR��7�?$�%�v��$�5'!��q,�m�d-w��ͨ`�&��QS�g�y������½⇦�w����	V[Ϧ,؋͌l�|����_\��sl��L6P���S��s�&�T&&����T����l7�>K;�+�#O1����-(	����Q�*���p?���؁��>��^�ֈ�ȳJ�|�ĄkV�)���\0aD�$�o�~!C4�zSf�9j�_���Oi�
�+���)��ڤ�P<$��}����9�������F��c#��L��m݇����A+�ݡ�iUeo!�u*P
��@Z���fl�"B���1 ����[ã�����PMU��m}0��:����kԮ2�م�֩�nf���@�F؃���8~��U��K�R�7ՙGoe(4�e���i�@��F�}�<�<�k�"'�@��;�ڰ:�!.\�ŝ�����Q�:$��x[Ur��&U9�$�Z�Y��A�����a)�#�]U�6\Dz}4&���a"1��Nu�&�`���Ŗ��w8���l��6w�^W�i�4V�h`G/V�&�_�L|�_R�M�[�[~dY��^n)�9 
$V��2-o;�T=U�P\h���c$Ԏ&��>	��PLo�fy�����9dl��Bٙ�z���4C1u��e� {{���jNITL�t��IP�o��F�� S���5h�^��0U.�G��&-��A�~TM�Z�f'W�P��*d��_�mH~�1��w�e�l_O���S0_FI'{u^D���0���H�k��ي7r����
��>N<}H�Q$�<�n�[|p�__�H���y �MҞ�r���z��A�ˮu|���k>�̥��fZ�`@��N̼����~V��7�W����ʿ����	�O2ãގ���f�T�@������j�;��y�Q��4X&�MZ��#����Ӊ:��:��Z�o-������ s�pYw���&5��I�RM��������|�����H0�V(n��n��:Z�E�lRǆ^�7 /`�e|�*0��0�eI����qڽN���uÞ�#W�	���G�
/i��h�2���vè���о��Ծl�7a5A���D�P�
ZP��W �}-i��hA�̪�042��e��k+�ɬ}Q��|\p�4.\�aֿ'����$4��&9�GAsL�A�ʹ�QK��BZ�B������ȴ.�z^��1��;^��	k����⫼��i��J�m�`�ڛ�~�bM/]c)��ջӒ� �	��;�X��L��=.�Lt���pK��;�I�L��l���bu��{��LcK�A-��|Sx0�^NJ�×1����\!R�j-�P�X�)M�P��:X�o�1tOXh>)3,� $��45X<�m���h�k�Qvy��ԛ��\�~�^m��3X��6�t]���Vn�����YUT��1/�?�n���2�~eׂ�Lj����=�}-��ʯ6�~��[��3� ۔�����R��������e��V\u�� 2��͕�߼Z$%m�L�KR�c�Q�(��y���Qv�'eG;>bc�>�ˇu�s�4+�����������{�)+�P����Ϸ�W����έ�z���>A�6��պaGd��@���oj�^���0<	M����(�����3��I����k毜1-�z����G��~S/�/��տo�N8���χ�x�ƪۈ�|��r8�	=ܚ��	���4��c&��p[�ZX���k�ў���e^F���	����v�6��6:��[yFl���:�A��F
N~EC�I��uz�ݛ�<���a�-��.^<o��/�u�{Ӥ�u���So��Ŕ��F޸�AR�z	1������S5��IīV������k ��4���!�����AEe>��[���p#h�/w�q�����2��M���ot��;ǌיpD�>���\d�ϙ�&�o�LS*K�WX� �t1�-�3u&�w�Z�5�Pt���.?u-+-����W�E�	zT�Ei�R3FD9;	���/_eHx�+5F�-��!��,r��p��<�p����3h2��E�>���34i��a�ݥcTY�o���������������=n.��/["�E�I��jR5�kÚ+�{��^�p�CŖW\d�v�[�k�,��BmRR��-�qҸ�����c�cUچ��ͱ�
{�L���:��
c�'����\��	ʸ��������^���o�G% ���O�5E9E��z�	�������^ ����d��~�1�m͑�X�[�p
SXb�]�4�
��
��&����d�y�(����
q�����aU.I�S/i�5��G6��**�G2>�M/񝆆Tf���Gd���X���#��yxz2Z���h�� ��g�Ȥ�_0��LiH�`��yV��[5k�A�;[��e�G@�e�2A��F��_�M\c�B����y�TEF�a�ڏ�UB~n�����c�����2Ŷ
vd�R�H"i�]�`�`��ۓA$�rs����o�P����x���L�|��^��4Q��d��f�!���aVY��	oዖ�n�}����~A��-�28*e�U{͑��TZ��sKnB���r=���Fw����7������.��!1�k����a6]������,�R��9+B�p�;�ޫ̵?���e��K�Q+w�]j��W�ff���i��3j׭R�+������%֮���?�W���}��.��T�Pa�&u��8�4J ��u����sF��u�p⛃T�t9�Bb�Kc)�7IY�bpﻧ�Gsh"��٫S���S����.꟟�k��kAI��G�]� YK��U�a���lO%L�����^ȷӤ`��� eo��֩�M�D��H<?���J������dA��6�nM�XYe��@,s���J���+����ߘ�E ���Q�sRM䖜c��Ŀs�y�J@�l�'#�fR�|�h����S�����Δ�k�7aI�����EA��b�ΰ��y��=U����;p�^Sdh�RQ~!��CK��K��_xv���)x.��)p�%<�}c��"���Z9�+y�E�R�1&S�<{������o�����)��[��tkSŽ	l쀛$��w(w~}�C�����ר1��Ѣ�ߘ���)&׵L'Ғ<�7YU���i-�� c��'DPT�E�u�s���X!���VO���^|��,Ja��g�D�ׇW�XV��O�Y%M�!}A\���6�����QF��[�=�ա��q"�o�D�hn�?�[�Y��/��`�w����&�0��- ��M�'�L��Ė����:�^�4d����ʼr��b�Ԅ`C���Yu� ��K��ޖ��M@��ܾ����}]u�7�LvU�IjJ�J��<E���3����"�j�{� �����/A�o&}�Y C����-t��E�C�|���W$δ���]�EA��\�׺�ݯ�3.�cv5�����_=�|"�1.�B�N�(����C0WT~{���U��������=�T璈��+i�~ի��p^<���`�Fx=���?Nr5_?k�����<&F��m��f&&�Dk;���Hj{���?;����F�o�q��Չ^j~�H�7���"�Ͼ8dNs|/����<{��(���,��K���י�&�O�����g�=̦ا�ޒ+�Z��_��PO�9/���\]�����\�KgY ]3E#1x.V+E��hՏ!��yX�����5�?b'�L�+����o6�Ki@F�B�BB�W3y��Gj����Q���w�~��[}^#]�v�q�o.�����oxY���!w���m�4k�1�\���N�s�ȸ���Y&�y��Y&?�����NBߏ�k�|��8��R��ȧ4n�:�i�zm�Q}�LBR{� EE2�@?5p��������ne�t�t	�H�tJ�twIwݭHww�C#�t���� �}��ܳ���_��z{��y~��"���J.��9t��ܪ<M�1h���_��7�W��)}N^�'�^"��S����XCV��@
�hf�mKt���w��%�
t�w<���k����Dኊ�P@�\E�h����w�C}����n�ܟȌ�	��عg�$'&�&!�
� ��]�C�Ê�k+�VzI����{Y���c;0V1pQ�Y�*��˺�}�O^��e��!~VHL^�p��X�������� =nnF�"�\*H�l�/��̔�NEu���坔r��[�[âu��/MY�_����qTu����s����+r6�mG9���p��/a<�ņ�ey�G��\�2Ͷ砹�F�dfeJE��t��y�G	xbXvM�Aš��+η9&��/���~Ѹ/�����؍� z��g]�6G�< |��&���CQ��{_83�z΂4#rj�WR������և�N��ֳS�V<Q��[�5�*��F�f�U4��R� ��/ۃ����]�p �J+G��� �ڭtg���敬�w�T�]��T�yXU��5iM���Z�v�qg���vvs���Z���6n��4���}�>d��xx|�m�P~:\�TWK6��>iu���1�G�V2��c>���rj����S�����$�K>�%����
��0�Ŭ�0��qV������j�Rh�����M5�;vp��R��d(���a�b��1�5(����9n��Q�\x���X�?�l��$|r��
�S���H��}��n��j@}_Ǖ@����j��shLE�bl��|P΃S�ùW���(:H���*̰����rc	���X�d1S��9�vrr��gg��mtr˻�1�e�����Z&�"��f㾉IXA�F����p�ס�h�=L�D�Ґq%7v*���`�f7�b��=A��A�)	����ȇ}����u��������z��8�-�}����z�c�]�t�s���ͯ=��gP��r-�\�y�g���>�l�W���#W�v#Dߊdd.�;o��Fd��>��X�R��] ��|w������RPogi�����nz�lͽW'�`'O!(�+oφ|Y�`�N������p��2����T8u�Kǒ�qg�v�j�fT�@5�.��hkC~Q8g>	�t��w+���4V+���"(��p�����K�����Z���ϗ�p�����_���юe����`��eI �]�ar'Y���Fi��͈��i'bE���X��L7����Uۍc.�!�A�ĵd�g�q��-�"�*�|{qu��$���m/�t�c�s���=U#;��J@��Yp_��[�0q�1R���C R	�%y���9�kB�j�!��g�ǫ�	�١�bU
ǹe\���J�7UUy�tS�C�w=ϤwK���&�O��qC�U��R��\/��!e5�nB�9��YA����:���u����(bi}¤�U�hf�//��\]�cT�/�9Y�uh�,D�%!ͧ��h��_�tX��^���O!�A@��kղE��!�Ѥ>��#������z��T((��_�J�;_m�V�j�;{LZ<��`�t4���jXgv�C �b4U+UD�k��X�z��̷��<�.�&�K������CS�u��e��a�	�[q'��c��R&��1в��jEz�K�IK�ÿS�1F����}�)��;ͽ��c�mWx� �R�i�K�K|l�����^4?G�����F�F3�&��E�|���hd��J�w���I7M#���vxj,�m=, VTV�*:$�i�(��b���Mg��(@6X%�
���:����~�xz�ǹ�&2�� �_7�wx�����5��#�Cu8���o�;���g!��
;ɑ��ջ'	�J3����"�_�@9\���\���z|��<��W���u���k��U�����؁�t@���_\�N�~>m�3j���M�'��H��{���iyݻ��J@ %����p����=����'W�2w�I�V�)'�ws�'N�	��6�d�!�ќ�g�a����r��Ϋ��9�}�ޫ�&�w+Z;g�>��3j����K��;���J'j�OO����(-vP(~�^���g�@��/��t��0g3]�
����?ҳG��oo8�	G0��|��S���rMQ��s�6?��o⹆�&���p��@&X%����s��Xj�ߚk���G�r�Rb��x��e\d.<���xy��ý��"���t�^���Ûo�O�N��=��paK/ӽ؄~LV8�g1��U߷4�R�̈3�X{H.��o}�VjV6���Q�rP��O>�	�Z�>���/�b�x��ƞ�]4�W���/k�B�R�i�i��s��(v�_���܊��*�S�������seʰ]ֳ#�_?�CJDr�b�"h�8�Z����`GU\��֎P�G��=K�%j�L�@����?	>M������Nb�4]Ƴ��*R1�9.��؞��YM����_95�S�y5�b����~0�+T��ޞ7���nn6���1oO�5Ln6m!�C���N����j����'���&�=�����4��Lh�"n���U�5�<��A�<�g<Q��Q�e�V��~v7��o��ZTv�y���k�"}��^垆�ֳ�I�vaŴhl l����g�2ڋ5_vɁ��*��&�����Rf�؞i�.��\���p�i��!����㣋����U_+X�ޣ�X4�ިDB��'�Zh�z�����C�\����)��E��>v�wW�֏�u$t�M�<�F�'���!����(�l:�����cE_�׾SF���jK�X��Be��B���n���MB�ju�)j|?\U���i��묧�"]��)
��I�t�����u� x��k�/E6�@���C��ܨa'�{���N���z�� +����L��1�y��z�� ���>Q��Fk�ϧ+x}�쓹���A|C�:z����М�]pf�Y}�{��x���'��Ķ��c�2!�����w����8���
:�+m��\Hb<���M���4��{tb�����z�7��8�t.�xiɥ=TZ�2� ?�s�+��:2�8�s>��$�0GM�M��_ZSQ�k�e�"�ewX�G�r�r���!w�.�s-��.��j�^{/��ܸ��ʺ�֦�A$�V���r��4ܚ�BA��"��{E�U.4ȓ�F?/����S���A:���_�5ْ���<�-�jh.?'x)h��o��DV>9Zl+����^������1�� )4Z��3��l�/��*kz}�ʫ�=H�$���2��k�Y���%�N��;5�S�}�>�h/ �'��W=��űt-9 i+�ᇖ<�����W�q����NF�P/ �A�Do�=(�V�SK�SD�Gr��]�������������,=��Bk���Cz-j|�[)9�ۅ�}��:	G�CW��!��ˆ��*z�U��b�³<��َ�#�������Gq����Cip%_[�(R�]~	����V�
��*������#�R��p޷���Z������RO��{���0����.D�k]me�E�Fy�V_�e�"ŧz�����8�D@[��k�&lQ�����B�Z�����j'�aϿ�z�7y�MZ��5��*5�V���-<}�#����F>%}'�=ŏo98��8�	59�v�O�x�j�Dz�S��A�]Y�	{�T�7d�����g7��U�,���>���
�"�b�P�J�lLq"߆�i�UO�����M��h6����H�!���O*��U��ҲC{E�����������O�PU*�Ul�}�}G^jH��6��*���Hz�	��m�m{ 
\b_��k�u��_�:��b��=UTص>e �	<�\
w�vL��1�-0�h+>nK�l۸�^����ݱ;�|`@}0�C�!pnIk��9�st:�c��D�������D��1�K��QoK=�e�'���Ui��]$��Z�rI�)��z77���� U�!�{S�}d�l=�����`�E��.�����x��\q��I��B��9��w4nم��"K�v�淋f4\Ѫb��	A�q�_4��H���bO�l�Tᇗ�b�w\a::ܤ2�8mױ�^������+`+5��n��_[���jA�qh��
�I��E9�M0cJ`2��r��Ph� �V���Q3s�,w5������V/o�D�?yh����Ӿ_����-N�� ��U��r{8�Ŋ�A���Rg�ջ�>zA��(pew=x��.�"�{?cd&ǯa*ΰ�cnF���WTdd:�&��>��+*v�S�,���|����V�w�I�u�W ��\\�3ױP�$W�ݮhǧ#N�hl��7����^�A�����Q��eN4�Dϯ����Q�1��7���g�=����pyYb|9��d�@�5*n��<2���{JmIra�7�����u�hV��:٫����8$�B��O��+����N|/�˛w�I�%���e[�.�8��wj}�p.c�K�#�Z�Gl똞���O�ܵW�~p,�y���2%�e��a_�%}L��^�N��6�����"��S�t��Ϛ��JPd�|%9R�����ܼM�_p����Z( �@t��5S���k#Amh�Z�éB��ONI�`������K��a�<�H7��z�kQ��"���6"D$v"�h���8��K]���	�Y�w��&JV�=R�*�F7�@�lR����4�3O���R�]�ɋ��-��}]"���l�A�+���~9�O@�7�'�8�!��ٞ�V9���q2�+��u�m��n|��c�O�0J�w$鳑V�v������$>��|��H%�ܓa0����G6�2�.��͵��/�6���8�R`0vK��z/}t����X���ͣP?� ���䜀�m�n��ws-��|�� �h�݄bΝ���5�xw���o�Ll�6�L�4F�:@A}>�q<����לd̒�ٮ������s�g�cfF�Z��5�$Z���`� z�����vHr���!ad �w4�*��0��q�e#Z�z�r���y��|H��N���Q��=()�/�l�Ժ�n.����5x��p�H���i5}�C4S������qRR�M������VO!:��/丳�s�G����Q�g��\���k9f1�*�Z\��p�����w�<
���Y�R�f�n����C��_8��}ER�.<ݨˤ��F��{ٹZG�<�D^��P����@�8����:T��v��] ��Y���Y1Geg���X����X�����������p�1���E�
�}޼���wHA��p��C6�z~����槦)��2��>0�*�xy9�������g��'��C �)q�h/�sM1gc��b��q�֔H뇊z��,�~9���8R���w�6�<� /"wx{��g}�1��FY~�ta�ڶ��(�d&�dFm�_=�-�،Il�3뼻��J]_}�h�Tvp������K��kYXȽ�8'pl���Yu��w�Mfq�
pE�m^�/������3ǧǷԾ�t�-ѹh����S\NT�;R�U��&�����#%_�\��?�\�5*��{��aK(���G�ݳ9YVy��]�n4�Y�[82�跨��Z0��y�����i��p���t9�C47���p,4�����t��I�f#T:�e���]���6��Mjw�G�1f�Q!�Y���[:��J�̴�؝،���5IBZ�Ke�:X����PK�W��<��я�(d=&����|�	���A����������^���X���#��3�D~~�����>�Of^��9�|tHe{�Ff]���N[fLT(Z�}���S��C��X<�Qbr�8Z&6� �LT1�/nz�6�b���^��3�WR������4n_����Q��k��Z�1R����R-�7_R4��a�k1�[�t���ܼQ-�콈�ɺ�q����H���4��?
�F��s,6��r)EJǍ�c��%���J}�$e��bC~y1:̘��@#++�kYZ�Ǭ��tWgmҤiP���M5��1AO��-���6�ܧBt�0�\��N���U*>#m�#��4�B�����������Oͯ�R}�a�7[�D�晳���H^��M\��R��E0x;[�\ǣ��_v^�ʡ�[B�Vc��Qk����x)�B�m���5���)6���
 Ճ�]VcO�v��>��)��`[c�M}���h�D'��c��\�S�;���yQ��J�L\����]9{�b���.������ LQ���J`#����T�2�S�ͪی4�2&����I���H
<bI����������g%K��6Cʻܹ�a.��|K����"��7mf���7_�]��b�|�@E�F��XN�}���Ndca�l��|�I�r2�Tq����[$��؂��������:�QD�(��aS��UJ�d0����x�)#���6�DgGGd�*��bc���\���\j����N�+�2��ͣo(u���QI�;B|Rw&O�;D)yif�q��Xv�����|�U��~lp�"�(Q{"��ι�W�9d���ޓaX���h�O4xZ%��'�[Ǡ_��Z�_�Q1�c��w&g�/}�q�m`��q:d�ET���3s
+�_S��`�����D��l�$�˦ꐀ��%�%�e;�0aK_G'�IU�@\���"*QV޾��j�^Z�y硫*H�����c��:HhWEy��;�V��a��}SS���L����!�{M���5ؗ쟶6��{\�>@��A���{��_\f��]X��)�6�tU.֎>��<�Z6�2����D���ۼxR�O �������G�C(�o����
���.�T�T���cJL��E����������2?O�M�W�v�6��6����I�(����fW��ST�DV����vDs(�B���m��H�;?�~���0�?�t/�XEK�B�cn��?5��u�Fb@h��z%��a^n��� �NbM���w.u�\a4^����'<NNtg�UX�~
���� ��i�vh���D��E(�Fo�X-���}����m�c��b����4�]�D��W���2�~ t	��)aP�~M�$&�cܻ!��X�9���@q~|o��v:7��XI��QQ��$�u��B�C��{�]%|(D�q	�	M�D���gdt����b��{b�(k��K#b�f%�fL%x��8�=Փ�� ؽ��׮P��;��q�Y�Y������
�1�M�+�3+�I�gɲ�ʚ�����pō��P��?q��_Ứ��S����Y����<�8�_�0��Ud��I��<q�;R���d[�ލ��$�L�co���QbS�׀n��~T�8 �j��f~�3x��媈����B�Yd��m��Ѐ�;���j��K���v���дГ�(v� � :c�7��Ja���x4��c���s���r��hr��\�n '$%�y"��,��Ş�
�j+|�X]Z�kA�Z2w`��횞�φd:�1��w�7փ	�W0DZ%�B��\Y�\uo�p
p�b�.��#F46Ʀ_^1����5�T�����L��y�j�k���;6��h��� �#!����654���}�O:�F.S��on��G]����J�{e��cY��M$H�%~H����8���k�ÿ����̇�OsE^���\'�o�Y��/{���z#l�AH�FK.�F�@����;�@<�����a"�nĞ�z��ݣ���*<�>�F��=1���#�xVG��p�����@�`kg�Z|:�x�*���ݚ�u�#�2��hJ���GRÃ>����-k�����J��ȕ8�5굎�Bq�/����i������l�N�ۙ+(��:��^8�fi����c����]/�D<�=�%�A�3��xx{ܸ�KïE��B_�Wȑ���Kѷ�'w�_"��'>����ԧ-���q���T�{�����6o�$N�x���S��3��[���?z?��V{"����<a��u
�%��P;��-����ͩ�"�b��R?��w:�.S0�xD��.|��y�5���9$��~d��0�Dt��7�`���=�DW�j���r_D��-+�o���W ��H'tg�6��*���q����x%�!bܗz0Ƌ-+(��S�}��^�����O������	�H�?񆄦�$A~8�=�g��Vr�-K5�g�v�a����.d�����Gl/��!����ha}N?ڧ�b�vO�{���6yG�0�ׯoauS8��t���v�$���b6�Z<,�Tׅ�Ћ�'v@�L�^|���3��c�fFͪ4�_�����$�i5�*�c����ܘ�Оr��&��'p�p]45��EG�E�oB���GS��������%g6�1Me��,uC���A��[[�V��n��P��R�Б>��6��^lx���x�4wd���bSE{��� Z����)�I�`��풒
�i��A��撡t��BzM[��k�8�O3B�
[1����-]r�#W^��7<�u&��	�s|/߃��$���
��#����Q�OS�X�'<��	���~.��ne�CW@�&��p��9Z?=MM$�W��eo�$r��Z��x�)��v�wB��J���DVfk ��M(QM����4��7�𰳚~D��Y�,�Q�C�N���-���}���1�'����z��v��6��7Oo�Y��nԙU��48^'t�w5F.i����eq�b`v�s[�����>z�Y囅1��y��/�$���L�r��߇��W01�4�c����=����{ O�u���s�lT��|��-w�)w�R����W����=�ί��]q{u�|�C.��mf�ꪪ�/�|��(Xo/�w���.�(���{@�tu���`,5��r(x>�6os+7PWl���c��As����rM�M���ht�D������%0����I��h<�m�r��[��D����� @��Ha�-����\�VO����&o���ܸ�m�����֞k�5�Ã%߅��v��s�DH �
���W��R��y�Qn�D��g^:�uL����ԁ	�N. ��9�`Ү
/!@�zU��-�z��ORx:�u��ˬᔬp�73b
8��F�V�i��w@�%]W�t�ĭ���j���ÖO
6�L������������4���G�SU��\�|Y����%%&��ݮ<����lݯ\��r%XK����7�B���5��d�� J�����ᣌA���O{�=��#BMuhu$�u������Y�oǃ�N�1�MpFY��&��!�?��r'Z<���66��6������b�6��n#=&;�Vh}�c��7���#�������^��MUl��e�m|�@��3p��zT	�Ok�J�`�j�Â��{	�c��R��Q	��Z�Շ����^���b[��3���Z�3���U�(qD�i����/��n�s|��f����`���7���-ϋQ��;>����O�2_t/?|�#�A�U<]H�r��x~FF�`����	@m�C��+;���4��<�,w�����K�4C� JL�c�ɰ�'��h���d�P�FA!���X�'�rs�H����V�,)����DA%��Ǟ��?��-�f-�8~���"r����k�4x������r͸ ��u�2zhO�C3{���<eJ�Q����������h]�M�|[[q�i�nm���#�G�l�SjǍ�/�'t:)R���ZU�y�ڠ X�M"����W_ ��<c�.ta"��� �6�����t>��?we#���o>-̠��$�`����t���p�z�1�qc����
QLA]}d��)y~\�vQ�,Tڍ{�1`��5�FoŤQW����ɗ�(�����,�++0cGC ��q�?[�:��@�p��V��	)"8�G��vC�u�n�7a/^D�Lq��{PdՑFfA�bw�X�#��)1e&�)���k�^[BZ��9&y��7�fK���zS�z6SEU���P�8y��t��C�����Ot��nE�{KJ����g/�%\0BԆ�n�%^G]/L�oR8�6�Ղ�c���8'�^V�m�3]_����xȮˮ-_%C4��G�?9-��.ex:f�$�E�����I�ӽ��'�"Cjh��b���l	u���ơʖ�ߖM�;O�W��u��!��R���m$"�愒�����N�*�.�����
81�6����s���1�gΨ/�Z?�5Ppft�y8�.7�uf�L@�?��آ0��e��щ��i_���,;{�J��&���m���mo\ß��E>�k�3����	���ʄ�oR�pu1h%9nv3�2x���bU��Ȳ*�O���H�������Q� F�3]2���{�G7%�G�n�}_����!}���7[ҭ
_���<��ͫ2kƱ��' �$<�Ez�7O�D?�g��eO0��:���@������������~o�J��I.��Fi��)1���'�2:!O���BHI�I��y�7�q��A��P���� f�{�m���~�^��@V;��T�P;����i�v�u:��:o$�@�ة�Os��S`%+c�w}7e3����zg�.��i�/�&Ae3.I���#ɹ��C���t��	�4A� ����_C;)}�sA��[��Mo=-[�Q�~��>͟fn��������Ө>��g;�t��n�H��+���תw�2�W9)�&����/�$�,T������Tܹ*�;g\ٜ�:]հ�|u0K�ġ�H�2��8�w�ة)4&u�����vgC����M;C'Q͌%�B{a��q�5&�nD�Ж��/�i��+�ؔ��=ժ����˩Ww�4�w0J��2�Vޕ�>���_2��6=U|b��~௱?��Y�9�_۰�q�q�C��\`�h��D���ZJs~���Ps(j&�kV��b��|���H��>��0��R|�^��?{.L�,�^"W�D�eW*~��DP�^�#��GX�Hc
��5b����&����R)���C��,woԑ����v�n����M��X3���:26���U��<�������L�������X�G��E,����k<��!����@�!�����Ī솵j�f�f���s�T#}T�㰅��rHu��D���3���~_h~�����K�r_,���С���$�X��P#����3^_��i����UO�|	�%/��vt��E�U����.�y�C�B�q���%ʥ.|��g7@�
/ޙC��p����WP�?�P�h��������Vr��	񪣝V I
���T��e�M��`tBL��kl�3��r9Ӷ�Q���&���@\w*����*H�+�i�����#�$��˂���W�(��:UT4ȼX�ݨ�V*M;��B�hF|��0S�*U��ഘs�_)�*�� ��v��]6��^}�+�����SK�n�Ɣ�dE�nc�e\++"��C'@A�� m:R���[**Jm�.8+�i'��B��X����Xk��_u�AO����8m9���W�Z�5��K���V<L���q��n�m����v��'�G�.�"W��2�"|h�Wj�F�:	�QS:)�@�t�����2B����o�j�A����7Ƨ'�f�,��j�at�B@�ƨ�.D"�H[N�<"��b�����_6�o�����HF�u�m��P�4G�fBo���NJ\�hH�Ѕ����RZ�G��/֦�����5���o:P)$}"����wzE�rQ���!�1�$�?�/v痁R2�+�A^��[?�X��[�R���܁s��R$��e�@�T�kl�5RH_�H8�/[�����âV�M �E|� v޶����5�7��Y���e�؆܀��*��QA���͆�i���W�4d`m%)	|���p��J5:�y�Ý[��-��d+pss�S�"��s���_U#2i�}�!���Z�w)�ncM�[�})p��>�-4kB��	79�Fj�R�1��>uu��iO"�-|&{Z��ɼ�q�n�[��R����8Q Vl�J����W��^�B)������vLת�Y��P'�Y��!�4��agu2%���[�SGg\d\t"�Ҫ|@��l�tR|Q�Yx"crk�㏅s��A��Adm\.щ��M�L�Y��d��Xq��7��G���rC�04KB�r7�J�5�� ��Ù���T��%��ͳ�����m
��c�
�`�k煳G�����
���9U�kVvW�z��e�1�*�q���[SWS�� b�8u��(˾�-�gx��H�\껯s�z�.��%��%�y<xѥn3������*c���htd��~��Dp��=� ���Ϳ�P�h��j��"��Y|{���������X������ߵ5$݁ӥ�A�vQO�X�ѫ�M��Vht63�U�L^z��(��#9�s�p;?}v:�P4����9��ue)���t.�6�{~a�.H�X�DW${�	����]C�����~�Щu�Րُk�n���{|��C `�85;*U��{:��������^oC�yu������L���nz R��.�����Dp��}��y�Ի��s柅��:J"q�J@�L X�h4s;g�����B�0�#uS3p����Cߦ_f�]L����U���5ޯc�֊Q������RחS�)gz/��<�%�rC�uW�@�67�_SnQ�	����� '���f� Mq�!���-�,�vje�1?J�\�) �{�RlT��J��}	%��[,��<O�P���CQ��R�k�S��_�yV�o��V��ndQ��}s��2��F4VCP`�X[>5}w��b.HNq�H�5;aZUE���uvƋ�J)���VS�ٿ�����#9tw� 1V�48(5��ʒ�k� ;�]x	��;~�2[�D=��p���Wt��V�!)��ÎX]���K/`4xee]	-��ޒB�X������}�☚��S6�%p�Eg;C�;��hڛ9D�^�]���[Y�u��G�&%���� �F"��KV�N�Շ�6����2�L��{���9��k�]۸@�eTJ���t4��X�5]����_�:�������#�[�u�5��u��|��b�l��S�,f����6}�1�y��k���"�OG⺭�����sD�	��U��	�e�GY=H��VK�KN!؊�e�`�/2���.mU�Ψ_|�Y�CO�"�����po�w�Y�9z+/�Y��	�u��%�6��W���:���=_6��K,"O>=�;?�%S�l��C�55wsס����V��0 ���T�k'Eaq��rb[ݗ+���"�X���ԩ�0R��� .�5���d�֏`���/@^�׽.���;��	�T5�w$�/Q�[v�����a<��������:ܪh������|{����{�{���Q�<��ʫm�>.�Su�ѐ�Z�����Bb�+")Bn
��t}�,$;S�F���<��-:C�~�1�i"����k4��{iJ3���#&�9M�Y?d"3EyF[k�.o*��K��4�ڹ�Mu~��=�}�G�'�|�#��Dd&��Q��1V%C+��!���kBp��w�ۮr�\��!:#A+�F��H��F�*���9f�cy������{9c�C�>�nj�l����6'��C��N_��;��*c�I��g�ʏ�So�����V��K�a����,����`��[0]mᏋ���a�*���;/k����j����S�'Ɯ��ҪՁ�c6�h�?}�4��P�?t�`�T�<��%��s;�G�稓�]�R.�u��HK�ew?A��WT���;) �x�_u?W"���q�IU�Cc�k�T�X�8�+��11��F&3�X�!��ɝQ�Ķг�*�I?�<�X�8���82]��g#�_~=~d3f`��Nϵ:����JU́7�4H�~4�9���~������ut�ѐ�)�_2{;�v/��TJp��ewoI��ބJ�IH�L䑥�wu�w�@O2bU�������f��4E�@�֮ڪ���iw%ü��8`��k1�
��"��/�825C�쌷�g�����]*����榭-�Դ�
�Mj����x�D��=�M8h��Yr51�%eD�:��k�OT�6S����ގ&�l}m����[�i����,}��IĈ�Z0˃Ǜ5�o�����!׵LԷ�::-���]�NXȫ
U5���y�ک`T��B�c�T����HL�2�"�Ø���(R��ؘ�*&ɘ����l��S�{m���tn��o�}�.?e�8Z~�S�ӝ��.gl�0�J	tl�k��F7bZ=O��v�2����E�u<1kr�4�݊u�Up�ţ����Hi:{2/gw��۽y���i�\�g���JH�+�Vk[Q���q�빼�ʶ\=F�c�Z�7s���?���;:��`�/�H���e}���8������fm���tm��'�I��?:���?C�l_ۉ.��~��#�7Y��^�|���f����

;Oz�k���>3�FO����
o(����Q�Q>H��Z�B.��5�Y5�xh��ړM?6q�9A[��A(�j��l��w�����!�u����E6y4�&�]p�r�u������8v7>:�&��]�&I�X�/���eU�͆�	��v��8}=�4��NY�jy��Qx	Q���=�b&C;D����2]���ã��w��s��	Ŷ�2��A<$�#"4|ʨTĀrlY�O�}K�nA���{g`���4Ҩlho�2�ĄoJI�Uݰ7�|}�]/��kր����t��`��cPW���|�����H�/��_��#979�4iQ�oB��
d���ج.����>y�C7���|�0?jq�b�C��f����^�WWΛ�)�-�M��$*�t��e��y�h�щ~�BF�GqZ�22J#�д��i1�%R�L$��-\;^�]�0Y�rw������D+�$y�� a�5u�x�J��'�̰"(�*��¯��?8�1� �s|1�#ZFb�3F'�WE\	��3%�b�nZ	34|�c�c���-o
?�3���6em��1���~r�8��ws�ğ���!�=fR���Fy7dUQۄV��jj���$��u!�]=��u���j�߳*d��,Wq�p
����?�)k9����3���P+VM+���yW
ʝ�ڟ���\&R?��Fg�xq=}P��A.�G�~Za@I�I��eF���w�9iAO][bZ�뫋�j6E���P�^}��Ԇ(��FWU2�	;�������Wx;��<�u08wT�&��[��9J�nK���qu��f��"�DT5n=bq��F|�{�ʎ����9[��������V�O�5�q(�h`�0<�s/���&��U{O&QUm���������?�C�=��P��ض|,�i)��B���r���n��;��)�sI�@�95��'�2�����V��o?���}C��˸z#����t��*#����EsEum*��-��Т�/�6},�Ф꾂�d,fw������z�=�oI*"��ZQ8�/W(��z�6���WZ��7�3A���9!*s^{|SH�Ɗ�6懾�P_+�����v�/��e�Ч�]��lm+�l���H��������sL~�ږ5��8k�ʧ���x�&��Ǵ;��j��%q�{S�z�}�^=ƈ�{��þ�v0$rK��>�`c]�d��=PpyRorIA�H"��xE�<{�8lmpaԘKZ1���Ò���7���!?��Xv�'�m��8�ra����]Ci�{�5���!xF��h���C�o�9�#����὾�&��SG~� ��]��o�<I!j�d��ƶ�27��5r��M�)��Վ�mw��U8Q��t�6�I��mo�hl���?,i���塢���: �53�>A�����UYХX��֞���[$�%��(%��Dptu���l_����`I�z]�������G%�װ���'���(�з�n�.��w@f^��M��J7O?��P+E�ͪ�ށ7������]U�{x����T�q50���?ߌ��7���R1 ��_�k�����u7��gg����w��u)�u�'������F<
�ɽ�^C+y���=���/�<7���3��'��G�"ޏh�mϘ�����3��� �]�ws�����`˗�%#���h�|��h���oH����&@(���E?��x��|)!��/�ힻu�Ƞ�k���`&�E�|ؔrT��s����Y'�{5�XP�����5�?��ٍE��[��P�-�z�\��z��"�;�OO'e��%Q@�x��G��q��	1������ ��vs��t�*��?�I=l����G��KUN���ѵq8x�1���ٻS�p�ue��d���Ǉ˴�Tb<0�-=:�ϥMy?u�LI9��rQ�]�S~qi�T�Oށk��c�����Z��6�k�w�]���^�t���t������]R�҂t7�#G��Rҥ��R�Q����h�6`�h��}���?��08�����+��\���\������HO��B!nU�T��f�b�^�,J�|�,�����y!R4�;��\��t�|Sb�gKK"ы�<�*��à���
S�Am��.��^tn	�	�}�x"~G%-;WP�T�B�60<;�(�ₑk�Ґ���C���+Q��`���o)�1�{Aj_ X~�p�^a��ѓfAt�N�=_�@"5va�j6""W1�g�hw�j�}�t?O�������������$�S2fw-.H�ԙ�f�e�)N��<`n�%��1��kl11�8����m�ȭu�Ģ��N�; j��i��J�I�	%�vR���P"�	�G#�;�Z��+���pڌB���6�{�$�d���O��
�<��q��-���D���, ߢ���ߩ�]_*D��o�L�7�eM��a��bce�~�ѡ;ڥ��i�u����-Fܖ���|�,<�ݴ��9���I�&����ڳ�(2�[`yr�Pե�#��:j���$wi/�1/�
�[��(���~�/dj1RY�S��W0��\ȧ����	��Ȗh���╺( h���`�_!��TO�c�&��\��=/�W��Ő��sct�[��`傴���˸LMO���U�Η�8)m+�[��p�s�@��k궷�9�-d���Dsr@�F&c�;}e�r{��<�H�os0;�q�K7�}e��W}�t7�͵�SW�P[�=i�64�ͭZ�.|qV[,Kɸ�Ɓ'��1�6�C����3�?61r=�p�v~���H�[=Vb|M�����B���P�U>şw����:=���)��xr��^Ѐi}M�u�L�L�P��R.E��s_X�on��*yK2a�r+��yە�6�~��OB[O>Fh����_�K-TH4Y�_��#�Jj�B�[ԭg������o�L�|�.���8���>����D�����W�B��x�0�1�r�}�p�d�>�L_�y)lgf���z������i�%.�H�@c��gR�x�8��c�L��ss�#���0�����e�^~���E�pK7��ԃ/�i�T{z�Ф߼19f�U����mG�?L�U%�E���4�L2���	$6��l(�p�QB�����{.�A�Q��ϖ�����&/���H4��^��8�;�b ��25F�7���׾`ߗ�W�pb�b�k�-��Ƥ��&q&`�Xk�Ky��2�����N���N'�S�,{�Un'|�q�o��S��I�/Kk��^m�R~�Ad.��wL���f�v݆��a��5�G��ľo�%�9�v��6M�"�i�A�e_�}��;K ��8�{_d��IO`�K��?O,����6�v�P�ЙYۙ���XY��īi<EFh�5K��FwG�gJ�G|���&3M���~P�[qW��g�g!�D�����uO*u�2�:|�_c���3�ٻ;3k-~;X��6l�C�5H$��#D��iwO�����.�
����:��~h���6N#� ���y:��$�����G㑛�d��d1Z�ۿ^�������ԓ@C�͆/�L>�\�0�^�@�D^�7�]��RM��R��2�Y����X2AV�o�(�:��߼!B3�zT'Mf�V�g�����lp�7},��m�U3��}o�EY�"�<�ɚ���0�D��b���43��q1v�
j�B���Ŋe�Y(.�:�ѧ��q���̌M�b!���~�f����������w�'��Q�����:|��� ��`�?n�&�OV�������T'��4��6��陥e�_`�Ӊb˷��ޗy�\dBs��%�]�1�4gb�-�Ğ�M���">�'2}ss�� - �#�R���F��sb�0�=L��4�pW��s�q���.�m�:�����)�3�_��u_��);�m�n�xL��N�WM�l��$A��֝4I]lH����$������%�1�-�"��3�})�h8��6����Y�^VP�nN��?���̫��%��u�#�K��F�@dt��1�=�.Ҋr���Y"<Tw���eK"6K���� &�]J<��_��&Dk��Jk.0nPc���4)�&�G��x]��գ��!�5�H��͠�(�nq���M�����`�v����r��+�8{*o��l���o���C��)�xy��s9�t�`�[���3��a���;>A���4n!�MQj���}8%>�M�`����b���f��*d-�Ւ��k{^�󌘏tn"�ڂ���:r2�3�����&�Ut1��0�����y�t;�/��'��m�k��@�V׈����=�F��fB�#ܣ˫p{��A�YAэ�|p�ո��3gBk� �
qAwg:ohȪ���B���knc����H����1^�{�]�z�c��x�����������iy&2z�ޗ�'�N]�6�l��~8V3h�S�S�?�n-�]:��Y_/.��U�Љӳ� 
�54	~�(}�����/�G`��[BB�Ĥ�e=�Nb�/I���&5�0��>��7��'"�W�l���f=q�L�	�R����+_��gBP:5���>��u�
�'�+��6���0!c��:�R!��{�v^R�C�%>Y��j�s�[.��?��3 `a52U�ͽ������C�2�#�n���9�Z�B>����~@���;���(bJ=7?(M���ɽ�gG��_����i���	��r#}Q��3�r?���	�� ;a�X��'�?�# ּo4r�)��C^i�'н�>hx�G��&o��w&�>)&3�0>r;Un09�&CT�d���;�A�y�j��de�����X�p25��� ��y�3�X(�zf�\\��Li��vW�,f�ɇ��"��	��;�I�!�>�(?{����h�n���7ί��_��&���R[��|i���^�:�:�Fz�yl�뷙��>�����+&t~�X��A�^��Z�,�1�,=uu!i����IC�PE�0ZR=;�a5�;�{Y�U9�Uu婭{{�� ��5��:$�Z���9眜���ۏ��ŝhɮ�\IV�g�K��(*)V�5�x�:J㕫͈����仟���K�N,'�\�1���t�GD�	'������t핳JA�e~Xk����Y(��?E\���i�<.?}u��a�i����#{1A]8""x�Z���!��4�Xv�����/�Y�E�t"���ڴ��FyӿL)�!�0����&��C>f�J�����
���~Q�c��FMͳ����#FӴ�kŹ��5p�W���k������~��n�zC����/� �m}@�H������+9@�bJtJ���C����4~���:�3��A���2Sӳ�`U���4�`�}���j���4�p�� �T��6'�o}~�_��
�?m��@�/&T���>�C~� &�Q�����p2RzΗ<��r�Ҹ�dT>;ӝ�w�d��S4��	k]�������^"�
��O�T��p������@�c21&Hij�`�O�C9���[��ɓU��w�֓�=���'�7�Y@pr�X�#�lf'ԽS����M��u'�V�Ե�>'r[8�a	�~��³����I���x��
,�{�w�h��QU�1���T��d�u���������rw��Z� knǤN^�j|1�+0�K������|���/t2r�k��q���v�e�#��o��M�ɣs�hV�c�8����Bơ��$���t�D`�|푡�v��/�3�_K�!��_��_������;������nM��
����+Ա-��!ܮ+���~�w�������Nl(�I�������j�o^&�h�Qj����ӟ�ڦ���E�/��ƑNCi/E���:��N���7�i�h2���M��������Ϯ}�U��}������B��-�ƺ;ᰕ]W� v�2u�q�n������l��p��f�#��:P0�}Q�D� �^}t�duN-��{j��R!
���`2)��"�?ow_u��-랿	����\�V_�j�Qv�����4z�5.���j��OqU�Z^�4�x~�ߨ���@e�7����E���汀��3�Y��&��Ny,NbF�i�^O/�%P�\v��i�����O���h*�����!6��0�h��,�3�Yf%��jhA�F>L�M\_�'g'�=��f8y$=���Vq�zM�0�X@�p)��������2@]u�"���lI��߲�I�ǰG�P�P�[�Ak����K����m]���z\k1���������V��V��}���g�r�l��O����p~�TJ�c�����R����
u���C �����Kxb��U��;�T�g��C���P�]��ü�x��+�rI��D�A�Ң�r��G+������;0j#%�R�d'\�^��ĕ��Žv�w\�i�m�Ǻܚ�N"�^τ�ȳ��1�o��v������XD&3x��:�S+*ذ��zD�:��r�䎓Yڊ��ҷQ\�ʛ֊&~�2�L\���<��8xlS:ʛ+[�L<ώ�(Tl�Ї?�#��231*��5�bf?<���̧��pw�s�����s��GS���w~,�n������uu�ș���39B��t
�['<����x�22�V�蠗m�����H�2�i+��Y�X�.��=P�	Q?�k\zay�47���կ�a(�X���z���+�'���_����4�:EfVA�[��	ғ¢��Do٧K��������C\2p�gh��?�`ݱ3��1܍-�ƵyM_1����.��-�-����բ��^��E���uD��ɿ������׏������v���"]r8�G�U�lI*W�2)L�w�Cj�w�r�.�
�,�]�V;�i�m��`^���S�(�#U���Ԅ\~������,S�E�5�QRI��*���cpٷ�8��օ�@+B�:ю�G�@��6
�91�w6�P�T��:�0s�-��~{�[��/�=ezx\�����)��苮�]��� ����zP��g�����b�^��׶��7���CN�h��?��kP���3�)
�m��7�י��_�0Z���{��,ʻ�~�4��o��9u^J9�Iʼ1e�b��=72�$�9#��@%��J�p��m�yQ.��p-͵�$���cU6DP�䴳�6!m	�/�P�p�Ѓ�!k]ｙK��+8b�P8\����q�as�l"1C�3�"����_w�J1;�O��r��[�2i����)"d�2ˏ��ù�d[C��X�N�*a̲gz�����!��`�|0c�R	
��E�H�BA��[�)����_��pW���i�i�G������7Z.n�p{����*�:VrmY��;Tß�p4� 2�"�w����x6�?2��V�R�l,/0m�mR5�c�A����bzZ�r��I� �5V��{d�zk�g�:&'�P9)EB����,�����m��s&vaH�Jo�y��x��1r�v}�˾IM�_`�oon����K��=�<㳫�lP5-��b������y�>JM���U�y�p�
�Nq=��t���}�b?�12BQ��K1�_�S�z`�䭾ė-
6{YD������DDFr9�<�����ۚ��2�3N[-�
��y��lp���z`���>��������&�q��}�"�oo���0	�F���!���K�hн<����a�f�yRH_�#g�R�y�ᗶ(�WI���ak"�Yj���U�̊���5l��xa}��sGq>Jih}�g��XZ�\��@��T�������8�2��4��G�O����w\����{�퉏�?���#��@`B�����EO���Fmˤ�������<͚�̺֚܆��_�fqI�D��X�:�:�����!�U��p3J@J�4���8=}ID����
��kp�@���]�]蚖P�iȵ���lk�� �l��5ؖß	�F)���О/�4��qQq{!���A F�7��NyU>s�������Q���[U�{���1��r��n.Sҝ>����_Tha�����x[���=�-�X����{�*�3�Q�t���_Z���I@���#�9��g\ɘ:�Nj6=	��z�$�� ��_��#�@B�l�­���ą#�U��=NZbݚ����d/��q�^J�G ��H�z�7n|p}]d������@q��T��8�%�g���3U%��a�����2�66��Α�!��
��k]��;G�5.Q�aIZ|-EM��Kv��$p�:/���cĂ�V�N�Ϲ��hO_�~͇ç��)3ۇ��[#�8�G�?��\x�ɥ�VFe����c_��̆�z)�>%�ft�+ƀw�*�pޚ����E\ѿ�c�!�̍�
�F�^��?��U f#ļ>7f�0�>���bL?�*�nt&]�m�/j����S����2�����L:��tv�Y�����R?>�娙Å�p���
���,V^r�\��:�0&ms[�o���0:"�~��]�DZ#�;F�?�>_s�����}c����@j���U�
H�5�,9���E	@K(࢖=<��'rW���������3Y����]���Z��Ci��s
��V���0�
>��3o�@AB.�̘0��zȭ�R�	U�Q,��?��)�����//`��D|b��r���q\ǡ4�`uz�%�rvM}J�C8J���!�I�/��H
N��"��VS\�,B��.�'��?`�������!J9���[���������2(>��=��*�û��On���nF��O���Ι�ǁ���t�<O�ǉ�v���8�'"���2n{�c]��?	�<�jq��/�A��k	���5.�B
tŭ <�}���x�[:G��.A�6n����7!ۆ��z&�+���(��m���_�s��nv���e饥 ?�S؏�-;W��*���	��ݑ-�o$A�t)�H^�Mr���3Ǆ��.����d
���\q��{�Y��~VH*w(QRH�̐3	Σ�R*Cz<�j�Z�PG6,t���5�����L�ۀ /9�̫� �f�F=���&ִ�}Ӹ���G�ZLr���qC���/JE���c����nw^�����J�s�g6�B^��ٽj�Y�=�Xe��߅�ͻ�n�d�>,�3	�
�
��2��o��]���<���q{鴕W]�豠`�?�ڕ��,!uҠ�LN9G�1ϡHnN�eJ�tw	F6�d�3C����m6������>��sE��*���͚	�9�E=���
�`�Zf)i���_ /1;]Z�l+����i�%�m��S2s4�ϙ Z�X���2u=����ъ����10߅�c�C��F����GF�?� KV�G��7zS�S:[����j��ǁ�ͥO��.������
cv�U^46��0#��)p����;Rud�d�/����f��Y}���5�����b\�x�L��*b�R R��������g!$f��A�?h=$G���^4��_<&�в��h�����h�T�3�M���?D��|�]\���`=�4�f���):B�B{c����st�1!b|�!���,α�KZoޞ�M�����7~�e2h�I�!�W�Z/�p��T6�Z�r�fػ��z�_'��uӶ\�_�[�R�B.��|	C�3�]ʚY�qN`��	)O�G�]s�qf�]F'r������.1&�@=Y��W֟���=]v�"�!1�?�m�^]��UG��oE�k3�ڔ�kQ��_��h�i��L&�d�+鱨�Y���qe���'f7}�k���I�	q0���]�����A��ߎӤY6��*�Id����ؠ���h��\3_A�{eJ��eUFh��<%j�+j���D⫑g�&��E����9����ӆ}g���(�7Dr]Xb���<棳�	��ԫ�Q���Je�%ÊW���+��8��CDL�i��6W{�l,�gm�Y���i3BW��8k��m�<��ql��qc�F�YV���${s�}���o#�M��0��h��N����9�܄�2�jV+��d� �s�]?��<��hzGH��z]^��3[�u\��Mu
rh���:��垟�p&����f�Л�i:�@`��Uz�B�W��W�*n���O��Ja��m�O�IF����P���>J����-��A8L�Z��ˣZ���VU��4�0�D���_�/'0DD�|��GO[b��.�Naf�L��!�{��%X��,>��	h���{��.�?�����,���w�8�� ��n�\��<�QB�J�/�{UX��c�YCGti��*����D��������X����y/��g����ĥ�g���Q]��:nR����nM���K�;+L��p]�,��qS���mt:��Թ�T�����|K���j`�Ĺ�aڿ��^�k�+� =�^^�C�-��������4���EK`�u��������F��������z�XF���k��,��=WA�����tgYS�sk����ے����"~�:��N$��~^x88�m�F=�|0<���Jv�/B�8~�3C��9_�rc�YՑ���W���l�^���\O�b���g(���4' �ө񋓹�����?��d$5���>.��o@ǉ�Ȳ���D���	�9��e�F����������4ۏ/���lC���sGV}�S�;|����ݣ
��)i!F�T��dKڃp\�4�:�H��c?�p֫�z��)��?@��{6��W3��^�jm�>w=���$�L՞S���Jۄj.	"�_Z�{S��U��R�����%2��Ap4w��|�B�s��Q1����ΪG��	m�y��r@草��b}���v��|Z�u��뵦�Y�b�r�M����%Kt������~E�ϝ��q�?t4	�Y�!Iñ8�Ė��[���(�l�<0��-�m����kU�N���<��7om����P�np�q���5��`Gn(�,s���J�ȁ),��o%�
�b鋈��a#r�o(��\��v�E��ņMw����(3��e�QԬ�q>`tft���&Ltln����A��|� ry���I�8�����+��"��X�� TT_�G�d�tW1���D��X=M'����}����}����Z��x=OՀ6|@�XޕT,Y�XX�O@!m7~xS'���5��A���/��*��w3-�'T\��V�_t����P�+�=+~Z���S�K��ٌ�c���e5�G��(y��U�-2�'[#,��zC�8���^��Y��l�wH.p�K&�p=�Wh�����MD�6��Ɩ���{T�Vf��%M�U��Y���a�W9ɩ��(�l����j�BDP܀.��8{�_��tHp��v����v��0�I��қm�h5�M�Y��1���x���oX#�cH_ϛ�Š�b\�jc���8c� �⍉e_�Ǎ�������S�V�n��]Ϻ��sw��h�Q
�+t�U�l����6��m�bզV=����������

�C����8����v ���\g�\�R|��
�F���{��N�����I��Xű�Y5�hy�/V9=���:"9�m�)�:��U�j6�l;_ _z5v� ��^��jn� ~��#��i� Y������QfIp�5�@��$`�䢷�I�JT�(]��?�`�Z���������re�I"a#���)���*�:Z:_��E>Ǣ��w��:w2\X�	���m���0����&c���*۸v�l럻����	_��>��}}߇���e�կ��:��҆[Z�=B���؀u��`kD��Y�0�Dݑ�5N���k`qt�g�e���r�N��M� 1(�W���Z�|�#>0�fV���1�@UG�C�>�1����llG���-ty�u��gٻ��Ա������՗�I����}����n�����v�]���2�p޵8�;�a��tڏ�嘸�Fx7�C"�D�nμ���8iMd���eL���9��Y�k��Y�U�S��(����cƟ�2q:O�h&f6�ӂ~h����!�-�]ؖFF���᳡��ùSj".k��_-�Ɲ-����\�U�G�:E�Ĩ�߸����������<
�gb�Y)�Π?��OMR?"�\�	�2F���1wf[�}����8&@��Y�&9�>U�&��]h��/�ɿ�5�+�-��㩜�B�v�c�7D8O����o��d��5���bѓ��{��\Z7^�ڻI��n��P*�is��8�p_4A.����j-ϼ�N����hb2��~h=^YШ���P�ȺV�W'3��Fbu�o��9��\�N5 ����t��i}|+ =:������w~p�s���PM>(m�Q��@0����c�+#aۿ���S�w߲�w���"������N��v�/��ܗ��=�zB��!���,*X�!0�O��П�΍�X.zMϘ�G����,M~��=�nѲ��|!�nא�:��O4�6�잢%X2Km�!|(x_@mk�
��B;]_O�e$m3���L�y0B;��������j��Ɂ���k��Cb�D�#�P��2�N���l��i�ZZh���~�d#��Ϭ�N�}{�}��������hT�|w����;���a�,UD�m"������ޛ�;�̾�tߪ8�>�b�����htϩa�bp��b'=h-sE���ţ����΃�)�s����V�Hu�Ꮵ�˽3ȥžl}aG\��"��++_M���-ҧ�xdL��H1��=d�Ә��X��|p��F�g7P���X���b�@D���n���&՘G]�iJ{�Ko�6J�O�p���a��#��=ضF7F�;�t�}`��M���m��T�0B����ɻ���rEÓ7��h� �\��G�ȋ�[���ގUN��Nπ$�*�����*�bp%��'N�a�������(�3��k;���-�b���Y|ڃ�{���b"tf�k�=\��ʾ�nLP�
D���
�K���Ţ�'��>,1s�~��+�A^�d��^�heK.��Hk��q����J��"���C��_5�^<�$�W��ޙ��~>#yx�|8�ȹ{��W��_�7��O�2h�K�����I.�x�_�@]tϻ��b �Ɂ�`6�=ˍ^���/�P%�	���l��_���c2�f�z��� u��BEWU
�l2˝�=5��X'hd�3R¼H�;�������A(���n��DZ���]K��Ӭc�ri��3������Q�� ��&�%]�7��
��D��+F'ߺ_�C줣�!��;�a�ՠ�W��AOCL*��Wu�!�hA��w�~	[��]�Wn;,|;�~v��6Bu�s�Dy��n�����u!��re{)Bb�x�e�Љ��|�(��X J��L����B�Vx�`�9\�Z��W�L}��n
�� WW��};�v��������SX�+�G�n���G�U�q�cN�W���k��b��z��O��z�b-��x�6�e�7��:�J����eꛞU���¡�q��<�3�Z��O;�v����Ӣ�s��� N�4��'a�}ɍ�l�`�an��9�l���{-|��;�33'�it#��ר���N��:��7���v�㒌o5�]�{UQ�EK?��ncե��s�=�@_�z�/�A]�ǹi�k▘��+7_'���N4���
��b�^&ŭ {)~?�q!M�A{�����L��?4�F�ۆ>��L�	Z n��i�2�)��qՎ����#z��	���(��ܨwKC�8Y�T+������h9��|��he�G��L1�
?x���}q46r'�=�`��B|�!\)��oh-q`�̝��ж�����"U�1����~�DxY9pP^'����P(�-�I,�����x����G^D�իմ�z&�Z�q ��J;jA�9�B�SU�b�KYI���g���{sH��h���C����/��_N�%��<Λ�Tú;�/��_�=�g�	��P�Jqѣ����a� G���ݧ���� ��>���n�7?�2g�R�1�4�i%U�eo��X��~8��Kn9�
9�3by�Ԕ�J����*��7甥@�tBD�;�����.oF�}v&%���;&�?f���֏�ܘ���}�q�^8�#����"��':�0��V��~��J,5)_>ӎ�&/�?-��ԟR.�dU?`��8a�	a�_զp���N	���{��_.�і�,"i���*
� �������Hw�̔�j��t�1g���]C�ݖ:	�����T�$��Y>7������+da>�,J����`.{�0���Ժ�s���r>y��v��N#�3����Q����ɩ����X��F����O�V׍������a�4�4\+	
�%�ш�����\�7N�%�b�?oH�;bL��5����+5h�T�/^^j�*���>�8?}�����(
��v�.Q(�G���WAi�.���?�5u��ޅʅ�g�4��h�o��1������{�����o��G���~KG*A�ܪ/g�n�+��hL}O󍵜S	{�J<Ck'��R[f|��'������^�\w�l ˽�NN ��]oah^��������=8+�����>9d�|TT�t['�����.�;�t8�vGp;�5�އH����8��������RR����i��67��J����9�@4F
�F��p��;� �tXFv��Xi�(*q�+�s7z��L��|��HA!�Վ��.j�Hh�v�Q`���~ �1��KL�w�G�(1�cGi�KfV��2��L��LhJ�����G�C��e����A$p��Uf��H��5�M�f%3�pQZ����g����z4���eLmQr 1�o��3�c)���R��`���&m�����/��X�{�qA��S�7�>O�9��p�@#����ֈ����I����Y��w~�ځ�U�X��ʹ����� �FبQ����QgX�^��1�{���	�I���EC~)�bÃ�a|�Q�,��'r���<�m�3-Sկߺ�"��8�o�V�j�.�ON�Q���]Q�<��M��G�*�T�g�0�S����Rt	��6����Lk;S�P;2@�3�9��Y�Fu��?ʂ��{V���Vu���[��'(��~���v#W��.��`�mu���ת���l�[i���"��;����+���~H�]�zZ��t���OI�o&V��!�餒ള�S��a�R��I��rL�j\VUqx�����G�0|��r�����P2�2pN���o�����3#P�"�������I�������B�d�3�n�xW�v�I~��CCM�����9*h�ܰ��O�z�"�i�4��(��a����g�S�P3�^����ƔԢm�o����Ы�lbX8������Dc?�C>d�2�V ��;	{�<	AvU}��FW;C����>O���;�7�a��A�T/~��v����^��]9v�r�|/\�����s��nZՎ�K�'�h��9\G��e.s�t��А���K8�`Yz	�2��J0̈�u�p��L�*�M�����rt�S�ǎ�׿m�wT�����M+nK�����U�����a��h|<���<EU�92�������9u��Ă��}����j�ȧ��s��	N�F�?�e�W����i
�y�M��K�����,�KNCw}�����5��X ��Yr�IW,��_��")[����%���l@�V�t.-�?��#���z�OD0��H�!��[d�����g�u�g���H�y���,�!,\̹�0H�U�NO�{RS�:�e�j�	},B�ʩ�7�*?-�s?��]m��|3�s|���.��ˈoO�	y��TR�ޞ�_f��'V"N�Dh��f��?���W�⪱�=����)7������:Q�r�H��\��#aXP��Yd�Æ�P�*㢲�w<?a�E_�_�������wu���P��A��qhhg�۫y7ٷ�K1���[�m=L�B��<�Y�,��#��ܠ~)�/Q@�2�P��G�p<���0}^����L��
"��m��L,Z�϶ɍ�:����kI��W5%Z6�;�V0�&!3w֞��űV6p_�4F��*�������\@�-�]���U�:�g��U]�G�٪}�]�\?�6ɘ0�h@[���KK�U�.tv�e^CY�4а<��<���v:\�E�v�cO�`��UT�󊦒�I'��%|-���dl��.�A�Κ����@��K�Q4�S�UB�@���\��	<
#i!��H�,�&���A��~4�~d�ueU  ���B}k�*xř'�n�wF�H��[}��HUE���lc��W緎)�i�˳������1�}���" V%pQ~X�k�|�ŭ��+r�?r�h��J"���-��bZ���9a���N�\wt�=��?��;3�̸h2�E���P2t͇��O
��Qc�b~��v��v3~�ޞ(��>Z��[δ�94d���L'U���wE�k�����}lE��N-ð�`�Q�M �����	����%���M���V��XO*O1�W���K�R �]�Xn���kQ��p�}�cB�3���o����^��	�-�	7���K�k���_��Ep�̈˯��:L��_Z�¤p=d�ϕ�Gi!v�9q�Ż;6%Hx÷��13:TqX�V���儎.��?�O�X+7��u�E��-}�v]�sjp��֣���8��������]੗斦*<����D���o�'?v����^�Umt�\�rWl���I��%S;�L���6h�Ql��rQ�1�ڣZx�]�FK!Q=M��&R�\E��W�O�f���
p ��.ޜ?�q�1@�ݓY���Y����-��{F��뷑�����K�(%E�cY
�Y0��Q��ޫ�+���\������,2��s�~3c����ibc��G��l5�Y��vڽe]YD���z�k��X����2��×Nt�w#��Q	E8.���1w�M�?�=��bϹ��M��7t��8|+(vn�:����O�@�B���
&q�!�3�;�#��ƴ"�jx�&�r�>u��ǁ.�Һ�a�Ԟ��^@��FU)��V�n�����'��L����=)�/$=+��N��H!q�8��Q)r8U�+��fb�uamU}�<W�wS�>�8�]"u�뼢X�1
8�JJ�ߠ#�
i�&�V�ۮ�ȍ�zb��~�f/�O8娴>2����1	�9�)���S�������t\:{�h髸��d��6����0����0�ы��i}0Ҁ�ӈ��'m����װ��;,nԅEj �@xV��J��I���';�L�a�Ef�<��^��wć�؈�(X� s�;d�u��CT���:�/nz	�c�&�ٰ��[�Dv����X�D"���bzp3z���& -xVӫ����D����Q�e�}M�����'�i�eI�y��޶a��g�]��botZ��G�n�&ںdY=ܔi������c �0�h� ����w#/�I6�,�Cƿ�Պ�2����H���l�\jý㇞��԰��=�͖!��K�طތ���~������x����vԀӼFX�R8?k�����ˇ0[	ϔ"tӾx�)�B��wg�6a�ލ�����۱w��8z��	��;i <h��?u>^�Іic�Y0��� �N��-��5��qs�~�z���X��zY?��)�SS��D����A�y�MH+�����Hڗ����C�}N�����81:��N��у�!t���>�P~'�dE+M!�2śd��v}aQE�	#"�	��X���2�C���<ٲ��e���S3�&������V5�l�+K���aaF[��oq�ADt���7{��c��q׵j�cڠyyFh������	|�}o���rD�1���r�4b�=S��B��x�{�f�j�	�	�
�
���ss���â!<�惺�w#2~1�D�#�Z��#m���U�E�:�p�C2�L8��*]斑 ��v��9͞�'J�<���w�@4�:���&U����ބ]<��K�k>������W��*����N�Qs1 uw�*�TX��pO����,�.��
��&��6�91XL��CG�\�$<��s#�	�=�1�eYgQ�u<�w�ks�A�k��cl��/��O9Τ@��k���t�6
�s��� �(ͳ<�-�r��+3?�������x饒��tT��Ղ@f�G��TƔ;㩆���9_YE�-��a�� ��א.��ˏ�m[`�'�]���x�A��(H��z@m��J+
�(�9��e�0��B{Y����i��n�����szFj*�v���|jb���LF�K	��Ś����o���-�L�Z�>�ن�li;)D��jg|�L�,$���n���!���i
��d]h��+��~X^�2�������O�0m{���]4H�d�N�;���xDe\�7�Sڕ���eV�b~��	�������@ĦN .,gUh���xu�[_��\�jYr|	VWy�w}�_ڑk=���J�<�w8����oT�5JkV�"Z{�a�5k��;�)UTQ{S�WP[l���-�g��b������\�/�u�y�s���y��s�E��n�s@t��L��y'�:[('�3ŀ 4Bq11C�����ů���AX.��
ą���v��;fn����*���.3v?�eq���L�S]�Z4DEcBN�^��N�xkt�Z�����Is���͂_/�l�n�=�8��9�r���߉�p�>j� صS]K���1�l^MY�N�tW����0�r<
�\$�^ $s9.��O���͵����MxՕǧ�=�\ɾ��>95vB3�o���������l~�f６���M�J�x���ii�ƀa{wr}�[hċ7��}�,�˙<���NQ'�^p��X�Kk�GYƲ���/ֻ�=F8tF�}��_e�\���(=�o���'���ĕ�<NV���[���P˯� ��&��AD�F����j����(5�v�Ζ鬜��@7
��~�1:(8n���˸��2�y��̎�_+9���2L7Gq9ܔB�݋��J��~4]M �����w�E���A�l5M�|��DҶ=Q�(���ޣR뾝V�N�Y��/g�Ǔ5�QuL�ԯ���)W���?�bU�4b��fP�'�a$�.����v9-�p抢j�^l4T�:�a
��d#ڱj�z�D'�E5��3�����dBJJ�12���*���T!B��T��on�k���"�j�׎ߜ��-�ch@;uy��������hq�chP�g�M�X���a�%o]'U�"	l�S�m�r���^��<΃Fѹ��~q�+}A��\�P���!t�k��]�H��h)`�I58��x���xaW�zz�α����r��f���ϸ�٩�LV�1b�j���^t� �8���~c����h8��8:>�W����үsDG�݅�U5� �J���/1���c�k^l��) �#!	���=C\���+wH��ɳ�8��9���0�/����E!)I�x����Awː��<��>��߆��lE��a���B��D�FX=��3���TĽ�����h�5�%0�̝{|��_F��(���S�9<$zhnnD乨,:���C�1�����Df�Vp[P(���~�����z���֚�\fr��ҟ!@~q�-Y��1�UfR�Y5f C�����A�����E9�_���[K`4�Y�p`���B�);s،`��z^�j:�{�L��lE�7Ʊ �xSg�l{���OQY[��x�~x�i���ћ^
0��·r�E[��K±,���}Hn3b��f����PN��`���B/O�37u�/�V�[M�f�v@���L?�Ѿe7ԄFf�̩��Ϋ	9��N�2L�d&�JJ����� @�V�z��|S$b9��>
�:�
�#_����J�޲����m�'/%r���Ɵ��
�sݚ��sW�������߮�S}КM�0���;����s��D������#���=�k�-��!s��@��p��-x��N=��$���I1Uܰ���^�E�������Q	���A�	Ԝ�ő�t�H䚦	�Ea(:���\�� !eip`$"7�)Us,C0X���H��J�ࡓ	�{E`�N�~��}�W9����JO�UF]�:;��8Z^�����'�tᗪK�`�3����1Bj��<NI��f��MW�<ֽ]��W�9��)��m�_�����Օ�^��-N��/�t�����A��2Eě܎ʲbN��>yY���1M�PvM�j5ғڼ9���6�a	
u��75y ��	�r<�bޅ��_�ޒ�A�_�u�Iz���ZL��(��CԱ�����{�;J޷ME#����P�A���\5rr���d�s+��T���.���뛽��".S��:�߿���L��"�,=`.?3��1i�Ao#�2���^9����f_�ߡ��\� `���'cͷ��a`��s�׮P����y�V[x�cp*�� �����!��W҃�G�'����D�I��hEK��M���*��&,%�n?���YS��}M܈�3����jʬJ�����t�mh�e��H;��w�c� ��8�'j9_+=|���+���+��2����X�j\�b�e���G����߭�v&C����B��YD�R��^����S�l"'?O���>�Y�(�Y�ـ��[�M�Ժ��3`��q���7�ê������T�����e�&����%�~i�j�`??�I��� C�(e��m�Hy�EX���h��C�1v�M����؈�����c�'�A5�j�7{f��#�f8q���D��ڠ�-֣��6p��BBf;jC����R=]]��O�Ξذ <o!�Qt���Ly3���gj��j�R�M��h����ϥފۋ�/�&�{�Tg-<����g,�)��.�c���4E�6x�U�d��N��T��g�T4I���n"^2�����I)�}�1؊��#�餔$~�.����$W��N|��&���U*]o������c�����XWpj�]�
���$?�-Gg{3�5�{���C���f����)���=�����-G&XP\�Ҕ%���9�l�{������j���>~�u�=w�C|ˉ�����))��g,oDa����ת}�m��S�Z��X����"ES|L)�9�ݠ��μ���+��E3�����[��F���SE�6
���ƛ�ޭ��BF}'B��I���e���<q��ߍ��?��3'��w�:��D�Cu�T��J�Ʉ��(M���m0T8�-$�1Y���_$�|w���2���S��67�(��UJ��<o�g�i��
�t<N�^
�k��Z�.{��eI�V��O�*�)�Q�_x+�u�G\L6���+
D�I%�p�D�	-�Q�~��?y�{�|��(��S����}�"K����ss�r�}2��2����\�ܒ@�- 4����w_��{77��>�oh
�������~REE~���}��|�J�p�1q�@�ͻ��7w�B������:��V�N�Ka`O����cnX�堤���� j����&����o���Y�~O��)�=v��1[�*/i4!M�b�^���>�la���	76��	L�.O����O�m�@����x&���L}���y��}ʰ��T? ��:�>����k�z��a���VR�=H�`#Q�$�flw�[gA�t��L[�u}u�|��{�V�������-L�;"�<��uc0��+��VL�b�F��\{C�\���Ht�U,�������{���ϑ�	��M�a�/םUt�����fM��N��$2sO^��V""y��t]��2fxC]����� ��D.��k���85 ������;�^��n��c���j�1j-{s�l��N)�����g����A�ų��k�Y&���6�*��d*��u��:��tA|�"Y� {�%BN��l����z�44
��Q���J���OtJ5���8��cy�VH&X�l�V�>�qt�
o�z
J�9�8[���ӅH��H��n�I�n!Q��ʘ>A
p�ʍ芌H��d��b�#<�:.�Ye
Bѥ���e��]���L�\�Y�Ch��SMQ����
"�ڛ�$+���\_ߖ�TF�i��k��_�AL�g)d%b�b'��t}�g�9D8dMmβ����7�/�d����8�R8�q���l[w��a!�������4�>Q�mcnX�.;�htm�gY�����Rw�}�4)a�<��{�]�Ox$��4\$d������9SIhI��ٖI�D���~!��0�NYn���.���z�+ڪ#`��O�}ȱ�`�'��CB'^�joi($��f��{j�w������U��L� S��w�Q~_Y̿G��(�#kvS�l�R�XG�8�!F�gQ����k�%�J�R��xL�(i�4���t�]{�-q���.!)m�����Nh�+�fkoZ�#�>5��b�N �W�_f��n_��8�P�x���&9g;z��hp�B�.Q�ͽ�İu
�����o��X�� ��<lL���m/1��bZ�Z��-��M�?���8�Q�݇ ����XW�<�{�;[�GH��qVq�D�����߼Z{H�W*-���IzERO����?x=��AS��^dA1���+�
;�m��Qa�E��$h[>����ż9���,q����uhO*�����̔�75t�ɑ��0�-�⡾׷���'i��o�OS�)i�ee?��wvY�����c��*�q}���*�rh�T���l۸�f4���$��<���A��h˚%!�#��U$7�Ͽ�ۢO�����	`Do&����U饅�ǅ�l2긘%:�k���"���;��D������(�
q��z(R�������!l2�3�{�P�
��*��*̩�R�J�����=���P��r�� �=�A��^��dl̤�N	 K���6F6	
Iw��i쟖�-���t�uI�,��/����	�8~'�ι[�+��\�F������o�i<��b��C��J���xBډ���?�xYE�쐝��z2P�+�~r_fE	�;���s�q1NU�.wp�2�����s��*�/���G�����7{�8Ga��ʹ����!?���k��KH����@����&_��Ɔ<N�?���#S,�O��3�I,yh����=�U���F���c�2�����b��3���%�4;;;W�T&V�	��_Q|4傕�1��t���S֞0u�>�-���ݤ'�(�o��x^AÖ������[~�|�����k7��B2a&�i0��?�]�3 j?}&�X�>ܼA\�����ĞM��t����T_���X����`$����O���]����/�� z�M��}e��L pV�L��3�
��U�؅��\�_�\��-�;����bϸ@���K����ۼ'��Լ�.����1$S��$j��̏R��_w�5_(EȝH&���1ay�$�a�&k�8hVA[eq����1C�z2!c�3��(���5+K�Z������&��]�J7�Y� ��+&Sc�1��˻y�������Qh?�{�z�g��.9l,xn��
�Ͱ�k����К��8k0�i ��ᶴj������>�h��v˄��"Y[5��_zV�ܗ�����.��MMf�u>���:��Bw�z�KqP��U�Q?��'�\?�9Q�Cȴ1��@�c0�c}5k��4�6��*�s]�h]���0�ZQYj����
����)�w�Ge75���1�)a���979ƭ`��V:���Z��65�M��&��� 2&H�{��؉�o6��{*�$�
E���,P��	���%N'*�9�U�b�߆�f!+���\<�h��߸JK_nޜTmਊ��Z�V�8u�Wzk��gϋ��/�P����ͣ�ԏ����
 �G]e��/$P���8�!q|�����Kg�}�|R�kݫ�U�I�j��=?=��_yR_=�	(��<5�O�߇L�U5�I�л^լ���=y�ظ� �-����Bh�qv�gA(�H!��4�?�	��~�Ul��o��~���9W����ÒA��IPd�P��5c�ca����=�:C�a���:a�ϨtCv��%��l��>����t�Ff�e�d�]�ڙ2�@/�<�G�^K=ґ̀Y*����N��q�¿..��N�ݛ��?-QM�2u����M�o���Ñ�'%>�1�P�ao�(�����.�P�����jW]M)k����n�^8�3���۸E��5�w�v;���t�"-��ۤ߫����a	oyvÚ�pB2�]s��2�f��9���C��� �[,��A��%�A^�Fox���?p�`R0�3~�y���a6���E�d�m��`s����ʾ�㥅�Gܧ����J�'�Ë�#�ݸ\������EQ�� ��N���w��8���ٞ1/{�D��<�_�X6���g!��!y��Y�qf��5ߞ4%�x	�1�
�KZ�2�;nr�;�}c�r~����dT�	I����>8�Tk1��@�������o���E�4��Օ��+�ᢗ��"�����T�]ŗ�4���:x0}qǩR�^|s�!�K��^�T2�~`]
�%����7�l�"E�Գ�X��>?��Q���`>�;�?q9����qW��ڗ�ȼ(�MR:������f��R���E�x���9tl�Ϳ�K���l��~FR�4�CW�3�NRwO}��#�ܾ-v��
�e^|���=4��j����J&ݕ�3�H Z�T��$et[�	X\�e�a0�9�	Lyn����.v��yO���%�	���<��+���Et#��9��R
r6|���4���˵D�6uS�1��F�l�ֽ���"��Ԙ�~��<δ��Ο���ԭ������L�v�l\U�2�Go���]18��?`;�b{��P{{�'�s9�#��d�8�])��F]�ߏ�G�K��n��~@Q������S��M�'k?:����@pT7f2:h08�����rۖ1�<L0	V��S��	!+q���2�>9y�n�N�oa�|���j�zGӑ�[z�aI��!\SDWk���S�
4eܰ\�L���{���;����#�AX���Z%��>�g��=���܉G�+�oH����WW�$�E}��y�,�I�\jg�"uI�X�4Y�1��+�ؙ����~!�'�ѦZ��>X��;�܋�{�ɻdl[�2.�_���qV"�䲌M��6T�"���|e� ��U5����K�?&�蠵�mw�2��7n+�
�3�8.(e���X)�s�B��6�OK�%z%�4g�S�<ꁮ�;Qʏ6KX*�����]=��v.�B;S-���e0S�p`+�S�@ǒ�t�9��lVx��S�T�L�_�wǴ�p����[__}B�KZ�7�^s��a���j/�:�K��C�lR��j
c�#����O�td�sk�׶�_���m�!�)*4�<������3����`�~[=+{��ڏ���H��V��n+,n�o�>�P�p��z[ɕ���h)tx��{_�4�r���*�w$VZQ��w�H��k�*�h<�:ۢ��Be�Ka�g��Wɘ��$�O��|���l�*!�a��Z��ʱ��c�k��(��a��OS��[�����Ic(>�>�,��H�/�}.�EVv�U_�k�h
���A��4'h&�W�������c"�ap���G�$�/������h�R���|�V���a~��
��&���T6��+������,� �Ul$$kj@�P?g%)=q�i m���){��Y����t�t����*iMd���Z��J���Q&]��{A�fO�AH��(
:e]��jU�⡗�����?X����4�~������в�Z[]��2R��3���}v�6�@cQ �DK�����1�{���_z�8�b e��t��n�[���&�2��=>�� ��ѵT6稔�Q��r?|8��kL��n��Kt46"�
��_�=����2������WA��Wh��a��v4L�Ƀ|l�?כ6��[�.�>y�ݥ�NRFVeV���g�f�U�)lh��R�#�#S��m��('��#��A�r-I��d�g`Q�Q����{؂>���h�V��d^r����}����;\��h0_\��2�aX{��.@��y�犍����;|?��)���]#�9CK���������|3�tυ2-C�e�kw�]��3����� R��#̥�u�Z�[�v��i����q؝ �����̏��	.(N����>�}��T�����Ӏ�>1�h,MܨK�'�Š����	/��o��[[O�jQ�Dէ1HҊ�Š���O ���?��0R��su�e�E�O-����	d .�oW�1,�e��j)�6�]sc_�1V}kl���Y�m�ʭ�hcO�Y�eȎ���a����L�ppT�3NǦ���֫%F?:a����ԏ��%.�{��(C�I3��&W�|�V=:�'ϗ�5��[w���i�����8HBr�����@'Ht�H�hX7�x�q�Oݢ����]I�x3ho���B���S�[Z��o��{pƉ]?YN�|i��|\�8:
1�y���`�l�'��I��Z����K�&���\C-�-{�T��Wյ��}�u�u�+9����1A��thj����n�z�x��6'�{%Yo�5@E�gZ?j�M�����e�O��Q�4�_ʋD������^0ed��ZP���n�9���F���(B���\`s;Z�%ͅ�2@�͏p�1RM/�Kʭ�_~|Io~�����#_O�^���3,z�'�܁4I	�����n�pp��6&z�}��a(��Į+-�4Z~�\�9�ڬ���j�W ^�'����6x�����UT��}�)�J9���'��Z&!�R�hʌ�>
��C�-Fc\dR�r*�P>P�Ā��k�*�hG�\t�j���fT��;j濲��3����S0O@��l׬h�4ɘ���� ������]�� �f��si�K{��g��5�K�53e�}ó+<K ��v��V�r������UXkxMwOL_P�*����lB�[�4�tJ��;^@b��1>N�-�Ԡڸ�}UXZ���ͷ�p�>)��sz�=�ŷO�^\��t��ߞ�}������mê�cv��c��H@}�;�L+(Cx�o�ω�G���Fx�/�Hߏ�X��!�L��`,��S{`$x�!l  �1�4���a���O���k{�"C���+麆2:#�b�4��u��[�"R��^�&�w4�7g=�ú�V�����L�\�e&9�6S���K���C�qimh5�e��@��`������lS
�~����#��X!BA�+Ӹ�J� �o�\���~�߿v�h�}D(�r�4	}1�,8	��m�,y�sj��6����|��!���噙��2�_t֥��AA�`�|�d�;7��yH!�-+3v�'�v~�G��68l���%S*�_&�T�
����N&�ا#��%�{�e�u=m�DHT_��y�5T���/��W5��$������\�e�ͶF�^'�R����ݨˊ�M��)W��'q(�p�b�Ϛj��(�:�Ǝ���֪�sF��9���/���=g_C��uL�	k��e���]z�#�I�����4��B)����Y�n��G�`2)h	�f`��!e��2^1;R"j@8[9{#[�t�3�%��j񐝧� ��  ݚ��Ӈt����az��z�l��2W���˞�"���b����>[��]�@���lb���׌�	ppX#..yᢳ;���=�%��;%ξ�+�ʂ�k�ˏ�"���^�pp�v0�ˏ���9�]L
1G��H�hүw�.�4me�f�;JQ��N�����6�ơ�]&�T��}A8����5�k���*��M��ee�W�c�:�'��+yY����^���i��~�;}y��MJ7s�޺b�<���#E�6C�H�UZ���|q���Q���㦅��&��d5��>�"w�R�S����*�hKt��(�����N�� ,s��4�;I1��^q{KcC\�96���%�}�4��I���|e;dW�>6���i/�<�U�89+_����n��=�z`~���mni���ș�?��;rW�c2<�����pRMAL��(�u�6ǿ���tO��Zq7<�� �f͒6ђBh��,���g��
���S+"�tq:��Y}�*�'�ͦ�?���̀��JB����gl+�߯�"�:���Ƶ�oP/���m��A%:��W��i=�ָ���FW0������,X���VQ)Q�ES��L����lJ�z���+�~��v��������d�eТ��D�q����~^������m���Ӏg�Q6
��ru^D�s �R_Xכ���.����}�et~?�9��Z��b�Z5�TR����]�&�=7V�I��[t�$���n5���G*s����E��J�ݲV������[��xӨ�}����t|A�9TOq�G2θ�>�V��E1���_���������gG��z�;�ݧ��ǜ"?a�.�7-�õ���R���~O9J��4ڤ��H�&WRW�[2b�"��0ф��mn������>k+�ML�^���]�	O(6�����Y��� �'<����;Qj��ߢ�]c�m�{;���$:����m��]	3���z^1����G�8���<�p8��p8�-�8�(�4ez�V��"��^m��$�+�m����]�y��Ś�9�L�9z���)1��6`�4���.�K�/�$���<��3���672�sV�!�Э��%�%���o��:���o"����3fך;
�����Y`Ҭ��g���� [�s������u�x"�y��N@��6]Tv�p��&vuQ=�~Ta�5�jx�LC�'�;�����fa�����N���u	0E��ˑJG'ž�O�]���!p��o<j�$%�d;�J�{�b���TpHg�t�a96|��0-PG6c1� O��{�_��a���\I��F��Z����Ʊ3?:�����b���O�Xy�U����K�4�e����^�bFH�	{�t��5{�����QpN����l�Պњ\'�A?}��#Y��5'6gl�b�=+��c
r6-���;9�P66gj�O��3�:pg,)���8������B�4�8�΃��r"A^ ^S}v�C�#,s����tM��'���u���*7����H�f�z4�,�-�����z]��ggK��TEK,�ˊ_*!�X�Z1Rqy6�s�Y�)}*R����v��|2vTD��ظ�5oH�� T���Z�+��;60��n<(	��C�&�^ش�|���A?��ao���V��?�Jsw�2�$���x��3�������`���f���6бLj�b��߿u��7)����YZZ��H[SW"����F�Z�??���5��6+Ȍ�!��`3e=`��L������]�[���K��w��pI7��������Kx�EÏz8vF�,��AZT����d��v(��1��՘Jۖ�#�����m٘����Q����j�g߁���j\�v<t07.r�(?�=��R�g�R��ͮ�Q]ӿ7]ù�U� D�m�wB��ѻl�t��(%S:jg
r
���"W3�ѝ�6���)3Z�@��_��|k?�~vh�gM�TE���M&���a;�H;�|�V�����=v�s�7[�UN��d�4��E��H��ܷ�^	x_�722|H�S$4<v5}v!g��)���f>ݯn��EN,�¸ ���7g5Ɵ2LEe�'gLxݴDJ���VO'�w��XR��{;��y@s{n��Avݠ7��p�Eu�^�t�Q��=0��9��aHJmA��wŷ�k;5��`i�y��b.bS݅Ӥ��88�X�p�}�uT+�k���Y���=f�42u��a"������1a�9��C�7}���zu#��ĕ����7x�,/�[�Z���)���#�"\L�pGH6R/0��p��'.���E9ǐM���lSٰemѬ=^��2S"�&2�8K�(�Z���{˻جZ��)Ԋ>ld�^t�Ӓ�0�s���f�F�؂���^-���^�J��2�����l�s�$�'��E��"��4;�Ǿ��>(��Uz��~!�_맋��X)����l���Ϸ{m2�����S�ً���R���j���'��Jx��r�d9��A+�v_iY���Q����a11�F�(�Hqe�7&�ox'g�&�������J�9f�e6���|�H������$J5���dD��o�qt,�	�q�]v��)�Y�+<�C��tU�%~�[��>���a��	�>�_�O�I�/�~Q����gPqCF�."��G��.���K�G������[����N�KR߯O�_�!T��
��R��\}r���Z�<�z�%��
eهZl*>��ܲ*QJ^��}L�}������Pptє��5�56h8���M�v-K�p�^�4L+_%(�|)�>i��5u��e�%?v\\	��7�P�������*�]�H`�PO!*�k;�3#(N���y�o������e��^ۋV�kf'�!e��ׅR�z�β�o���8[�"u�-Y6Xֻ@U�V�d-( �(	�&^7��Q�iU��=�^��q0�6`���&%O���Eף��`�Ӌ0�1����M���0�O���p�б�����{l��S#,�:�*��=J)por"�ؑF	��$.��2�H�A���E�<�@�h�0�t�������+���������?_�Y�n���~��Z�[T�b�?��C�f����^�R�Ʌ��V��賛ۅ�j�a�8��)룫7�Ϳ�={5���*��v"��#�"{a�ﶣ�FN��(˓�#/5��[��Mܞ��L���$0B{^^c�`�	���$��,#Q::�M]��I��&��8hoѽ|�^%�֧��_n|�@�(�Mlb/��|����n�J�G���%5bՐ���
��Z�T`�Y����Ͽ/�0��X{��״A��F���a��.���s�!ݍ{8���d���ǧ>0�G���J2�z*]�4>w\�]ӂט�[yX�r�G~�x�jgN�3\ȍq�>`,01;�凫⿙d�.j�;�>y����L�^Ϸ����ۊRO�MxVm�$�Ȯ'��{��$}�/.$��94��1���#�LP!������y_��C�2wa 4���Ic RrX�t� ����eR�Nwˤ�ߵ��"�/VzacĞ��9��Ez:|gw���Ge`TCg �&#���<�,��� xv���̌�2l9t�ĺ"��Gl{z�E�'�3���c ���T��ck�(�a�Իs��1ЦT#eYYɭ������fG�wv?IyH����/���lm&v�ռ�'�����R�*���7S���ϸPw0[����G��<o��A������>"A�b�Q��4"�)�"@a`�z0ۏ?�L�"��2�ג�-A9�|6W���
�hfK8fU��"[5����\ֽ��f���� �A�_��S�M�i�h/'�c9���B� �L�:�u=���ʞ�N���x,�a�=2M��*X�ۍ*y@2
/<�S�إ<�ע"��=E����^0���\��FX�GHP6ڟ���(��@��Ԙ��x��A�w�~�QoL����qm����e�i�%�MO�TR8?�D��$�����O����I�׶�	�b?x�(;�G�+��M�;� ������-�|A��	_���D�Y�Ri�aW7��U[;4������u}1p�i��CY���r~��mw��$���1Y���;eC���M�������G�|S"���١-Ri>t��y���F&<�8���j2��	��]:��(��iKK�@&�+�Ԙ��2;ͦ��1�nHP�.���GRm�j�}`��:;�aX�ᧉ�i�������7�Y|����d�\���/��9��y�ӦE�e��Z���r�n�*Q%���P��^�RQE��ڼV�_�_�%8���6�"BK[��p��&�� +�KբX&Yk���38�׃��&��Z]2�c�5�	q*�z��oJ�����BP-H9�>�+?ݲ^G>��螖���Bf�{����;mv���|��Q���IQ�`Lܐ|N��
��7<������Q^�`����_H�<�ir�$����&�u�󺩍"/ftV�w�B��R�*R�;�%����L�� ��v��6��6������.q�۪f��(=-;/�m�L�x��J�Ֆ��y����H���ǃս+�Ѩ3J��%�z���c�A't��ꖸ�@���g�}���n���?n�:�����4P�'��$�O�%AX�oo7(?��'!��%��p��8��S��ǎc���j�D>���dgZ 	z��j�5�'*�CX�Q�k�r�=On����` ��J\B�2G֟[�������-�&�R�;�bi�p�O%W�}����nc����ce�X�.��LQ̎���3�ժ�[x�i������^@L��G�.h���<�(�8b��K#\W#�h��'ի"Fʱ��R�S�~Tg���̉442G.��^t�\u-Q�J����^�8]eԗ���K<l�IPg�~u߯ĭ���{�G����^�f�(��	���{#�6�9t�2�=Sh��n�M4i����x^p�eQT��������+���P�7y�j���$���Ek����c�G�H-b�ܿo3�a�P��L+wX��9��_yh��t
8��D�8~Hc��!O��� �v��'�]'�r������vY7�Vr���ܕ)���Y�;�$�W�dߝzh�O	i�!\<��]�
�+��(��ms�!9A'�r��C��=?q�X��4$_#�!��q`Fl�]E9 u]_P	g�X��_S��J�;#���Ң�܎��7ZV��#��{��F%X�4QSX7�y��@q����\ʶ>��Ւ�r�XW���=�G�*�Hjj�zg�vyZ����a�
���4���M�]CO���M�%+뻎�)q�G9OY5�!�Jy�}~�!���� y�m��� �6Ce�$�9�sc��(�J�i)�w++4�+�j�m�Q~{��U7�zTk��Y��P�D ���]�k�1�@˷4KLoϲ3�ĥ29��K����d՞�NI�m��:��S���iF:��i	���j4���*_�֯�� �O�;N�jD׾�"�$�� ����o��$YN���-��'������7������������1:.�.�3)�:ZK�Q
6����U�_��V@��(+Xe���!��z�O�b~��p�6N���M8�<d����O���7����0,Q���y\�R A\�6�"����SW#�j�P��N�o���1] ؍{�m��\?��=KpGܮXC��ā{��d{Ý�^��J:����e�uL��烩��j<.����L������e=J��<��X�A\�N#��osʊ�(�7$�����a�w�9q]�0'���ݸ��E�a�bt��t��c����]�ƕ��(ϵy|�c	8���8�*==+M}-�,��Ȥ��B�Un��v�����)�PH8�@of#7Jn�I�T� ��r�pWiS�����J�j2�T4�V�()x�ċ%�7_L���	�Ut~�����"������s'��H�}����Z�։��˦����?���
ج��B�R���Fws,�eov�k����ר��:zv�^Z b:ɚ�kz���_Y���{r�d�<���B��l�8���DE7U�]�]��,Ȧ��)�WƆ�dWX�u�Oڃ��?��g����N� $ ~��������{�hP��[*���sq�}߮��N��x�;���4�K� B�Vt���d�#��/���*�rJC:~lQ?��{z>��*���9#��
�\���?!D�bL�y��6`v$lSOY$�J �(Z�@(�X�Ĩ���/����[,�q��{+
��DȔJqߧ{�
��K�?��0O&*u����&򧫌H`_JNʨ�8CL<^I�?�"cP��E��R,j�k<ȉlX�R�������O�l-�j�?VM^KڮW����иI���-���S
� $Mϕp����b�cJ'�����#�����7�E��k�U~��~�ŰU�q���X�N�d�7pkH㎌�������4�Ҟ��yŐ��\�{���x�.jc%)>�~9BwvEtO����jm����E�%~\��)J����鳚����w2� ����ȑ��ܬ|��G~����C��Ĝd� ��(ߖC,b����y�J)���~����z5J�GҴr��'��Ey��.��$����p����m?K�w��J�� �p�@��#���O4����V�J��i�K�X��qJĺh[�t�	������yXф-��n\m��y�?����t#F��B\bG��^�%ڇd�@� id)S��H7�
`��Ƥ�����ys�M��eq�6E�ph�k$�6��J2�����u)#X�F_��9�����̖혥�c���o�<�9�?T6���4[7\��AO�d�OD��vk�5��ԫQ-�����׺�<c���$��[N��9��Z���&I��������h�y��f���r7�F��z`7��.t�j�4N��O�l�����(L�n�;^8��z(k�y��2=�D<�"�����(������� r����;2X��_���˻Pxi����o(��F*T�g�J+]Ȁ��l��g�t՘-I��*b����@|u�|7R�]�[$hH��:����!4[�4������5Q��o���@p�j��R���h��v|�v0���C8����{�IVb�l�͕���|}�ٍͮ����f���i���XO�Q�#,x��D�,I_��㣵�Y./�[JH��3X�n0�VF.f��7$6�nV8h-��vŻ�{����KBAB�D��E�Q$:!z/ѣ�6%D�;�(�{��d���3�0�1<#'�s��~����g�g���GȞ����O�{����.�'����*�V�7
'��np���w���t�}/��:���� 	�ݓ�� Ң�'��ٻ>�8��f)p��x��Fdk��)�lTh��,qZ�"Y��_)y?���)�9d���-X˄���Uj+sYg�����z�F��f�@@��n��j��6��:�2+���Cj����(kf�`�:=�c��z���b
܃�K#'w�|�a
1<��jԙ䩚�_f��El��*�\0R�l��>�L��E�ْ��o+�&�mڸ-�v$	�ȣ��}�pV��ĝ���r�v��=��w�w�1��­|MՍܒ��6*�L���*�,A��#M�[�V<�) �����=�hpy�?�8�` q��|8�̄9�xn�{Q��MYsC��y��ɞ,�-Rͥ�>6�U9�kq�;�&�����O�V�,O�:������$[-~�@r��ұ���|�4�������/�1��g�����7��ꭃ�ށ&��� �-�h��9K::�Y'+�{�Y�.#��Τ�<{GD���W�5���e���7�%��E��p�UZ�X��+W�*�q3ۭ�٨�[5w*޶��!�a��|�{1��x�.�f�Z0�G�cRBc�]�CEr��=���|������/��qG�r/{o֋���=�8�M�g�v#UWs+j�&P�N��Y8���MɚG�֞c}�Q:ߎ%n���eP�ec����}�$f�g�P��b�r@IT����x|�2�'.d�S\��f��^�ɝ���AUՂL�4��7(�n�{䤾u��4���	�}S(]�!��E�缟��F��*8:e�x �AL�b,Xx8!m�y�P�=�lW����f�7}+(p�↭�\���=����v����l*�p�As��Y�*�22-�Yώ?4Gel�ɵ�h� _m�ß����r�=���}�ך~aGһ���`s2+%�a�#>� /&!��m����v触/��t�`�T%��w���s?��F��,�t��	>�-�,�<��GE3 3'��c\�-q�٣��p�/�Qv "W��C^4�h$�d�Ě��0��*-����O�A��>���K�����K��"[!��:����E�O�p�<�<��5��p�"q�mK����܃����3��Sς�Tܒ1�Jq9���N����S��-�{FL��Ǟ����e���ב�8�c�h��K2�|�@��^����b�����L���a����-�>����Nh�B�<^P ��f�B��l��gü�C����D�?s	OO�u�Pc�6ƺ�H%xZɑc�2F2�{',p��`2H"��jټ�F�[��
�E?���;�|�Ň���G�����w�k�g�B��6Br3n�6�y�^ϙ��O���ԗ�̙;c�F���Rc�����\ڨˁ�j?�7FA�4�?�`&iR����Z})��]�����2�WOu� DU �9i��k�WV�1��4��I�0-;q^Ϙ����{ax���6�kJ`).Ԁ��l�p��*��(����#�����ڍ2g.��gftIhLɈi�aT�w��3ˉ�GQN�ɕ@��o������S*0JF�۲j��K�O�W�L�T���K�����>�!ۍKT_'��f�M�]��m���f�\�����k!���غT��o�&�$Ol��u��S(%I>��e�1�k{��#�����,>�j���mL���
�-H�`��RLp�։E���ʱ�9%걯&�V
5D��=��A��-��Y鶒u�>p�mņ�|��M���;ɛ�SW�7��iN�ֱ�v��
T�����ȟE\�/f��!D�]t�)E��!&����YL�����Rj�do��k҈ǹJXS�Z=n"v��
y�Z�h�`���4��J��e7�G�t�G�#�i��S�����^��R�m(U��^�q��J^��.�8�=+ՄI��Œq�� �k幊v.��f��\)���s�Dӥ�U�q�ڤo�g���>�N�{l�oy� Z:�#w]�*M;�i�FS�0"�9�����-s�F�ίr�m9��w}b/�v
T�W��N7ip��`�:�A��]���JHZr���P�а���*X2knTi>�ֺxv
��s~R��d�c��tN�o��UJ
�e�B5�
:��%�s�V��4�B�m������#AX�E�Q!ʾ<g��`[���Po@*�*�����F��8O$-:�ō�+���(&��dP�����m3��U��z���7�ܑ}�A唙~��;�`���sf6����o*n�R��)�����[^��hf��M�蔯��o����%�Q%��X�2B+��,�ct{�O��xèKC5'E$q�vK���>�)�r����Dp������W�ҺЗ��>��wZ��5]��c�M��yɪ�#I�8S߆���B�s9	.�����[K��E�R��B��S;�}<4瘄w�:�X3V)0�xt���~�]���I�U}�Vp�q�-�eE��j&�#����k�$w��qK�X�:������{6��nt��/�1�z�E�+�u����P���j8���ˁ}Z��uK��ڴ�hEo�ߔ��fQϡ��K�+p�"��,y�nnm�y����B{��J7�i�)�@i<�*w�$��!2c�tÛ�Z�̉�t��>SG��U�H��wVڰeѺX�a�N±L�R@`=,Y�ýq�_p��V�*1��yJ���$�L�@P,�E�l��Wik�d##�!ϳ�%_��w�4����͕s\٧5u<ʗ_�C����u��j�m����͎��P��߂��g�U����f���)�q��b�א�ϕ�}���f���L�3m&S�o��*W��N.�z��S0�R�f��Q6��Z��$�O�re���e�ݡ�~�5�JqPo�ˑ�.�X��oԵRE��xp��@��3���\�+K�]�E7�`D���0eܲW�͎x�kA_�@����l�ͅ�۶-'8����(���6� �d�[^�c�>x�i���m��=�OwITq�*���ζ�㿌��H<\��Sl�%�3}�r��p�-��3����FwW�R?S"����RA�UC^����ۇy�=I��o��`�E�dh�?�n�[�iF�hY\YZqIK����[��s������5\�wז�q�0�͌uP[
�:���QB��E���!��9��.w(�
b2�'��/`�$�-��4yW��?�@���B�*���w?�?w����)��8h�M�V�Ҧ����c����w|�$�QǞmR��/e[|�v�<?Ϧd���<�Sߣ=�A���wKY K@D��LqN�v��]܃N9�T��R����F�?��_A^�͋O)9)�'�勛�xxAw!��x�2����4��+UJ��VK���tl U�0��uk��k��6"Pk��)i
��0
��a7�)]�q�@�s�9K :�`�OA���M*y�5��2�wA9���E��s��-�H{�H8��w9�Yk��-�������T�F��']�終qw~j'�)H4c���q���0;�X�1������(p��C�P�~�mT��n���*cwc8�G[�C3�c�'�@[Q��ņ�Э��c�_�m��k�^�Zq	�h.j�<�3�O�f�-.I��?���-F;�b-�%�O`�A�������V_^�nz2����V�wq
��k�_�Q�g��J�8��L��b����S:�I�%�AY>'�1`�)_\��r<�M]��e�����6�p#��+l�;96�V�:E�WZ�R����@¸�⪨���6��ŕ��Ÿ�Q9��� �ވ�ȿ^"�|&fY@�⊬"٨فF�*;-5�n��3i*�4�FU�R7�0(G�"�-N!�l�N�?J�kc?����@ۧ��_X�}x�M]�m�d��!�Y��SW���Ӑ��nن߱��<�Nߗh�`I<�8Tv$s�4�_3�\����?Y�d�4bw��"Jա e_\M?�n2>��p����_R$�^w iɥEݫ���F�<�-��C	�i��EQ4�Eof�{-7�	����=@Q^�h�y��oL�=�&y��|p�����I��u(t�(z4cz�ЙKv%��m�
[?F��B�I��ؘK,`1�3��.����#[(��#��j1J�;,1���GwY!�@(��v�3�H�z-��E�����׮�$�I�8%g���s�/�k{�B�C��[��9�>����h�~�ͧsψ݉ڊ�G\A$x|�AҤ?����v�b�g,�U�=���N�[�zˉ���ӂؑ�m���P��8� =6,��^8?�j?br�?�1�<�|�n �08�4�ѩ��2��"'P�*yT�w�Vnp�%��>n9�s�Wtu�"&�4�&�y��)�����^s,�WCe(:��#~�X��Z<�� �I% \ތj�	�]~��CRr�8ǯ����(]x��w���F'�ի��K;VƊ8]U��:쟭�n06wI��,Sq/
��1�Xq�D����	Ο.+�V��2��m���'�OJ>&�$���K�*����&Uŵ<�LШeY��QĬ�s86��H��C\�S�L��m��خ�ᜩ�1o;��܁�i[�M� 
������4A���6n�����V���2�T,b��B_�9ܼ�W %2�w�T���w����T;[�ά�C9�=���!���nm&t?��{���C;?G� �W����?^��@Ӈ?KH3��ۚ�%¼�����L�Y�.OzFh���گ��w�]4�q�<�F��}s�\��	��MX�����{����&Z�Cu-c�f���м�T�A����8��X/�8Tl������o:i���KE��oQ�^��

]0*�n7��t#u@e�@�5��4��z qt�y}d�Fp�� _���D@�
Ԣ��p�ڡ���h�V�\�O���|���-��`�d'�Dڎ�M�Ʋ7Ԏ���5����u�����d=e��?|g��;]�_��$֨��jol�{%J�J�b�O&������۸onTC��%G�1n~��p�Н��W_��������V���\Q�8��wش�w��۔��lNj�7j�7����p�*��%��e���F���n*f�5Ľ�T����nQD~�Cpu]�$�FǠ&"�������=�>�)ڋ/GX�xҘ�R�Ts�������Ȕ5�]���?4:	&ǫ2�|^Ѽ��#Pr���d����6��X�igמ~�▪�)����+��kf�o���u�g�_���8%�\0W^0�<|�������Unn�E�pD�{_�u��bU3�T�sVx$��j�X+����F/.�!Ƀ]���c�ފ]��R%dcF����t�W�7RR�R3A��j/_�����'�ԩ�)9�
Pqkx�A�v�^��ÿ��o�+N���2��?^:�~����ȍ:�� 3t����PךK�/�nȩ X���<�}�4op�,āk��[�O8���'?uv�zSޖi�u^X]��_�.?IЉ�m�^)���ے��ԍ�+x�Ť��-:����QP���p&俾||�S%���C{�FV�(���~���_�@r�/���4�Ő�ő~�,q�Ӌ�\1���-�xxnx�­�����/{���V%ɿ{�{p�@�{D���_a~��iH�kC�_�堮$��!g0���=R�`�{w�F#��\�/Ay_L��w�������.Ns�]���
�o��O��i���!��.M��6�4�V����P�QkG���0��?r�HI֪�:��ك��lY��R����%��0��ݛ8��8�ǹ�ŋ����[�����l �����
o�ߠ�>��L�q��#�@cB>|���,��=yݞ��.å��@����H�r
�ܴ���pz0=��j",�)�����7����۸���⣘�|� ��oZ��w�?/��Կ������y3f��֭���A�:��^���տB�+4/ ���M��ܐL�P5t���seBymd���_����8r�?���C�&|z$ߪ�Y%4I\).� �SV�*Y�|��ikѭ���wM=S�FE�6��XѮ�H,���]R��w�o��?�z�	��ёW~�-F��e�)�������]��I t���K��Շo�/z�u�_&��FPL�^�G��ڹ����zf�eyF��O}�OT��g(=�v�������8�c�e��D���ΑE7tό�G,Pjz>���*1$}��uk_�0���y���i�z�k*��[��3<�ி#����5!K�I�t�t@9�6xi�N$�m���\�k%[�Ћ����d��a��'ɺ� ���a�)2�ʒӉ��R���\&�F"�k�O�ה���EU���Q�?��7E�Y�O�'&����)Ț���&��Y%cM-�j����k�De[�	���Tcv���UJPv�7��i@�R�'^ϐ5��˸��\�,�Oh&��	oh�5gD�D ��P�y6	�����d]��Ϯ����f��� �\��j�e�~���K�֢�c����"�Z���P�Գ}*H�|sչS�M�}g�w��Rk1��jFl���yt��&��y��J��k��Mw'�ݓf����\|���{�%�X?u%c�X�Y�ע�B�;�4r��WI����n�s�@u�$�_�G�2��j�֭ěf�T1JV�*�1@���0sړO�K�\%�����_���2L�ȡ�+i����6��63��)/�G��Z'$Gt��t�J����lC�w�/e����	��"��>�3���$V��/: �8��حN\�Be"�?��2�{�[G�9y��g4\�L
v�V�wd���뮞J�(ň-�?T��s�*1H�NaG��[� ӕ��������g���7�y�w
\�e#���g�{JyԞ;���e�_�E[���2��s�,@ ���a�z�[.���l��{�r\��]2b7��������OYJPc@$w���|��:�Ɖ�i���KC>?��<8y���ݿ�?f���5��mJ{wz�$ҒXK��-q�a��O� K�9�!�*����B5�����/���S�n�����`����돜�)�[bI�2��Ů�ova�]�3�{m���܌v�����K8����[�d��h����+u�z�Ƕ@��ې��2�>������E��^�Ġ�"9Y:x���U�����Z�ޒY[��9�������^x��t����H��k
�S3����ߖ�O�4C[GU��W0��n�_~{ll�)&�ٮ|���,XM`�7�n�S��즡���L��k��I�3S��������.�aE����MB���ƃ�MZUCs�<�&{u���j�|n�谘���'�q6��H�?^�zedF�[����.R��dY9���'��z_�����o.9d��2��dh�p5�d7I>�0�|ig�U�HW�h>���Kp�L���?�`���/�F�������G�^����0r�Vr$��j�]o�I�M���%�tl�B���ٝ��ۢn�9=�?I�Iڪ��o�8SS� �L"C��<A������:D�������uѡ���t.�42�k���4���'y�O�Ths\�o����wi ��ի�m��.^<eM�8�{$&Ӷi�H7�VTJ:��f��#�ܳ-6Y?�=o����37�{^à���gs3�p�l�Uk�4�n��n�]N/�84t������2ZMۓ���Nm--���Z:!:Flp�t�x�L�	fg�A�e�%��N2�B8�x�O��Y��i�Zܗ(��u�4坉��t
t������]���4T���w&�7��7M�VM��c ���ٺ�S�nY���kE���O?�+}����$�c��t�;Q��U>y1Z� �̻s&H�@�L�G*�k��akW{��lnbK���I�%��&g�]��u�й����m�}�<�m@���}�{�y1���/	����[�l�Omo���t.��䧈���[��2�Q���d8҈˽����~mT���(+��z�޸� ݟ٘�匦*�d��}�;��D�K�������R�N���5�Έ~��m��1kr%;�#J�i�3��|�֩��I��̼�A�K��R� ��
 ]����T@��b%�?�Se�5M`��G�'f��vo	��f�_z(�..%�����a�c����S�
^�����R��|�(K�)�c��b�zo���N*B09�=!�7��<߅�恙s���|�g���C�P��r���a�7�NQ���m�OI�]h�;�i<�n�0^K��L�SZ��W#��Fŝw̝C��r0��9�F��E`g襸�����j2�[� }�w�ؖ"�7�s�w,�Y�Dl*����"�o}&�ܥq�%����S�?p庽��qq6�^���]�9'��[�=D}28��ϛ�	ϿJ�^�g�ʵ*�S�c; ����G4��5K`����(�麓ue�W�ӻj��ft_K˚��TM�t����N�/��"$Rwj7��@���\+~�XFR�DPbN�&LdQp��#��|�s>k�;���:n7G퉜����f<pt�^�{'�OI+\ck��P�ݙ؉s2��S��L�C<eON�٥:���\Jk�z�x�+��i�H����c��Ƿ�3����R��T�f���l5p\�?9.M���v~7�rS~*r_|�UG��e*���ꂉu�P��������H/�`��Q�ͩVY��ƥ�v��G��dA��F���,�{���>,e"�3h���X@��y�p����}b��sڡ���IOS��JV�d��Zm�?�^�{ˊ�y�����[�������~�l筫�W=E[�Ug┫��A[7��*�'=��.�T�X;��]�S����J;���A��"H�he���	N"�����yM��޻n{���e���;�f�[Ug�
�q�=��q����ڝ� ��Ά���s&ץhqW�n��YK"FV3�3H�^�*��8�_�0;cr����Nʿ>���4�H��K��`�Y��KD�6�Jթxs0�B)~ޠ�AB Z�������'i�,�O��|�[i�m�޵�؏�&sB� r3qF�Y|Z h滙H�c�e�,{�������s;�ɻ��v�����s���L�H�@7����. @z�X7�,�����z�*W!6�O;�n�Ԯ��8�Ӻ�!�ш(�S��h��qT-<����?�R,���w~s~��!S�.���U}�K���fLǫT�XU�8��{Yk�"7�F�rw�_��H%��gE�>y�E�i���Rz#��K��[����TR_���F{�	-"b����?�N����QU�R3���D�׏I:��Vd�,'�Z�XY�y=a�,�>�2n�?��]�.��iv%&��I�.�&��`�R�m����Bn�~�k��I��LG?�|�	�qd��C*`��nd��+�7�dz~����UX%؉"�ݧ����KMU��w��ț�pMc2`�l4ǭ��0ʩvA��ϡ�ݴY�1�dbV�~�#��\P�/��*����E�
��ܲ�dn���-N_8�����eFX�9�d�Pb��m��%��ր^�p��f����>��"q��DԮb�"���@#:'9��A�s%7�����9ޜk�=N4�//����$���+?�#A~�b���t���2� 	����(~u����@���3���U�/���y���+��hL;�C܏�m�5�F��A��%�1uo�0lE��׻�3��!z'G��L��d�ނ'�XnL݅��َ:1�:��1����Ƃ�3%� v痙�%���yo���b���������M��	�|�y����\�H�=L���'إr��U���1R��e��� �T��7Q�Q��f� s~��բz�g���ҏ_�ᬁuؑ��qRb[%�\�����K\pZ���$X΍����""Z�x�ַ붙d��p��v�_)x�	v�Y���|�y�u�����-To��L.���}l��lL��)�&����aA[�H�i��Q�viǶ`� ��R�A���|�.@ܴ�M{�i�5�d�dU�������mt�����u+�2v|L�6��Nlnf'`��b跥5|�Λ�v�n0d�}`#�05<�~�D�9�i��ì!9�u�,*64�*L�l/h�p&�ϑ�@$��g�1�m�&Żm�������^l����m�����`�4�cC�#\;W�UC�������18��@�-�*��m�:�vp �ON���N��������K=����%!�3�_*(�[��D�V����"�(�m(#�:��./�ER�s�{�4��K�����FG��5
�N���Y�{�^<������}��q���0z�d�=�[h!Gc��ЎeA��i�������G��q�
8�Jf��$�������	����)�B�b��=X�^R��a�	6�(���&�vm����Z����2�����6��V� v�'�u%/goo
�ݘ�ߝ�PU�;�^5�G���w��[ї�!�ka_
7c�O�St�)�g�	�1�^��c�$횁���������k�+�&aa�tG���X ]aL���e�����c=өr�ݼ�n�w���zP��횵Dʨ�/�QR3)38Q*�	\�}U���(!�b��L.�sFNH�<�/����*�
)����d�����.(^���Q�ܮ�[<d���gؚ ̉���n�с
2�PM��{X���0]e��Ӡ;��ʥ�� V�:m�iH��h�L���Z#�S4}�Xjj�&�Vۼ*Eu]��#�u���n5^�0}�E�V=/"m�{xh����oKmxx;�?6|�,8D@v,��N�v���n��?�͗����UE@.>&�Y��-?>u6
U~-��l�� 3��Y��eK��_���N��{��yO���@�0���&�w|�*���֨ך�yWGQ�N�����u�n�n~�I�!����������,��Ð�[N;�����^zi��Kb�û�F�{c�+&h/�d\��Ű�����qx�\^�.�����e��Є$�ߊU��.do��҅�V��dP͜Ax}�R,]�VRQ*mt�ѕhE�Za���[�j�X���������_vvj�3�*�tf�ٻ�� 0��_z-�*\)�e��k�8Ͼ䄖h��g(W�0;\�2)�TϺ���ׂ�霰�)�ـ^�5c����`Z��pD)F��P+�z��[��5#�A|�M��{A��^⍥�('T�|3��S���[�t]��_��N�ݦ��H�c�=t�5�i�u�Qٚ,L�SV�~?k���^�!�.��~��6�_�ɗ����I9y\�X�/�r���B��f����.5�o����g|�c=�.��$T����q�m����I���$y_�����2�����b=ݺ=X0/�6�Z��+��2N�bN,m�܅B�wS�V��Ɠ�o�w�<�a�JF��r�Z)ǆ��{�gc�3OH��? ��;wTq-��D������%�8&{�	�c�p�h㐿<���?�tqY�|hn�+��ԕ��HhF��m��j8�^�IR(����s�ĺ L:�[�c���ݜ�3JNىfb��NЂ��ٱ9z��]|�L@�h�z�u�WP����J�o��H������eN2���5��:��*-v�e[��W��7�ϸ�ҳ��Eo���E��H���.���A.o���O�C�s��E�}�h�M�_L(���Nu�"�&�5֟?훮���}Z<�#x�q�d~*3+f� � �,?c`�Ȇ���(R��C�xo>#j�zs��>Nݘ�U5+w�Ml�t��-�Հ��N8AK�jp8{��0�R�c�/o�+���e@Б��
�tŢ�ُZk�O������
�n��9Iާ\~*�yw��7�L�h��_c�{��W�Mc!kreg�|��`��g�
��΃8_�o����Y~�7md��v��x2����{\L:�g#�_�u��8���=���`���u|P���a[��ʬ�Ge����s�%�>�0!Xs��������D�IOT[F*�o�0(����%wc9�k�(��>����}|�y]�+!�_9�b$��od���Y���G{@�g����4�xO�Զ�`j����1c?ě|M܂�O� <��SbM���ΧU�_+mF��|_�i���	{����Z&���<'VR��C��=�z{�!�+��.���)a{ݾ����i��U�sĝ#�pS�X���0�W���e��qb;�m��ʛe�_/�S��.>�/����֐CX%����z�[Zç�!�>G�~u�����ũ�M��餵\_}A��-H��'R��2w�x�i�}=p��0��m���@F��/����}6�~����F������n��9��XŞZ�ވ��kW�b"KO�eUlN"f�ě@� �q���ͭmvGYAX�xF�^�m#�bgW���ߊIG'�U�Z�����5I��Dz; ���1�U?۫F��=�_EE��6��J�����;��U«ׯ�o\{b��*�-pʴ)�3Q�K�m2�WP�'z�}��'��Z�ݮ��M���-���H/���K�I�zLF�yAy떾��5�v�Q�׼I*��� ���c?2�db�R����fwN&������'�9�{:���S�s�^wԛ{6r�B�p)���g����4v�6X��F�0&�S	������M4�|V�{�����($oę�@u�=Ǽ����8���z�|���3p<0}�����K��m��	�PöQ��|p��ii}=��g��[���@�ޢ�ީ�zթA/�r_�޺7�}9�1�T��v��7̎��ov�pÚ�S�P醾���Y�)�%��Q�s�g�#HZ��d��o6,N^������.����|ek��jU�� [[&z�D��:�u	x�l+�+����鄗�|>��E$��e�H$�v��$�)����Um+,�/'�9�E�����+�}Et/G�����dԻ���7����2����RT>�?r��lM̅g�b�~�����}�I�_�z���G�9�Q��_�2V n�����(��U�4�nQ�
/��k
DXE&��s�X��N���Ac����w�"����2/���jJ�йD� Q��+�q��� \�n[���xw'b?;t=(��PL�fX4�n��k	q!��9�\��ߐ���|�Y��P��s�/��e�k�g�5\�|l�sf�0�k���4m00�] ��܃���rt�R��	��YQ����q����׉/��WR�ڝ�D�.��$Wب-Dl�����7�������H]{ZK�<������7�z?�ZDE��q�D�*wo�O:�����v���Zk��w�r�2�V�a=hLV���{e���>��@љ{��L��,o]W0�xR��i��gg�����VAro���")��a���K�5N�g�r��hg��r��k%J�IsJK�\'�M4�m����Y��֎"&u���@�zbR�i�|b��@e+�H��#��#OUy��&�N�!b�����F���䭛��lL��Bay���o[������d�����������Ks&6	�Ef�ܰ����A�&g�j�~"j*��>�"|9(u�)� �E.� @FRo�M"���28�)=y�0��	�*�3eC�9��yWϔ��k3���x�Y;O`�x��*�={X��nb�.b'<��jkd�R�!���q�������m���k�!J֫yށ�)�,�v2�*'���s��Lt�[AVVKmdR��!�����~xs23��yx��iK���WmPid��)�c.�%�}�$ǫ�����>o��j��v�ɕ#�V�
�q�
(JR�Tk��D�ü8�*+qC �S5K���;�����8a�8�*l��vz*��#L�PYD(	c����\�|�,R(_���x݅���d84���9�֩x$�H,KN8L/�R��6�;'ϭ�y:������<�S#�Z/B�����+6{=ھ�|)�u�^>�d�U��H��KrdK���o��!��#�p��7��ze�yh�"�'�������,V�D4/��W��Y7�z����t�t����V+d [�?6�0T)ݮ2�RYw6K̰_���W���,��|ˣ�%W�S#�Yņ���a�����p�w������ZK�j,� Y����*�u���<���t�F^x:o�w�d�ڧ��d�͑[v�K��x�`��Ln�~���"��r;��k[�;곱�r]SL�<n�ie�z�#鑬� �?�5��O���pQȮ�wC�J���������HM�B\�{��ΊY��tӊ�x�E=�#�G^r:1��x!D�[�g��$\�Z-]���J�φ����8�<�4��	�9*&Ψ�AҮ�Ic.0������)�p8�N`��U)�!{�E�Z�X�C��8�G�2<[�J��_���B��G�~����|5�U�ZoWm���Ҕ�O���i� ���O�^�c��i'?��\�v�q:`R���]� z��P�*�<�Ⱥ!ۈO��
H{D�C���sb�j�os�A��PwgY#*���\��l��Ul�ya�'y��{�c�F�_������x r퐫�Eu+���"|*]6���e�Z]�#��@-�}X�[���z���ɥ��#�!'i}�|�T���ɂ\����H?�E :I;��r�s��Bˤ��>$^�1h9hf;Q8]m��Xr����%**@^�ϋ���on�bk�Q�j>�)��h�@a�^��W�6���!��� >&6�Y.P�-U�i$e2>��.�NܿO�P�.,'���C��Q����4�5, ����5�{��!�{��oƿc/���K49�]���8f_�{��M�,���9��=�@������@���Ϫ���@��G��kӥ7H٧�_�,��.In�������a9y��AV��.�3�*�;.��Zݙ�c��<	�Sc�a?��Ո�t��d]I�MpZ4��E6�Ȁ�}r�d��l��Q�[f�Oͽy3X�Vldf�ɵ�
w߿�����6�Kzk �WE�~�S�Ѝ_���\��������mg^����PR��!���3e�۟VM����D�5)_�E���6������l��@���7ԧ8J�G��Q��9O��en�ܯ<�?�/r�Y&�Xlv&�Вs�W�ה��a!aur���k堖T�@v�$�#��]�!�x��O�Op�m[���5��0�U\�̾�˪�7K��u���S��~�{[U[�h���SR2b�]�bo�T��cx��!�)d��������Zbzf�}��sw䱍��(7�֯%�����Z�9�$X�����"�k?��W����� 篋���χ�2���DEG`F�R_)���y���y	Y�À�vP��'oɶ2���ƀx�Z�˦�K6�!_��Q�e�|���ޚ��n���V̑�_�G�yvr~&0��@шظۀT%G�o߄l�6W�{��=�=�>e��))�G�~��.��4�3���3 #�WD"G�Ѿ�����&f|cƠ�/�F���U���ط�S�����2C_*R]�{u��o���9m�1ȩ���io�y*�� J�Ye@�6�E(��iHS��8y �^K��N���*�Q���fS'%����H�x��[vx�ª�TQcLíӦ�u�aC-��풇�b��=�+��"�ck�s� �5��L�M���[���3\g2����{H#��VBt�Rw|U6��t�,A�JJx>���2�"~��T�R_������^5��eXY1���<Pt��%���O����!��������{G7��0��O���)N�������S7r�y.�E9S�}b8��Z�,�h�y}�u��^k~M�`�6�����D��bt��9����R}�Kzy�wב�Q�0�A��7�&E���Zƀ�$3輸�~"ցJ/�n�F/��A�EL	��H3h9Z�Fp��*��3sw�_'�5�?�x���c	ڣb�9��c?��JX�]��TRup)67�����yiyʦ��z�b�醶�����ܭ�|��k��kq�j��X���,�G�g�Fj��>�ICj��&?Y�R;��sH[}���ƙ��T9}'����1y��hת��U7u��$����I_N)$�.���1N��BN:{묂l����S_-X� ������r纖hB.���
��,�V+׫��F��.�%��\�V5�t7oF��<�(�9����x����E��B�/����rj��E�����!<J6
���|��	n�IAq�m |�S�_ y)7#P~�ۏ���;~������&���b褽�
�x}v;���,gA�=%l�Ŀ�LÐ=�`kD�R��+xM�+�� �k44x�
�ɥ"Z�[���r�<+n�Y���[�.����e����-���@ ��o�1z�ھl!G�y�0� ���&����/1��f\�IH�M@��]�G��ԏMx$�\i�nSM��Pn�iv�N�녎�c�%?e~Ҫ�*N��&���W�*z�#������z��Z��Z�����*�Eyr3�9��Q'�$,9u���}���MmG��]��=4���%�E�Ʈ�􄾹��n;[������]i����,v8嫉�yHa:pj�M����K'��E���U�s��:s�{�YK���֭�ukF�S ���94e���}^�}�1S��SA*VN�sT�о�QlH��ܡ�!�[����!�H�<�o�Q��U��C.v1
r��~S9k^�<�U�QB�-��D�b_!�O.�P��r��vBm���)?����щH�F��j���km�tY�R���� ���ڇGPR	AR���T@����S��niJr��;�c��a`����+�������[k���מ5���teW�^fණ�I)�
�柌�)ƺ�z��&�|kň�h���M���@�TXQv+>���^l�����m|u��"��ۖ�Ďϖ[�j}�fӳ���2o�>+�������|�&"����͸��'ݩ�3��ΑbQmפ��KD��������0ðׯU���r�(s 0� K�q�6##������*�����$#�OIM�JN=�C��GחOV��hW���HZ)QP>&/����`�tHZ�[@�_Q��Nr$�dDl(IH����%�-�K� %8�C�[�J��U2��6�V6��_{4U��%��Bkd: ���2��j��w~�lƵr���|z��)����l�2`K�O��3iSp�ސ�Ԟq̈��.��p���(�ϼ�k(�-P�Y=�k	��+g��+��]���	��)3]���쎑K�|J��y\nh���c�₭9\�o�)jD�ՙ�Udl�O��;I�E�~|;f����Z5�9K��oǋ���'`?)����S@�O����@�S8�~v�D}�J�k�Srrqww�^%$}�P	��o�I���z�[�*<�x��/}�S�j
~S��>�Gd�fٞ�l�hv՜���G�*9�יmGK� )ģ�%[�O�JFy	H���|%���c~�X��yˣ/�>m��|�X�!5��Yd�%��깿��rVt�u4J9b�w]��NZ��p�,�s 4�PI���쏢�*�m�����?�1"��|&eg緆M%m'��
+�cs����������=��'�w�r�x�&�i���)#C�s��|W8��v<}����d�DO��@7:��Q���Z�1�g	d�܋1�J'Cx�p�?��ѱ%}�v �� ����U���,\;�-�l.n���Zv ?`�"��ܽ&�:�d��3�Y���-H,�q�?=ԍ����J$���X�w��y�����p��kM��{���\�� ���0=}L:��`>Z��X^rvL�4�-z_ȁ����p�íqdrz�Y��.N�CL��.�**s�<{�፟_����F�x2���		�!Dr�v%�YT"a�p�����R���D.y���*G����ۇݦ]gK@�d����FU���l��>wV4��`s`o�����4�e�'[Y��ߣߔ'�z�C�?�u(0'�L=tpz8�v`�6�i:�'Ku��;ҮkmD7[Y0�O����M��2E�1����-��Չ<��/�f_L��&���e�j,�*�n:��er��9��7�
G�������rg��0��뎙�����픏�|e ����o�?��A��"��ɇ��5H.A��!`�I�d��t(5P#�2��SSk�&ѫ)L+v���ӄCr�w1]�d�.:?���In<⡦�M�����	k>���5�|�F�&�(C�5Yr�@Fr^pν-=��������c��?�g�<BN���o��-�?Ƌ��Qf���o|�m�����o�vFhp��|�R�؍\lX���������d�K�Q��m+��_1�$q҅<��ӘZ���-�1� ����p��o!<[](æ3�����a�ɟ�(m���ɗ���܄�E����}���c��vR�"�'�5�/���?����n� �&(�H3D�y#ʃ�WQ��Yɗ1�0����/����)6�:2e�	��.fY �N|y[�/�^�[5��gbN�V&0ok�6T�C$+�@�J�W�Eϯ�)����]���mN��~O.n��~S79��1����f�!��D@ ��p��>!��zY{��[�����&x�/'���V�k��Q�Td8\��b�Oxy��~H���f�t�9��n(�+�W`rF���@�!�b�P�)�^b{ �GaL�-��N��F��b�S��1�Z�v����3���699��5�RP&�p��;_#����o|�TM�7_��z��)����G(�m��ֽ&vR����^
�LLO�5�Ь<�S����n��Z��3jW���W�l���@��Ψ׮3w��J�k�?B��]H�枋�WG��4��Iݧ[����� �����Q�_�%cӌWj�����!�����u�v�%2����&��"��~.�2~H6�.9�aW'Z�~L'b�;Zr>GC�&�J�/�w~��L�;:�Hj��}<����9���K!:��¯���äA�n1�9@��������
�)���]�R�%���K0��g6^�����x=��*p4�]�2��i;��2"(;Yi*\�׆W��^V|̤��N��,�q,n��~�mH�8��H�p��r4�<�;�\�
��7m�Y���t�ɦ̰��E�S\w�~}\7���S�\Jݑ�o*�^Vu��.�v��M���O�:�P�������O����Ս�|��TE[\�L\�N8Ƞ��5�h���ì/��뜍��BE)�װ��1A-C,V�rѽpxa�h}bc�#j�q��"�*?etV��yV�D My�����(���6���O�d=�i���<��҇&%;������v�|~ɵ��A�ށ��츛\�U��,_�u�t�l�`�y��^���s{nA��ѳ��O$�����$���=e�}�,K��=�*���~f�`+�io�tk!"�?G� �D(��[	J��IDÁ��ٺ��]�g���ri�l�;���E�;s|ő�����Y�����2#d"a�`'���ec1���B���4�3�Ȁ�\��lc�b0�v�Z�2q������8�א_[�
73�#������c�J�-�!���'���u_!ӜUP�J�ڮ�8:(���\��B�1�g�zw1C�'J,��Y��+ѰM�-'�VH�Z����J���
x20�nh�B���]42�)�v�҃��h�ە@�� l�s�_.�}iv	&:D�h_�p�PT����)+�T�p��Y����?�F��Rd�6��R��cr��[��DpD�&G��I����-GZ���C��!�-�e�/o��D]81ߑ���� �+�W�Y�56g��`*cR�g&]]Sg��O��}F9JP¾|�U�[2���ƃ�c�KĹ�Ҋ�E}cezu�	�_��ɏ�]ޝ��7͛�l3�{,ש]�,J���ߦ�>�gXߠ��D�Զb���L���(���-�� ���Y����ڳ�Wj3i��������H�c�H���7�qnu3�|�ւ��/'kM7c�MX�:P�\Ø<}҄�X�P���<*"���$�'؇]h'��Z��H�>5��	,������i1�.T|=0�+7{��Ӱ=�$[zջ;��w�6S��|���%\�3bqz�'�r�(NY��Y崾��z�=Q`Z�O��pc�Q�ȯna�Z6�����U�D�4+�~f�A��2�E����?�G��!�F�f��������^V2�_?��8p'~�����W]Brv渚�CE����_�ۥ*��|[b�H��_�p���e�|��P^�����P��Y����0����*�� ĕ�hH�s=	�>��/�R�1���&Y�|N��[�;�	ed��p�̝+����y�J����|ӳ1�_. ��K:v-��b�*��o�aUKs��5���ry܆�Bo���/�m�M�,Y4�B���ՙ��q��퍑5X��&ЪL 7e���ֶڎ6k4L��]��D��K�L6޶��z-HEѹYM�#�'ڂfٶ�;�\��r�W�H�SQP��bb��$T�)�?L�n�I�Xu���9V5/����Ef��#0+P&�O����<�9���o�c���W��]#�l���潻 ����Y39̎P�4y(ʆ{������x%9�v�a�*0�j-�L�7�Զwxo��w0E$R��<�K�
s��������ax�xӖy,)!�����"L_�z#�ӭ֌_��ٰ������Q?}?yr��9�SC�\��yj�|�Iz�P8$�&l��F)|��"�//y���(�M4
~cjjl-Q2#<�$w�#��U�d�Uj�UA����� [
1e4�[���?ⱽ�~��l���8	��7�[��/i�8���AZ&BC̛��<��ꚝ|�+�
�Y��h�-u4|���O�PG�����?g}SD?J�"�{@6M����Ҫ�	����� ��ǁ\�ZY��c?؆�]/$�&�{����l�P�u��1p�Đ��kY'���]B��w3�(�%�;�7��X��̑u�1�N0w3Y��!j�.n�;���?%Ec牓�kk.��^����E���W�m�Ѹ��wo�曦� �����϶��5�	�5q,�2S�����s�/����|�����4��Rp�/V��2�y1u�@Q@�����pp�p�ޣ\��j0!�Ķ:\@.05Q�ނ�;-��~�ʉi�V��7{!�i?&����=�5ۂ%^1�=�V�8��jԃ@�k���Pm��	uRK�Bn���-��?�he]�(t�8s��Z8���d�:!Z\օ���H�}�`tt��f���(娊ʥ�J��|Է~Y�ᔞ4�'^�
�_zq[n�c��XX�~�||��"!��5�*{�VL�c-7c��5�^��;:��ڈ%�aK�s��I�e�%��S}AR�R1?��[Km9�r0B�p��U�D����	y�[����w���K�؁4bL�گ7�U�[���!��V���12K^��tUQ�4O��U*�T��fU�{́��A�c	��q	�o�ެ�E��U�LF�y�_H�>׃��s�P~Sxn�~l ���*�LN����ȅn��	�E�QMr-���o�W0�o[���\���VY2�~�B�<N�o"Q�`�U_H��OD-1��$﫩�r҄�*�!x�������dM;�Hi��M�o�Gl�yB�2����R���\M�������\����'Wxֆ��ɩw���+���m�����^!���_���<c�?�9Y_+�������S����My���~ŕWRzs�����  ���f�F���,������;
]����)=u�)�D��ǭa'b%�Bֈ�R�5���T���N=�L�=t p�Q5ð5׺���DOD��K���t@����3�A��Ԡ
B	���2h�ʟ�G� �>D�l{��.xR�+�����N����ßN'�Ǹ�E�R���A9�������yt�!�_qE���҉}��Yv9y��;��^\��n�S�� ���X*��r��d6���{g�����\z ���4!)i̳g��2�(�r:��)=���a��7j�����r�  �'�(ٵ���ۨs?����B7(�kd�(M�ma5l\��z���̕ �߅u���◠�z5�E��3�K�_(��rAGJA�os����!a%~<uvi�  �� 9 ���*w�O�ʦ���(�va���zZ+��%��E�nUޛTSb��.<�*��8W��fP����Q��a�miE[Ҹ��́p��ʇ��7�W� �P�
�L�����՜��$�Lֳ����$�q-�|�c����ع_/W2��;��#��@84���+6:[Ţ(U_]�u?����
�} ����^ں�EQ�N��PW$����UH��R�6�H�]?�M��m��K��[���r��8��Z�il�p�.P@��C��ɴ��;��@�p�"���(�) �T�Ȕ�$�R��Uo��"4�Z~�I�H0u�o$�Z�M7�� P���C�g.�s��S��X��0��S���]�)N�K�x�4?��[��6o9�q2�eV�Gv�ƩC��n�6j���ܵ�rQ�-�����$�F�I&�U"�f�+�,��N}��e��x�Jf9�5*
�8s������]?  ���e��at ,hby�-&Y��r>W��GW,�;�,�d�k$�޷��!v\e��S���q6~򇀱wX{��'�J}����~�*'��.vNޟ�,�3�RO��T̏�,=�o�� -�K'J��s��������(ըI\�����B:��<�zt�yb����T���@��:�Eh^B}^���sQ_��W�����/���xH/6M��@��O$x��F۔%��ָ��[�9cG���7_�!��|)\��\t�x�c�p���A�gZ����u:?�܆(͔!�wۃh�n�ʂ�s����*Hy�m'��ml|����noҷ���eJ ��n]`��z�[8�p�c�?	�XJ�#q����Ul7W�﯆��.�h�M7O�MTZZY)"R7j�=aL ��:L�p���}Њ���槼ը��	W�CBN:��!�xiB��1��&>��+��Ua���=�x��x �	M��4�� ���t:ޖ��d��Co�V��+^���ӛ�\\Q�I{Y�{�&���bB��6��#]�D���V��T �`l�(!�����R�\�� �1�1���v�E��%w��2]5f�B��u��e��^�>"�b4���h���[N����D)��� �.��'�I'@��0�����6/*5�$?����\���Y�#�H�-=����� NE��s�K�(�]� q;匦6q~�n2�&E�]~땕�ڛ�xD$-����7_β�x~���Y��Z��A��O�ɛ����,�s��-j��B��4��m��ԃ�aoS��J��۠����ܲ�l���%�Xز��w=t'ݯb}�(������}Wf��	}KY�+�>��h�>x��_����]�
}��SW"�]rC��.� Ȉ��'�v��
��ٴ/辟-	�����;��ԍ��U����c�q���+��0D��7�G�g�!�"y�]�g��3���M]"�b�7�C�農�j�ׂ0���{�f�>W
#茂�7��龫��8�Me�	_��wώp��R���9I_�4潉���p���@�T�m̜o>6���v�Y�h���*�W�\���!vd'��;,p�Z��+8�]��<
7���D�3��x�l��N��/s�4����[��5?@��U��z[��>��#{�"��x!�k���છ��c�[�j�9U�&���$W����%�@O�8&�c��W~� bF����n����ƪƆ����vm�5��lN�T ���ns��.]M�k����{��:;
�V�М��n���em3_�y�I���4kcn����2y��Z�$\�i]�# ��8���<�#o#p�*�2�a�ȇ2����\n�6W7�����u�쯓��e�'!�6�7���Zg�,e�?S�i��Y�z+z�
��Vm��?%S41�蒪����9:3����@D�����鐞n��s,�2.���N���UX��"���8��k�f�U���xf��c���|���T=f��㕌��b��7`�8v9��������GQl,O��4ld�s�Z3c�/�Hqg0j���1�e0��as�:���i�9�I�ϗ�~��å����˞(xϚx�J�F_/՝w��ߡ�I�F�s�﨟:1ܪ�� �=cU�-�z|b?%y��jm.�g̜��t��W�#al�����dE1��0�A�Q b��J���ugT��"O�����e��+_����n���q��po򶒝Z�Wm��X� Q�CbN~8I���nx^ϭ�Z���B?���ǫ����A,�[O�j��	E/e�P�y(���ǂ�S|�"ώa�)*�S>�Hѱ������MC�&+����,I�SO�2�̀������칑7��6�7G�R�cfJ���C����X�)vK�~����$�#�c:�G�q����}�	���Y�QI �g�b{��D�]R�]z`�\fK�!����'EI�C ���_*�b��H�Ao*Ф�S��آ��uB)���A��
 Hn��w��cU�y�-U�Z�L����h�ߊV(!�[�]��h���>U�0��y^�kzt����t=lWjtuA2���ξk����,#k5w��n�z�	���qD<	�/Bv��w�-5�Q?�u&o����N��j�]�[�M���"ӄ��-_c��[!�����m����J�<���?E��(�Ɲ�5	�hZ\��1��y(0>��g 4���l��w��  2�v��޺ӎ[BOm�2=�&����O��?�˻�C*�wf�QJ8�e���hI��Y݇ˆ�5��1��|S�&��5� S*r#����_{LcƮ&�Ve��֖Y�I��.l����4R�[�;��h4�j<Y?�m}�t��@WU����c"��eP�M����|��6��/��{GT�1�F�|n�3��5��[SGtB�;B�(�^�%X�	��_��,f�s��b"�>���V�X��6e�P�"��x
r,Q����P���~�J$�ɫR_$���@y.�e�(a�O�wU����$�ԋYwy�p�>yD'z�e"�V����F��יy�^WpO��J�Th�Y�T^n�����Vd�?s�������Z.�\��'�T�A2o�6�G���ה`��r5]'�t�k����[-��|�fMLA�����Ŝ�����o�K�����.Ρ�
�TOx�oF����C�bP]�W������u�p[��rn��S��GXi5��`�+�m�ӆ��6l�H�u���|�E�J�{�)�le�+\ꕩ�*o�z/���y�3�� ����PG�iEκZ����[�`�+h�!�}:1��o� DHL�"�ŉ4�P����
���do	����	�'^��YY��M��cu-��Oׅ�`�97�hJ����Y�E�.C�I?�7
P���Q�y����;���W7�!����8�B�*��n�H�	�G��Wy\����͓|㡐�gi��&���9�\�~v�ۍ�����f��L�BǷD��7�����z(��Ex��尐ʩ��tw��6J��As�'����b��j��6{DW��skE�۳��O6�'DO�E��I"]V)0v��j3*��%v8�߈�=Jn�T�'%�.ADO�1E@�~�v��S��	��{�,;�V����qPiey;�o�K��\�P�N��"p��5��>xq�o�w�2x)��~�׵4C�-�t���h|F7��	��ьI1�I��'��$a�ߵF�س~eA|帹�T؇O�f��mp�6��	�AE��;�����T[t� �PU��S'��7�l��r��m$�C=�LS+Q��=�Z8�7s��Ι��/>�{�O(X�&,�=j㽋�4o�M��|�o��*�#�]�䇳���;)���,FWUW$�ȺW�d�3U+���̫�v	��6���*r�Y�������eB�&���6M����$>H�ݺ1SC��,s��B��H�jR�kA�=e��}�d�qW�0;]����W�js5���"����y��؅��n�kZ��'���	W�v��
-��s0��E��q�D�.d͚c)x��'c�	�*�,d��%w��*�;�xK�U�76��u���c~T8��%|R�D䄇ԔB�<���d_��f��UHۓ�5�slC���=�	�0Mq�O�cT�'M�$�So黫L	]f�2e�����P!O?�5���o��*���߭`�\�g����Ye__;�H<6Gة�,Ļ���5o//j�k@�#�N�V0������U�X�s���~fbǛ>�u󏊙U|��9��bgȲ�qe��MZ�\!�Q�V饽�Nn_��M�ަ��̡龪�y-��1�.AO�&Lt��ܼ�CQ��0ڂTvr̀�o�r�/�Rj[�-��n�鐘{�5̂z��&�F�g{�4�:��ջ�c��`�N�-�!q6�UZ 
�W4��i���q"�,��P@�������W�_Zh�$��l�˕ᐳ�r�:�v�@z�ؒ�\������!�6΋hwl`N�iݣ��+⼰ȾU��y�,���`ui��vl~>m����Ku[X������R��[jQx��ӻH��J
ۚ6��l��,����KuD��'�EaM�!��|2�
�Wk�;����AŶO��K���8|��9 ���Ua/q�y�"rT� ׳�E��UZ��C�K���f\�ު�|Y6��h�N�@D���C��Hv�V�h�2�O{�
-1N�7��"��+@X�F\e���l ��y�B����
�1hC�{1��\,�
8��	�H�J5��vPw0��}�����x�}���C���C�b�ꅺ�v���
[ljv7K| �p���1qx��գKuCA-B�F���O���}{}*lZ��F��6���2$���+� ��n���!�+	�V3�EIxȌ��mi�6<H��]�]'�
�,�Ix&��י��N��8%rO���t����܅�d�L�4;Kq�.O<�t��V�����:,P�\H��;w��ȿ�cC�j�ww[$vMA����?�I��&//O�')�x���0 ���QA�m_6�>�o��Et�ײ|bN�i�l,���k�t[��X!��S�tG1�ٛ�안}�	�'�d��Ϯ�g�KrB�A�Ovvy�9c."�d=���1��;!ځL_GoƱ�������Rڋ���u�8?� h��i�|�:kS���>\80ڲ�6p���ڧ��}�]������բ/�/�S#xc�a�ox�8=I���)��ɷ��\w�7�8�P(��W��
��m�\��y(�8W�5Wu+�C���b�3�%��yk��Vm|bn`{s�t���E�9�[�@8Wa��OR�	S�	���)���m^[Sb*:����� lp^C�8���!�3�T� �3�	����n�e�,ݛn5B�� ?�� �zrP/K���h�4H�{�y�(�~ԅ���q�tY3M���|�����ݪ���Ma�/Lj�u�Z'!��lU�����⡽�%t�HocV���]2H���1[%�����}�KT+�\��b*��M	5�n��譔���f��Cy�{?v���Ԕ1ѐ�n��"ﶲ^�`@Զ_i�c��4l�67o���e��I�X��Xg�7�u��m�\���	�����J*�^a�=�X�$b7S�B�)+�Q}�)6���n�d6���e_78�	;��C�m��Y9H{��Zw����̲�T��cK�C
��;��R�x#1�`��X���o<��A��������,e|�{<�>?��+̍x�>������z�"��F� e�/qN*Jy����k�4�c���g�B!��>ۖ��VQ��*�'i����[9���{��h��d��6F�5(�IN�X�*�o���.�f{��Y�e�Q��m�����u��p��N�m����WO���U�4��K�
��gt��J��:Vե�����=)L���>+4(ZT�GOV{ W]�2�4m�dN�!�4�����?M���t���ɒ��AŞ���=���sIZ��ܧ����qd�r�Ӹ �)�"��8��n�=nV�2 �� 
�zچ9"��@�� h$�\񳄊��9&�)�РL9ߟ� ��}v��D���z�ؽ[<�zk�.7[����%�b��
��㇊=u�ٹ���M�wG������WM���5��f`E�� ��$�MO��=�0�-�2��_z�Y�("�29��U����~c�Zu�J�����DQ�n�5{G�I���1 �X�2�1~K�î��14���>�E:�v�IO�1c�c���RϽ����!-`mu�۸>��$�MZb���}��<�Z��e��\��v]nԗ���3��q�;�FI����^GG�||��P�:�WI-�H��nظ:�PVf\s_|���_(K�Hc�����Б�A�-({�uGb�Df\���H`���T=����3�� R��剩b��T���K?�D���G�O�j�o�8��R�����T�а��s�(}�Y���[�㖤��)Ĥ��"r5Y[.@��M�ɸ��r�5a8�)�֧Y\�=J�G@L:���m��(}w[������E��Ĭ����]��b�%����bug��ܯ(����M�8^G�D��0��r �"�r�76I���W�0�����;�C����G�N��
{�l��B�����a	�}b� �V��4�G�<��h���䨀���p���%�����
	�HAz�ˇ�q��b���c��FJ7|�+��ӱ�"�\o�Yx(c,���Lu�Ѕ&�f���p�V�!s��E����o,����SJ�5��)J���3J���/�$v�Q�z�0XT�e!���>�72�8�4��V�d�-7��p�6�%���:�ؼ��o�y2�HpQ����P9��h�'�ֺԏs�궞>i�k��妬�]��Z�$�^�4a�};y[��ydkq� ����n�~�\�"d�3�_F�B4C��87�,��E�����á-k�{�ſ�}:/��t�j�/����*5)����ۀ"�~uMN-��������
���9���+�����g��q�P'5�~��;��EB|>W�c��������6���p�}������t)`���VC_��=�GAkSl͒�3O�5�44����!H����z`P���Z9�-_�[�u��R�+�d��9ޢ��f��*Q�dC�ၻK~� %�i��	y�~��W�V��d8s�ϟ�� ,!��|�$R'h����ܖ�҂E?�%m*Mr�I��pl1�]�jTq���ɯ�#Q�������H�#��[W�jh�X���������[@�
���m��ɩX;٫�<s����*�\�r>)J�
���&)/O�F�A�6x���Y'oAj�1�OJ���ـ�����l��N6�Z�1���(P�����^��=��ti�g�T�N�B(�6��l�����_$��
�,��4�qjl$�ƙ��v{$�ak`��"A�	q��/��-N�l�+���i�A@np�	o�^��`wsq�l#έj>�� F�<������������3����fd�BNjZ�fgY������|F�Mh�R�j�Փq�����|���_;�c7�'&N^�p������QayF��KM2�*N|,⍸ϋ���IX;�6��|^.�C:�[ڻ�����2�����g�^��w�w������qk���pC�ƃ��N�S(趏�ӑ�48�N�~��ǣ--mtuu�t�	d�GL��#1r�-�b�}c@t��$�5kO��u��:�%˺&���sL�YnZ�RG�3뵻ۼ�����8�x��[�ws���G���;*n0����+��A�ͪ���B^������,��]fY�|�<yl���*��&6�F/ �d�	��Ҋ(��RL;n�CB. �֛�ŷGF�E���M�fC�*��f�X��RX;ωhx��������8���S^ih����>_�N�{r�����dIK������HQz
���W9����bz64�ɔ�IT��ԑ�_���U���%s��T��$0s1���s�9��.n ������ԃ�Bݕ��h�����:x4ý�A-����ct��$sMG��G��$r2�X�����grB孚��j*l !!�O�s�"��b޽���ń&А���z��XK1�Ԍ����Z`Y�e�C|�wr�fͳq�������h�>'�YRA-�pKq^M]G�.�O*��ʾ�U�al���i(GeVP�~�n�~O-�YZ(?g��Y���-A��~O�n�U����f�2�p0~Y��ш���(X�v�F�E;���P91D��Xb�y��um��G_���㹤ƺ���j$�&>6��0���2�D�.j��4R�8�\w�q��Fݓ�ѾKz�d,�,�S�����t/c� �v�����o��<(f�}�����U�JIk��M����&�2����j��o)�y���g�#o���19?;�������Xܒ�5��T4+��S��+�,C��˩������;7??3�[����y���3�G&s��9g<��KP��lWe/$C�L���j�T��L2��K`҆���Z�7���F��w������py��92�">��«:Ԍs���%\��������a���FEw29aj�ԹL�7;�fǷ����?�9��3ӗBČL@�~yD�0KJ��)<�;Q�=���z���@�P���������l$C� �{�6����lzF�A)�O6������C4����ʸOBA����b1��`��Q�.徼
p}~��@�@4l���[������&#��`�#aW�U�#��������D��b���&�hj_�d4�z�7�� g��{���0�e�O6��#���cP��$̫���I�\���7��[�K�19�32�ن�boQ������}�[ZT�G/�ԇu�=�NV��Z����-�Қ�$��j��?���I�n��j|�m����`A)<���aJ�a3�q�
�S�X���W<��ϗ|��F �%j����Z)��
�w�W"�/u��뇮����k�L��'�S�u�(�?�K*r�*��3�J�;`Fh&e��s,���f��sBt�A�b�W0<yS�'�^�������(r��}�}"	(bb�9�G�p���Ux3��~28-D�@��`b:�S�I��V��͜q@.�<�z�Bɾj)�儗��Y�^8�~���S+[^���o'����k�	�@
 ���X[ o��c��=�YW㗟��<o樂����r���Ug������,kh�w���w������!S\�)��(�v�&h�hں�8ggb,�%��-���J����<�Bbj��ޭ���?��K����\�C����f
[�I���!C��~hV�V��}��|ڊ�:�o��oz��-Ջ(���Ԙ�лC���>ژK{����0k╫��\��k�"5-�~Q��+��]��[f ��_=���x&g�d*6�^�9B��i�'o�P��K��Sܟ�>8���t��a�VZ.uQ�i�����w$�e�Ǚ/����:�x��y��($�Ws7Q���`j$D8��H�?�ɮ5-��ƾ|F��L��djD9��V�\%1P؅8���B"�I��ɹ�����[�G?L����=���I�4�80׺o�� 򖒫�h���+��b-5c5F�(�_�E���A�.C:��煹u���AɤA��k'��&sH<N�Z����J���,��C�NJ�"t�;Ԙ�|�/	γWpB:�v!�?��hk<y��7ΐ_��Uӓ��sqh�ѱ�ɩ�C��}�m����i�u�@�w6�(�w�'�k�$̸o��rKp)⿢&�}I�����H�x3 ��&��(��,�>S�:��t�e̅��'����''��r�Sq�-̫�K��煆?����|9/^z�#ʿ��yb#[ b�ت�xN�d37-\Όk{��^���1gӹ,����8+�>�y<Ǿ	hp��%ZB6%�E��\� �����j���{Z �8&Z���d�$UeR��1�o.�.����M���6��NN�>��9���|�����Ԙ��� �Ff'K7����t�����'7�������{�k~Id�2� N�qR��/���g�bȜ���A��(W��Ҽq�WFד^��[��d_D��kx9f_M�����LH�c��M�j�v;�p��?����q���a>�����9��i�9��ߒ�P-2o�v�V�����V�X�](�o�w�����Dbڞ,n:vV�7���˫!�_��?�2hք?J{�	���%��fE)d8��-�������[�����+N ��La­���@x�8�e�.v����þ�:ԋ� �yRY%���d��H$;�ݜl�t��)󮆨�:��bi�{��Nc������;�'��Ѷ��o1i�""�$��[��_�:s-� h�NA���Q�Ի-�z8���,��ST
�D���(D�l�7���"��X� �<�¦�I�!��O�Ǥ����N��Q��pu4���6T(3����t�I ����(I7e>-���&؀���Yy����& ��I�2R�%�0�Q�q�7��s�ij&Ih����Ss| s���FU�F�@��qߵ�h�t����|l�ΫТ'�B܄����o���3J71ͷ���z�אg��W�c���^,p�Կc,I>�e!#e���ⴔD^D-S���w�4�)�q�������7��{��<���<b��ҍd�{B��_�\�FE�swv �^��U;.�X2�VZ��N�5ל�U�w'���b�p�e DK�v�/�@��{#�Z�l)be�1�!��0f�z�70�Y5�/rd�ɨn09�t��M��p�!Y�a�b�P�roK������B��1���Ƕ$
�m����L��%r�©s��G5����(7?p��eWT���W)�|���%���.ߚ�R����#]�Ad�Y������SQi�h�f.�(!�L諌��٫����|ݗ����t�C�;TZ�^ꖦ�'��*��0�y�%�d�86X��c]�g�G[�t����-s���=�qp�&o�0H�`����~��;�UM% D�Dݷv.͹Ωω��,R�	X}�M?�]�-���h@=��i�¬UQ��s:�U���"�?Q7��� 
+�� ��Uhm}��v�Ǡ����,:;�(��0�H��(��K8��aWK��<~^�}b�q��q�ޙt���X���2%/���潴�ơ���~�q�n�؍n�؆�F<t�/L�8:��iC���F
����GDri�R��D�G��kǽkG}[g`���a��8b,`�٧�������ϔ�����K�J}kvU��ed!K�q����_� �˾�F�v~3;�Ot�[�vK�`@��sw�U�렷��+�����'�#Nxj�AB�"�Ϙ�}&����|��5��ɽ����98#�`�������QQo��0H*
RR��tw�(Jw�t7� H# �tw7�%]C�0��3x������k�k�s�ٯ���]�,G���쭨��GS�T�;K�/KT/��b8Uj����[�/���Fu����)���3�^�{���� z�g�fgk<x��%f;{w
;-���\!=/4㙐���/D+� J�	������y�ܪ�b�`1M5�M��z��0��j���b�h�Z&��8�E͞o�R.��_�Q���<���,=_E[ʋFr��A��F������2f�zǗ�}Gn�ME������mN*g�y��4r}i`�a*P�������8�9fT���4����;)�O��gM6��{��ƠDΆ�B����-� �ޛ��A\x�5"� ��(7����<Wt�Q��z�J�g�/0Ihpz:��ΛX�k�<��8�-�MRV����0����}��
�֒R�>�v|�>�o�'ʯ��E��&x�h��*\�n^����?��>*Fm��q���}e��&]�U�h���h�֨_���+f���ɬ���ᐘ-�� ��>�����<�6�c�$Q�7s�ʁ)>&;��XP]��
S��A���Y� Kl�2���D�-_���^���u2�E��Q����;���L��B�kv��ң��-��n{��o,����� ���cR��O-g[��b$�UpШ\���RE%97Y��n�A�$^�����v�y���PU�W��^��<ݢ�Se�]�!��ϯ�R}��$=$@���y���V�0iv�����Bv��O�@3�ϧx��2v�ï3�<�Q����)�/�e_��vĿ�C5ek\;~1�=�Ի3?!L���>�z�c�ƭ�N���C�|�!^�Ȏe��������L���<)�?��AX՜���`����.����~ZrrV'F��s��}8SQ
h<�gX�1H6��d!O(1���_93����֒�������\-6�̛����`�,�L[?��G�b�X86n����p��CɆO����o�Ǯ����m��+Q�왹�C���b�U<���8��QI������:o+ݾk@Ktk��7�GƘ���nX���H�����nl!{����_sFN�?9���<&Z)��枅Bణ|�T\5xk&�f�h5{8q�I���Q��y�[f�w6�E즊�[���h���:�X�)�x璏/�@��A8�>'?��=��baDC�@����]j�i��
�(fz��x#�D�/췾�{�߸5�N|{ �5��Δt���n�C�a�/��15�R�7Z�A:�E� {�ف�������_���O�reK���6�a)�V΀'[��[
����P�cF�fi����2��3��.�V�mX�P��vڌ���Ǖ�u����sv�E˕~��	Q?.�ÑYc��3(3d����#3���t=>����pw{� e��<;�a� ��G׉mu�{��R���T�b-qjʃ�"KO�����荖ġ'��e)�v�!z�W�(�K$���yf�������i���f!��h|AQ���%�Q=]�;��
�����6���G%���ڡ�ȵ�T�T��;:��|J�},���yi�C4��H��g�r�����I��f��N�w?ʕ���E�� 1Ǳʦl,������S�%�gul#�[��ߝ����(�&�ïn��Ǡ)ʦM�n���8�O����oN��=��ohy{�"Y��Q+��C%���**5665���i�T(/��k
���qx�ִ�������I�r(��"$X�p�#ZZ��'osY�z<!��>Y>��O���~n�Bt�F\�२��m���Ub��� G��B�5�}����{�>ewX��?�n9O��LI�)��abJx��l_\��qSūȖW���H߼x�����u��e��G���Ⱦʜ�Rٶ!�X���V�6<�`��za�;�p�6�e�;�ͮ�~�Θ�m�na!RE��~:���~& <Q�'%Zsp�����EN)X�~8����"�+���SB�bl�)(�aW����R[�<#e���,-d�|��$X��=����� ���u���ۨ�,��$$�A���ɶ��s����2��d�tcr$������b����[�I�xʜB��KQ�z}7g���{ro�r��sx��rML�n�2��r$;���_�Ơ���V�iz�2Z�B�����r6O�]���A���k��M���m���}�_^-���5�x>	B[K����7� g*�v����:�ݚ�@�T��!�q��i�<;�^{�8y�I�4>2�������cy��mp�[PȺq&����6�֧I���|�Q�����k_/���#d6ex<�}n�~���=�C~|�����oj���=�.>�,A[���J�mA ��FA὆���!���3�����P�w��Ǜ��uL,�u���FM�g��R�@O2��f 6!>�\��������} ��Ge�c�b�c��^�8����뫇��������V��h�w�=a���*���$B��Щ���!����
"�$��]Ku��9�=�uY��1

ҟHc���+^��b)\b9�0|��h2[��+�<��c�uy�kBrOܽ��ѹ暰�}�8���������gm֨#��B�@�ڄl��NF3�E�D�<WY񽆃�M�á{fV�	�Mq˔X֢=��s9��gκY
_��"�^�k.�� hjڿ �N�L�/�3��Eߏ.t�{OL~�hYiٴ�Bg���NN�*�S�U�I��s������\�c�Ko_��A�^�})bD�������!�%��|�ۦr���H�D�tdB�����f^��!"[@Ck
�)i�rx��
�������A+E��/�k��u��Л���>����T�|��/,x��Ί*����>�%��/;΄Ҟ�����9&��:>�W!f9�_)U���2^v�$_���7�T�r%������\�n����l
�#\N�݄�A݋p���R�>ȹ�O2c�etͭ���I�(죥�iAg���T3�~�5y�^�gj��
RB~xʥ��nN;�t�s��c�|��u\"��;j=�{M}!�=Fpw6
��R ���ԉ�T4�}5?D��I1�|$�aV���˯ۅX����6b�D�T���%����<���֤k�*��һ��6:��*�ߕw�|�06᝕c�)��I;k���GG����fm������+�S�/p��x�=���*��������s��2���y��w�:t� 8�4u���-6y��8������`&�b΢Id0��W�v���&���9e�!N� ��r8Bjq���
�|�
n>bn߆l�;��|ҜG��1}#չ��"�R�N�����X��iTI�5��Ю#=��zY�P��hd���E���qrA�R�Ş{Z�,��B5�b�����6TެTN����U��A�9���4�t��~��)y� ��pX�h�}+C�_pJiT�W��)�����(�>��r���<��0?M���oR��S�v#��%m���1_쯦m�4���{��t?�i��>��}Ʋ8�C��g�V��J3�r5���[�g�:P@��҂�#L�{�ߖ���Q���jQC>���|;�>�a *��Aϋ�k�ю3҉��B�^қ�Q�[�I^��c�7���;����88^%U�2o� 
�8>L��R��S4����:�O�^%]��@g3x����I�����K-{�2�}�޵ČyW�_�����Ϧ���!��.���2�(�=(\i�.댡����t9��M񜐋�s��h�O���=�s*�: }r����}��r\�IJ*S�=��)�O�/'��նN�$?�6$��Ъ�ka=�j�Z���Yٳ�PKdb�5g�Ma�f�?�KɝY�+�7��'�R� ǰ{~=��|A�{�����m1ɃC����8-�������..�ǡw�/f̻�i����z��!������R����J/]
��9W<�BX�� )�����ϴ/ �{�1%�.��9���RPg�K=��o�Y�%����éu�bj��{m3�p���D�r�7�!�٫ �㶴~�sþ4/u�4�ȯ����7p�]Bͦ��~�����-3vcش�b��~����␿w��!&z ���I�C|j�ϭ~�"�2V��%����|�C8|�ߪ�%�V+�{̇����.�⛝.Y��L���r�%7�:��L_
��ܛ-X����!A3��/�q3Z8s�����lS���k�N(1� �?O��G��**�-��k�����ԍȧO����َ&�mzcd�A��Uy7��i���Ϧ��%.��� sÈ̔�GVe��Qc�lFcp�ZޅC8��=�^\�y�)R�q��}W����l����`�x{�O��A���Ū���C�'~�eA�Q3������3E�ܞY^�`6��9�8:r��C�ʗu�|-x�����,JV_�c���?�E�I�>4�P�2d�����1t��i�4��t*�����3�ir����R��ߤŔU^�m��b��x�az��~��|)=��iua�h���������GQ���=���ݺ�ӗ�G�ĺY��t���W<ٙ�46@<�v=�M���i��&��C��jE��+��a׶���L�=n�G:�K����`���D�%i�i � �ݎ�����]�m��Z%�&��?�P ݨ�<V�.3𻪍T��
�UGDO�I�3�w�8ke鿈�&��0�'��B�n>J�U��0�� \b�R���ޜXXp�����ˌ�Y�:7��__P�{'��&�^e��?%-�'
=��-s\�#�t�����T��0����M�(2s^�E���#{:p���(�.�fx���_dW	~��.=��t�xb26�� i�C)�F��Ʊ���W��L��D�n@/X]E4��M��]��]�r�="��>x�;J�xgWv��~Y��Nfs��qé���J���f��1]�����q�]���x����c���TD�F��$!J0�Oth_�U|~v����7h;l�-3��������?s����ꉤN���="%u�h�sڜ2!#J.�C����v���E���������?^.�Ru�������w�ޣ����8^iAgy=�4u���:��)�^E�����F���7��UɃ��>Ծ.#a�x��+�͖d���Z���A|<q�ا�}��4J�����ƳO�O�+2��'�*ȟ�@�S=WBټ����d5�Q�����]7V0z-�d^�-To�u1�s��)��j��Q[U����J���K?�L�&mX7����U3ݗ����^�Q{�0��>Ԛi��
<[k c�n�3 �?��Z�~U����,b���`�  �5�����i��c>���H�:�I������ �zA������-�9���8�ܤ\u3/ȃQQ(ް=f�k�g�Ph����wL���-�O���x��V��=�s�?�&A�E�D�c4����m~�.D�@-�+&v�C����@���f��BL��~�gQ��A�FW�O�%km�쟴�~1I�BHE��#kD75�k��+/�L���P�վ|넀Y��=F���<+�p���>�c�K�-�	wz��[���e��$TM��	�<!
���~����ð�J���4�4�E7Vb�}�y%��T�M.S":�A�= bߢ~�q�X�H�K�_-�@�Ь���r�!���ׇ^����E�/���D����<#��-�&�Ov�P��^Lf���-ˣ���>�A��&�sg���v���íL/v_��~��zi�gH���Stk�B�����d��Q4��ۗ���iQ3���D0��I��a�M�9Զ7FC�j�5�!c-�J�l��=s1MoT��.{��5;C�L�y==�*�c���qk���"g�zme�㢨�ǚ�=8��!�bw:n�;P����ʥD�@�}�w��ᑋ�m&�	:33.j����V:�q���&�^K�|E���S>��3�+`��szc��B]�Z��q֜�d���eMH�{�����)�a���Q~����yғ�����r��Eɹ�'7�ͮ�,c�	p�$���A��"�b���>��2�}�n����?6Q��%V���-��ȥ��7\à�?��ar����	?j�p��*�FO�ku������Eo����)x���Ý�h΍��7o��I_��Z��Q�E�t�RLzTpN����qfv渰z8I������dZ;qֹ�.y7��"�	�'Щ�,[���J-^�`2�_�G�իX�����Gq���VG��j����
��[�A����7�6����䂉=j�4��Fj�����5q�Z�	�|�����+�|�g�b��7���j��Z�?:6>��� 7����\';.��T��$�v�.���;�Kb�G?}<��$���AaD����=��gp9�� �����p�N=��gZ�����ɭ%���'.��P�qdF���7���go;��0f�3��_��hs����m33,rfWE�}I��C&ʴ�S�
 ��<��_���H���u��{���:��L�'�MtZ�����}�^{y��R�����>6�8ڐY��j��P��*.�&	1��L/�$&vGW9|C �mec4�ె���,��u�Ǝ5<h�3�c�}�| �g'��\#�}*�#s�?�bbKK>A�]�2z*�r��쿻��G��Z؉�m����j�|��D��"�?�������keƧ+f� #��\���A˧�R�]b�zh�uu���}��g�ߥto�Q��~=�lx�q]v�?��1o#w����f�R�N������[�>������5w��ιQ5��*I��0>0i�C��Q�~�n:����BA�t�NSH�����>!Y�G���e�[�O��J*+Y>����4��OE����>�9W��f0����؛*X�����	]/��U���ЩR�*�Y�1 ��c5Wze�±����u��-��ז[|�G��n�^�;Az}�D�)oR;S3z8�lAJ?.E��Η ~�ߋZ������?�r&�dO���M�d�2t���uń��svqA�#T|�u�}��p8u�π"��-a���J��WM��+�`��sX�g�X�]��bs��� %��^�lZJ��!��m�|��}�ި?�j������.�B�As7PTз�<�oZp������i����@�.�,��-�����ar*Q\����;_v%���hFBRbS�u��u:��,r����,dF�֙��\i����M�fK�xp#L=?6���n[q[A"�?io�F_CV�W��@������h	�)	,��\���n��4]��#�^��b��ܘ�~Al�B ]`o��/?��\>�e?���Ln����|WQ�ψ���_� ��.W�k��3�?�*��q���\-KH��?�R�f�Z�2���9\Zy�ji��c�RcI��D���J'n�y-v�Z^�[L�����2�qӅ>='��(���bQ��̄�����g�T�{���d�"�ϡ�tK��)���T�f؁��'�9rT�QL�M������7�j�%/�Ÿ0"���v�Q����ϸ���i)��I6吉����y��+/���=�f7��G�ms�+��~�I�
��t��(C���3g��w�i��j*�hӻ?M�����^o��K-8���{��?�lG<ɿ���x8t�S����ɻ��P{M�"vo0r5n���[���$������]�P]ئZg9�o��޾��o��w���w��wl���C®菨���dE�C����M)���0�����M*�-���f��4;��C�[�S�2U��I��q��ɚq�����9V�;Nq��Dn�:��XG7�Q��ώ�Y�q%���߿Z����Y��0`�W���b5�h�K?�� �^hDts�V��č�-H��(��pZ����f�E�<cU����t�=��j�Xk+��ۙ��Mv��<�V]�	��A�9s���iG'�3c��u��o^�{�>�ԱE��1�K�t[�{�N�C�MTi_m����%e�RK-�ۀ��gm�QpJv�ģ�?:�:����3�VZhQ|���|;#���E+�c�.UZ��ڗkX���ل'��9���=Ѣ���j��~���r�M}�ᯔ�ԫ�NX��XYֽkiD3�����}�⠧4��~�H�q���d��=1����cxsP�Q��O��f�9J���l�U"�!)b�/�y�@��T�'Xz�^2��¸�������e}��R"sOP�� p���0�1�|���n�~|��uVR��
�����7V�̂F܍� q$.�Bqۨm}2���\��������'��v�����Zm�☒sμf'}J�FOkhH�l�V�RA�.�A[W�赒'_��}}����K�&%��l�غb7��Q7Au��L����obR"$���G�޼����3�j��c��?H�}:3u�����= |����I�[Q�L����b+[0F��fA���.v��r𔁁��%����,�y��?�h7K�T�s�7���k
�V���.s�1y��X��6�$����4w���q�}��jpP�G���g���o��ju��',h69��BڀzuǜԄ@I~8��6��k?L�Gu;������~Tm�z����� (�u��³��u"_�E�toX��V��qօ��	�p���J{na�e����:��y�n&&~��΍(���y�E2G����L�O6Վ�j�U<�%�Z�y�ǜ��=h��ocdo�%o�*��dR����ZI�c�q]o>m%�"�(n��r+��'����G��_la��#Y^��9�Y���b�<*]l���`�I-�y��*�� Q�����Y�`�y�5��/m�>�3p$Z�s8$��6�^�'BϚhQ�z��c��k��'L�E�8~�Y Le���vUe��q�J�4s��i ʔ��d/(�;�a�ըRm���-��X�x�a��!���i<:[��S���L��VN��3]:>��?�o�����e3s��Q�غ6�4�RVݤEjG��tV�@~� xr�޵j2��h~_[W�c��8er&!.���2��U��V���[� �J]x$���/[�~w�.}�|*<���Z�n��t�B;�jK<��~����pU3�Ԁ�h��,�`��@捞��U>b�[��𷢕��D�%�ͨ���V�Y�7]�1O9��ku����Y�I�U�������[,)/�ٽ�����S��1�\�ۭ�B۶�g�\&��MCS�i��P���/��J�l?��uB�ś�ɠ�q������R5*N����ن�
9���⁑�}Q��k����k����a��CNĊU~1|K�]�Y|o���v�t��#;��9��RGu�Im&N�f��f�b����Ë������j�|;o_V�T�����S��w˯&2dOoN/�e8�ڻz;V��K��,��x��S	�w�G����6}��&ː�j�V�>@���	�����f���3��Dn�>��q`�Q��o��M�{��xn�mx�I�zA�/�4�+�=��J�)����q��P���,�/2~��e���w�P`ՙ5q��iz���+σFɜQ�'g�����PmX���,�213G�J�V�Pӡ��uP�*9i��ۯ���nW��+��珧�Uj1P�C-��t���y)h��J�&���J���E���
4���oy���	vU[��'�|����16�w���K�ꐨ�_O�����/�9��7�f_��T��-�=ۡ�-��g�h[*�kG5�g���Ἑ�)��81��c(K� ������|q��7�W�  �N��u����$�;��v�kߜXX(�F�j�۝R��>������́7Y'{�`[��烝�S�w��$ܟ�D�h
��m٢���/��T�V���`�(fY�z�:پ|��<]}|`*��q��.ߗ�e�41�cj�:�����6]��]dF�}:��J/:#Ir�n�~�joSP�}�e��nrͽ�����a䞁0�����<P�s�(�ЁcDI�vMѨ�gg�Ǉs��K�HrO��Z�ϗ����)���i�C'�AY�d���w����b�����x`P�PQx�9C�S,E�!�%���k���7O��ށup��q�A��̼��[C<u���t.#��<i���]!��;Ī�<W�<*Z�WM�������(��k=�C<���؜����q�;��g���䖉��a8��0��5!��U ����Q$^_��#���θ�ضk�hWK}h�@F8-���n�[�:U��u�:�'�!�(��=�/�GEpӅ��[W��k�oH2>R��NH�K�f��^�Q��+]�����4��Ex�Ŝ�FU�"�!S9� OǾݼ��˒�X'PL��h�ә=��}�I���J��}IV���E�+1�K����e�������W��:k��m��}�C�A�ڃ�h�ͼDD�����\�BXB��W_:�=3�;r��pV�4I���,��N�!^�f��L	_V�o���T�<��2�w$���D�zhZ�j7۪�ZɎ����/5���#�.�<{?hG���5U#FĹm}�A��8���1:���%��F����\��������Df�+0��	ۯ��
(*k��Az��+��ɾO�{��A�J������rm�����=��l���@qFy5^@�����2���Q4�G����OBV�6��1����.���f�ޏ�p����P<.py�'�!XT;]2g�ydܾfbR;w����ی�1��a����2�&��<��<)^]�x��#�A�%���e�{��Z�.��*{��(Ĭ1�ݩ� ��	x'�9�HS�i��.Ȩ�m��t<����5������5�,�����������U�G��Y�ߢEYW�k���o1�Q���c#ѺO�4"3D�CA�C��{Ϋ���cs��8�,��+�^~q>3_�lu��>�ti2ZbKF��Ny��T˗*������: �W4S��|��τ9���4��l%�u��/�k>	�ޅ9��*((TQ7�pq�)���]n<�P�PM��&I|���C�d#G7���DN���BIPЀ��V��N?ٚ-�w��l���!T�	�{',�{3����2��
]��V[�/N�އty�-�A�bѸ6u!tJz��GM.�PLibx�z(�����yL v������|@f���m��&���7{@xw}�aYȈ"ȉ�i!��"�R��F�k6�4l
�%W�d[�
����cP6	����v:�MW�.3e�P��)xq�q�cRrt�{�-�tm-j��Ւ:C���V_��σ/�G�%��D 3���vt�
�n΁��/:?����Hy����:Z�ǹ�E
���Pm��l�-�Ow+�ATRK�D�MB�r�>Z\+�϶��`�)zsC> h��nıyH��ep�ݾ7��go#���������L�ؑc��ҧ�l�@
��ړxX?�vֶ�H��~�0�%9o���.ik���a�Tӭ�GW��1 M�}�%�QJ»^~�ϭ,�*�ww�Vc^����̸>�ό�X�d�t�M��h�wP�CY0�Xj�9kC޲��	�(�PG{& $!͆�t(�ᗚ�]��bF��ug2s�!��A|OM�$�<�K_v���=�x�]]�@e���'E��#tj�dÄ�(��."����`����Q��)������h�J��ͳW��w� �+!���ڌF|�$���K,PZ�l�y���`��d�zۆ�u��5~��|�M�������L�Ł��b�Y�r9�t���,c�Q���y����������hM��[�r)Ϙ/�	�|�-�e  t�a �Ybx:]IQ�`��GL�VWUwαS��s�ï�^bO9J?��2��m�-a�=��t��:Z�[a���wF$�[�K�y)/�:Bg�6n+���V�ޛݔ��;�1��d��(f��"����uk��n8�;y���@>�]�w�����8���}@�kH��68W�ڟ4����ͫ�q�w��#{��(��}�������M~Pߵ-�i)��}��x��������0�X�n���1&�\��m��*m(9��B�3��S2��(B��>L+��p�)�B��O�Y��m/���Aw=�	.��j�B�?f?�n��EV�{�k���N�^lx�Iq%vF��G0��J�ĺl%@P0�1�cԏ�d~�S��F$a�ij
T�5�cj��z-\=�� q�y�8-�+m�cLk�]�}�j��sf��D9��+�#������4����yX���㳧u@7v#�b;:@�>�����[�!7+s�X�+z<�jX=Ȍ�H������0�C_�:�M&�?����1�-'#��ǲS���N/I����F#ZJ�U�8�:?��&��y�R�����S�e-�������j�$��]��UW��ҡ�O��bZd2c&^�J�0B5�o�| ��b�S��f{g���h�3��	`汍��2�}捚�Yq�����3q7�R��u�ڍ7�` �������.'M���.��C��k��Q#e�},��a|�XX�S9H��:E�r��0碉�ĵ�_�㰣��%�������|�7ʯFs݊�0�Qz�6�nk$3�ü��w-�>bT<�>��4C����]zZ�ۧ�dT�$h�����ȗj�\�TD�0��w��>4�\�d��<�2�L��k]@���I�ŀ9k55�h�X��2��{�z�)��ԃ-������b�2'e�`*X���56�:,f�+�Nn���'���6F�M�9���^X�~�㛤MuS�P�ml���c�LM>�k�5 ��G�w�Ʌ�#H�C"��[y��S�7�G�5R=�J��d�::1���MtТ����RT�g��`�y+~���A��탣��J7��a߆5���}\{��&��"W��c�v��άO�=�>�����^y�0�.Sf@)U;�C�W�ۼ��U�ˮ�Ȗ�8��D�/ze�S��
��[�����.79�5��dJ�>���$>g[�
۸�"�i�^﯇=/�'��ù�/ݼ��%.�9��ʭ "�0��B���;�U��Ŵ��~�� ���mM���4gJ��s٩[iIK���Va���+u%"��/����X[,l`�2û�'N��X�W�l�f|QU�x����]���U��_ox+l�Bk�o�|��ؘ���X�� ����DMzvi:Qy��Cl�#Ӌ��:��݇��e"L�W޺�c�tP��mW<�	2�Piɤ�5���
%�p��޸l?ýC�8�T�9jbQ$�-���L��)Ж�����i�j�M�0��KĤ��<?�z��C)iYY�x�w�ثȶ:�̱���j$�jn@D��Q�% ��G�!�tu2�����qa��/�t�چ��+��-^Ξ�~�y�������"��!\<�!N
�R7��*�f�����(XN[���?��6���9�
Pt�'r��+
�0&�*������fc�DV.KU1����p��(rb�H��g4��~�՚�1qr+�UDk~I��W<6q�==�Ƙ'�w��N���HE��S�+�G���F<_P���.� �}�~e�׉Q-6i_�K�h����?�BZ=bب�D�%������H
HϔIx3|/*�������禆�_��n߇��jX������,gŨtQy���!������3��"n|� ��5W�,�[�X�B�ua�ɞ�+����4�� �t��B��h?!�n��J�Fş����4���ѹ�XA�v�C��5#F�Y���U"��n��~�\��l�L/UB�%U1�-�|X�L�\��}��WQzTI������,+�/[]V������*��L�'A��_v᤹\D��yE?�7�6ͱ}v�5��eN�M3P�-y�*���/��x��d,x�<�2���y�c���^Fd\l�I�~Q���5�D(�C�[j��n�J^a���������#�/r� �������=��E��9^��(�If�ӕf���Ȭ�Ui�Z&O��YS�y*3�tp�U�h��M>��u�kN�����3�Kg�3/�\>F�J�i{o������t�x:�I]���6Az���ht���mҏ����ќ��iV<缺��e���9J`]�٢b���|y-�$��zk(u`�cW-�̥w	�I�im���ʷ� �w��ٹ�Ɖ�׮���+W�j[( �=����Uk�T-�x.�[="���kD')���fX�Ie�2^pWU�$	�n��#�Z�3D�a���~�P�0_�$ �fml�|��躗��O}�f�T��A����>�B�*����5�S��E�a�6F$h�'-~?0����������op/��M�_�=���3#W��h�kiC����4^]���.��ީ�\:�Z���I�F��S:��`4�ii����t}ڦ���J�BXm���rW�&��\L�R�=޵�`�,.l]����rwO	|��[�N ���mm{���M.-g0wh��6�u�W��9���BĈט�>����'��©���u#�ENr��x��D_мk
��w�s����Eu�҆����j�O��u�w'���T�����#]���9�F��K�0�fW�J��,~z���U3]�X�h���R]w'9c�~=�PV��a�U4M�it��;A��D�����a�&��:9�MY1RK��72�����w`O�-��S���6�jW$��[)��k=b��նl�	�S^����K�p��������
h��5��>k�5y��J�������@�oPå,��^s�U"�-vS��[ȥ����tn����J�-S��͟|h���:Z�zI9�?FBGyӲo�� a�ԟ(4~�;�����������T���q�L|D����v�������Y"}���;�Y>�l�?;�+tH�i�'y�{3�����i;&��ǎ�4ƞ	)�
�75���0��٫�����Aץ�>���8~>"X0u�b���y�@�kEK��ț1�o���$���a�w��*�SmH�{�aR�}a�x����N���J�3�����x��c����#�`��L�mbvк^�{qʁ���0_Nm�����v�����qz��n���+��a�_{�Ոh�6�ș{׸��n�+�*�ɚ=���( H�?�ٽ��x֖D�& P鳝����@�8����h�R�eX��F^���!]�6�o^׏���QN�� d$z�������Fs#새�[��/P(��Ur۠�r��Լ�-n`;�nT����5�l:Z��-$�r9���!��qd���m�-	�ċ�~�ې�h^��n��,��V�.e��u~S����{�?y,s�ǘ^�ҏ�{/_V�W����;h�	"4�*Q׭3�o��r�iX��*G�,;$T�깥�Ǌԩ�V2���M�:`h��S�M>
M�>˷�;�(��t3H�z�A�/X"��m�E��!g����D�g�z����˚�#v��M�J�V%iڐ��vo��Y~�z,xS�9�nq����������\��{����������X_i�u��)�{�Ķ`A������~Ƌ�t�34q?Uru3��������އxc�������ll!���m-gJ�)x��k4O�7I�ޘ-�ښ��t"G-H>�s�[�֨��h��l�jM���ٵ t�����{�+��������I:U��((xT�-\(Ɏ1ł�b 6���Q��Qm���)1V������F�g%�w =��1_y5��"7�K#kgvR��<��]*v t/edP�$�w�f�o4u�|O6a�bg`�K��=o��Kr-�n	�o��'��£��ڞ��8a���^MY�����	@�v���ť򱓇��Ӑ�Gzd�̲��:o��m/�KP���ָ�l��ة˫Ku{ו"2�{�Y�v��L-��Ĺ85v]4�^[�xe=���S��HOm��%fP��5C�ʚ�m�����g���K�/N�
�C��a�t��o�i��E�K?�M�c�:c����k'������U�.����˂�Q.�؉Tۓ�kc��Cը�[�`�w���D�<�9
܀�Wq�u�81F�Vv��EGv���\��i��#������Fo�c���yĮ�^ �~�o�<͉]z�/��cE���t�(������o瓹�o�.S�'Ma>mML~������y�5v�.N�a����]�UM}_��đ|�_|i/��1��u	��-B;Aq�E��B-nA=l�{E~�~��|�#i.��<#�4�����U�C��`蚙@K7�ܪ���i��V-~�0מΨ�R��-QI��%���ΥPtf��{{oj���$��e��� a4����8MSM�|$�ɾ��~�Vw��8�����c����p��0�42�/1g����n���j�3MGD毺�+m��柭��xl\m��g�#���*s���n�zZ��e��̕��ޯep���GRڒ���5>L�˸�[��ߗ(��U����x�p4��[B�(L}@�}r�|C��[w ��]�˶[O�ƽS���:Q��m����/~�k2��sp�����x�{�7�;�es{M��j�:�sw�/��T�P+����1韜��O=E�c)��m£Y� Je1ZX��@�m6����Nk������^s��I)d?q����*�N���.��gҪ��O݃/���CBU_ yF�����{�?��e�.$h�YӰ�}����km�y�W�	��9��i�Y�S��<{�3B��^Ǝ�Ӳ�g_�����"|�_V���͵E��v*�^?�Oև�8D�Z�T��]!f�2�Ke���?3L�@F	��սr}����\ؤ �e1/ �[oW�u�!�4���Bp���A���,����K�{������������t�[���}���8˴F�E~/+k����J@�r�i�,H�Ϻj�i#��[�D`�װY��nCP�"X��z�?ލ�铖y;�������(Ƭ�;2�Q�8�+�I��;ln�M�����W]:�-&��M�� ��m�y�vT�Eϒ͠�|�<�:F1e�%��ѐw�~�:���^�^�[��;{�l>;���ԉ9�[�m��|��^տ�#����Y������0"S�R�C�����>R��-�&����mm��ޜj�{��Rl�vQ�h�j/=Qo����Q�$��숺�մ���b�,���"��O�Ά=nL�3���������x��g�7�$��O%Y!sqˎf�2�E�#9񜈚m�=R��_C3�a���H��*���v(ݫ��ݡ�
�q$}~Q���l��� ��
�&[�����ѻͯ�f|FYQ`.o"O���`}1m��#55���������'r,L�x�|^V2���N��$����xg��ʑoGv�[)�[?r1B7[��e�z՟�V<]1ؖ���	��c]Yi�"qt��I����l�B���i������:��T���ڸ�@��&�yt5R=+�;#D^N�v�f�׻L�L%n���l�ѯ�^����K�}S/_�[k�M�(8�GJ����)b9�3,�� ���͇Bx��[݅^�� z��ү	F���gđ��� �M˭�����&���"���a�pT�A��rå�zb��Y��^8�1�d��G�g�_�%e:���K�#�IYB@o�j�U��"{��%}�|�P!�7;uA7����~�7	3��=ڜ��&��G٪-"�����b��ί`�x	���:���q7���Fg��>`�h<W�&��� �r��J8�=$_������&���B��՜��:mt��!/?�(�ψ��?��J��n�w��"-�	rg�~IӥPg��j�(j����z�lQ 9�.���8%*k�i6�����ɯ���m@����b@��(_��$J�h�8'������.��ņ`��ˡ?h�[�b�u�?����K��TƵ�88���x-�}vJ0�(�9�D��]�_�<�1l�m��6@��k��*p���ld#c	�{�l�Sѐ�`Z������2�l���%н��;[�b\��r��+��Ml
U�C��n����i(Z=|3�YM(���-نE�CM�Ok����߅�z��G��m�C;,cE��&)q���i�"��*N���Z5m��@+6�єO�*�ޖH��L�v� @��W�l���</�֭��i�o�ϥb��iQ���%�gß!�N�#K�ݭhgS�)*� �?n^�8܊��y]���:��w���(��^H�(��	��Z/q�$!s�F�l��n���b�~����;����Sq�ʊ�p��'ea�+��D�)�]���������̴����(E�Blx�g�h�/>��AH��Z�����,��:�QP��Wi���^�����'�� ����O�k����R�v�������~F�'��=E�_�O�/F���k#Ͳj�]����Y�4�z؇��]��Ć� ���S���s�t�X����T�ߏ}=�蘙�;Bqn���o3�<䴕���T)�mۈu��mc�>riz5Cϗk�_��:c��AH��S��0�&/�p��o0V�;�y}}��q��1h��C����m�)����������T�W��l&�K�m�~��_ۥ��:6�_9����#2�bN	�U�j�B�vXOweݭ��.y�0�6�|KgeJwٍ=]�}	�������+�_Yb������C��m_aX�P79ܟ[�2d�3$k��>},gKм2�#g�=�j)g5[e��R_=�B��� ��}�%��z�`N�V�+�[r왃�ǷqW�%.F�w'?��I��U���?Xp�<�,�J{���PZQV_�=>��O�;o��qy8�����Po�P��cW;ԙ<���J�V>3^9��AZ�(����P��f�+�*S��%�.]"�6���WT9�ᑀ+b�k'O�k9Prj�G&L�4|@�D�D=�X������4���A �.�!<�O���Z��$�l3��A��(� ��Jr|�s�3�D�Ĳ&��[��t�wg��W!F�Fp@bj��������~�<�%�'��O���� xN��b�,���s	hd��yo��e�mCD�'�h8���rE$�/�RУL������2�]���2^�ڿM�� �����v�?�o �q��w��(X�EG+]�ב�
����"�g�}!F=�xd�<����]�!�JqM�����ۗ�]LČ��/	�q�5��R[Nf�:bd�e�J�k_
e�ɞ=�~����ڦ*ߺ��VF��:��}��/���+r�F�.Q &�����9�K�=H�}��rF�\W$����Z��F��
tV�^�;���o���'xK�."l�]_ ����
(Iߞ�\�4�����j�Ez�;;=�;K�����S�0V��]��Ik+J� G&Uk�ߋ{{c�}m��;+�gc^�q#�%��0����=����織,���]�t�i���m���BN-�����Wdg�"��g�?��	��\�B<R$�jKgdPMf	�8Z��2���2���xG�w;>�<�-騷�i1z��ໂ�0��;�N
��̲T�l:t�Uz���@�U����Hn������$xl�Zz&�L|ן���걛�K��H�[����|���o���u���|{fY�wv��ت��p��{O���N�J�b	��M,X_������y���_��<���ŀ�)N����f���_3�;�����$��>�u�8xxʭm^D�g��5������x�T
�~��\���'�^��x��������#B����jqD�c�٤kՐ���������,���_4���y��QVlA�y�gD]R>�,ȿ}��w��Qi��� ����� V<����}�K؜Ax����6|�=��Y���߃ES�S����35��i��}:��Ӏ�Ā辟bI��[5,�6���l~�tM4�r�U��� A@����CL����b�wA{z��i�k]��u#e�OL�sWg�\�h0�>�xn���!8���&:
�x����ϔ�7�m�r�7����=m큂�|r��cΕ���������x��U���rR�x>t��v�<��L�y�����r��(����(ܒ���XB�J�jq�z]��,R�|J�T�6iAC�������=l���6�V��=!�:�>5���v��P�r�+yb����^���n���F��V�A���n�5.G�����p���������x��	����
��|��qL�_���Mi�8g�f%�&^t��{q��GBN���q��9#�8��z�K&f+��?��cQ�֫�<q��_�ϿK���u�9���.,�w�m̗��T�P�Utӆ�܆�����60@�x@e�����X�_�������A��'v��|�d�k�ܼ?�=d�p��x��ʮ�nL/�9���"�֎��P ��ٺ�l`��Y�����~�p^�F��n�����l�5����;�>c�K99��d����AС�ī2�eC��}L-��	��8�}��*pg1f����#��·g/ߟ�^��[�r��<�^M�?��a��F�e�?*m�Z|�j3Oq�l�b� �W�2���^vH�_��b#��MxZ�Ѻ؊5$��;�r�,�T�w�50m/��[�i
�>\� G�\�
�o�K	�H�Z�֒|�
����-��,:P��U\xo�uk#��C	�oAe��a�(�a"Wa⣅�g&�l�g���܋������n��S�N��~�=�J^���$�^�mK�⡙<	�Qs�j}�\�J�@U��x+�� �E$ANE��Lx��=N����Q��x�f}q㠹����#���gf����z`�9���{��{�0�?��w*�~9[4�~[dt�����B��7�EaĬ��@b����:� �5���N� C�%���/}��V�M2���el�H�!n{�n�8��Y�$�H�~��7N��g�ح]��.��� �{`�d60<1۠?d���xv�}��HE�=k���o�� �cX���m�n���).������Q���t\�>��K�����g�|�{s��B���0���s�v�]wrO._o��.G~���&ƺtV�F��N`���d	��o�{*�e�[V��#7��a�q�~��j� �"����}��A�{����ˈ��+n≅��R� �N�]����A������u�͋TF`W6ؼ��4�����)�ʌ�y�N�CR���,�q��P�^����i��g�J�E�[�65M�,X�vfs%��� '�S��� ~�%�X����q��L+�߮��ǿi���T�䅑h�P ݃o}�ؾ?t���������^������tz=��TP����T������%ר��i���a�/���nbF���������9�0� �LQ_���o��"���"��WE秲�۞����yjl.������I�_s]q ���hQt�D*�AQ�f�PJ�D�b���g0X���͈��|�^ʻ�u��{�v�7�ѻ�ޓ���E~��j���/6Dro�tٸ4]��9����a�z�G��Ita�g:2j��?|m�Ƴ�-(�G�k��c��йrg��3��Kȓ�AZ���]�c}}��O�\��E�]��>�T�'FJ�Ai�A������GH�&s���+�j.G g.��a�����1���o߄h����j,��;
"����.rJLЀ0Ż��jיjl�=2oߙ��JCX�xM�`3��e����p�r�մ��i����'���&�]8�jV:��6ծ|�[��܊Hc��,7z@'��m;O{YE�"R�[� ��+��]�Tit�BM@O�!6ߺ![����kA7;%;���GMRA��Ko�d�f=�N$s�W��ǭ����+WA#	��`�fCk����ㇳ�`z�8܎��\���ux�1zĴM�D!�ߡ��c��?Y"�,�d�W��%w�ugu�*sd>����F��4���
N���B8�"G���e�#�f(�U�*�&����F�������-]�d��M�x��2�Qo�r_x��Ɂt�p�?�2��,��(0�u��q8���#QT�O#�Ж������U)�y1J䶲���xvF4�棠 *�@
���pa{�}mm�^��d
�.�.�z*q��D�;8=�Ȅ��*�J�;�8�5Q�>��*�1� ��埻Ǩ��c�_k����L5��hbE�B�����3.i��b��h�7!�u�	�&W8"{502x�؊��t6��U�/P���'63=1K���4��B�l��#���vI�kY�4����հ]|0H�}V�u^籇��x))?%-t����6���\�IJ��Ls��P�`�h?��C0��n�`9�Ȑz��y�P��!�S�	�@t��<6 �VH�?�nJ��i^��ҢX%]��r�p'XBvz�㔍�f/|덬p���M�!�ϰJ"32���� �g��(�_Z��]�4�7�?:.��V�AS �y�����Y����8U� t���<��@PX�Zo
V�����p��I����g)��,
;(�M���l��<舺n�ٜ�[Z�4m�垕����SQ���\#͈�����M���V���O���ZkŃ-��T{�cs/7�1W#�{�v���>�ڏ�Qj%�O|>ѿ.�6a�=x?�`N�Dv���c�c" I������&e�J��_���5�12�����H%��a�� ��z��QDT�B�a�J�=�(���������ZXp���'ڀ�`vRo~	�_%y �Ud�n\�4>5R�&X$C�n��Q��Јǫ�PG����9��Z��U8-ȑ����K�t�񋋷p�aL������6�*��ƽo߾e,�<�~� "��y��J9_�����%�uۧ�$�3u�<l�ε�P���Ye9��;h�7 A̙�
�h�oc��������A����,nc�`�!�(��T{ش�����/��cF[<P���3���Ʈq⚂�K>~V�JOC�:R�ƪ��PDb1I �;?[=���*����
~�o�E S�Y������l2���z���/ݾ�^Ͽ'�r4�~6X��v-��o��}z�����ü��p=K�� �	��tk�1ɼ�x� `��W�}"17_O�����L>�GH����%�p~xT�q)��\!ۧӛv��V^�W��ɉ{�Χ��o���V�h�%9H��ѝ��!�)il^�}������yd9����n��Z�o`����V�j�˿J�C�M���Ǥi6�"Q	��'��0h�	]�>O����H�&q&J/��j���*��i޾zI'�� ��w����"��}�[E�V]���7Uk�T;���-2��e㴏�r�űr�����fa���t�D�v7�F�tt�4�D����쐙Z+�s��U�[���[̳~�|��D�(!t���CJ���5���x���L��+
�Y�nE�	���au�$�fHH4��_%�d�UO.^���lls+���Aꎯ^��.��~R����<�iԮx�P�IZ���Q�R���oa܍m��������K�b�k�D�LmrPμ�T��>��a9�g8 \@�s�K��ٙ�x�U_�i5�#�|}	�HRa_���øv�sFC� ���1[���W�}��=�rΉ�*��� �dl��X�`z1Dc�>���Q��a*lia�P��W9�|��5^�n��+�ON�:����MJ��*���X�*�"�w�m�'[�;`�֫�8q,�c����&�f���;N�j��<l�4�w|1�oz����/�}xd���hA��$W�\�F#��}t?�.�Y��b���b���&[�t%�8p��u�]����w4Z���)���l6� D�,ծ�VP'��'?h����X���b:qɩ�A�D���F̼ؗ���DD
��q9����&U���K�i��vӋ6��� �����=���������3щx9���Z�w;�Ѓ<��=���nY������uĔ���>_��sq��c���S�����j��Ϲ|O�^jl����'�&9�o����fe�H���d��ʠ���q�D��L��n��"N�����6��DQ_ȌL7�N]��g���k�r���+@���{��殳�b���~���������^��엌\�Qo�"�Y.�#M�L�$�?[{^,г��kM�q3���t#��k��C�ӿ5~BO�A��4�!����9�d+��z���V���e;%�����6�S��V�]VbbtΖ^��΍�������[��o5� �6�=�G�^Ҫs��k�e~{��[�X��h~��r�g��:	ۍwۍ��o��;F��Ң(%���sk�{����g���K�05Q�w�b�8|��t�����-5�c�S���{��?\��
��;�P��;�L,�N������>O8����Iuc�^{RL������������Q};���,�ͻl�!N�ܰ�׃��#|ʧ�ӝnt�O�tX�,>��a�K�&D�Fn*
KKCΔ����!��z���d�,D�	�L�`���6��Xk��;2Bl2-/]���"k��lr���VjV��ږ?�º��4IZ�'d�L���β������{�eJK��]�l�ů���s �I-n��������Z���]���"
�d�(���Lj,����b�A�Iɠ��!��u�'	�L�����#.�����������!�6��Zd��m�w��|�ٽ|j�7��UY�4�m0"�򃃽>�bd��]��n�ڷt����23(1`ⷎ� ����^%�e�p}Pݷ<��Cσ���
N�j �_wyu���;�b���<F:��8��2�����牓D��	O�^�����nx�s��˥��Ey��.N��6���o�a!FI�e���q�1HH���*���3/�{���,�ˌ��Ѳ�q�\|�T�5z���ɘx#�i�l΀�Go��/��E�[�*���E�-1��-�tE˿�9I�e?v����t�jT���/#mҨT�R�a�����[�+
�հT�>������bQGEC6�n���PGn^�I����7E�.�S��k�],��{�����nV"�O�W�@ YM���∡6Ĳ	jdes�Yo���8��ȨC�cE=|G�l��ixe]y�7ˆ5������*���B .\Ʉ�����9����RwX2%0	'n���G�?��K���y��Z�$�1�s�/޳�
#觔a7�8�D��!�P�/ѵ����aI"!k7�18�x��~> ���j����`�P�����%u�N����`n�O��?vC9v��Lŵ���9�4�^D:��l圼�pj���q)W�l��D�2jmfE1T��ۋ�@��Ţ?� y��wL�_��_�����b�,��G�c��[/^�苤�GM;ejf������@�s�[�L �����h^x�?�T��`v��q5`��f�&����r��:Xp��e΄�n�?-�Z��]�5\����b,[�Ej���ױ�FI헪_1��ɮ�mlm%�/DtmA:γ�NN��݇����G���-\~kC����+P��~	�����R��4 �כ{%�<�_�����__��ԔD8@��i<�2��������������^���'��GKAl�U��m�Vy`:F�n{�B�]ts8~:�[��P�^�����1<�jJ�rҜ.c��,�)Hi� |O �6���ݥ��qNZ��z�
�������N>�c8�g�?[�5jSl~j��I*�������s\nk������س�#��)����'�����E�5���'��Y�0���4YYcG������c,
�}�d[�񡟔����J�~ۡ�w��Ң;"����D=��A����xU�q�ř�o5әW��E�:�@٬Z��\p�R!\�����%H&�v��.#Fs�J�:M0Z�ެ���.�����G)�dU�b��AD2�:f��9m��4��o����T�!H=4�6sm� A���e�eQ�I�sd�y�F��"sa�ދV�\t�A��\MY$ʓ��a��(?k)��m���Ф��7����~�)�ߔ,����z$��[��L�Z*�>�ǖ+�ǣi�&����$**�8\�O�$uۆ�rg5|P�ٙb��avF*��V�𾷤����[��P������`�Ы�$����&�s��b��S�����Mxg�1*>�KB�y}.�ȉ.���e:n�hy���&�/�\�(&v}��B�j係��L��Y��wɖ����w�f��o-�
��݋��xlұ�iU��Br��9|����P��[���&��ϵ%{�a��1���5��9�_�,�n;�jA��LOr�O�d�x�y����w�fҵ��V/P�>�xתJ�m}©(�?���Õ�҆�{`N���z��_/�B����Q�r{�K¿K+r`|v1�xv<zi���0�Tv��)d������a���Ǻ�NZ<���c4S��b��'♌2������;s�$�OM�ǖ1=kv
���g[9���q�RR�
CϗM|�v0��K��i%]�^�]���(�nf�B���A�q�K�L[]8��3Q����l �cы&�_�J�}ٟ;��\Q��@f�OZ����ĵ�U�ƇE���ʎ�t��f��j�:݄�v,z0��(8Q���l��{<�(;��3��7��ٍ/!�|����Ds��S��S������Z������C�j0m�r�f�a���h�d5RP� bv)`�|����U8wlV����nˌaK�Z��J<�K�\���W�jx�p���t������3��X��d7�y��gDS�G'�Ⱦ�m��7;;.�q߳�[���X�)z7�������`��r�"9�C����%	^�ꤞ�t'0�q�4坾���9n��i�Ւ�}h�#퓉'ݜZv����R���Y��-��4�z{%Y�g=���C�¥�"�͓�U�
M��/����GH� ;MH�:b�y�[�rH�к?�#O��A�	xgJ�NǙ61S����a��4ei��I�>�?J\��w�
�3�f,�V��W1���@���,%����t0����'���{�O�U��!��-�9A���}Q�p���U��P�Ѓ^K��bR���z=@!��1��@�	���i_�h��$��Ԣ����pɪ~�@�����f!�:N�@J7�N��������- ���i����O��.|5��@6́�o5��A��P�7dIW�E�^(�jқWe�'�ņ2�R�-g'q9�ECGǺ��,�8IL��t����g��{�ˏ��VS���h����=+�m�׸��,���i-(䀦{��򧒭����v�;C�er���[Â��2�����ى�O+�U�^{}"�!3?lII�b%*[Y7s���#����<_C6?K������`&+��g�;�����Q��ok<Xl�Pl�0y3�\[����J"���Ն)���݅ub�	k�+�袲�������X'����`J�u���)���P !��Qt=�]Q(���EzA�E#)	���@C���;|�_T\4z�,��Ƕ�0��!���A4�l�0����q�6�M+~*����"���П{>��Fo�Ϝ^�lw݁�n�ġ����{�ܨv�&W��r�l��vj܁�����sG�4:,��R��Z6
��o��`�� Q�$�Qċ�l��A�u�4!^�/7Ӏ��5�&}�I	t�G�>�k��&��{2[���g��%�y���,{b����b����mF�I9���,��Ұ�-��hf�D�\���b�����ƹ��5��gq���t�w_���`�o���z4	�
��jЙc��W��^	��
Ac진�[�֏�CD70����_�-wA�7����W<����g2Ю�Rff��{����4H�DE��>gK�[ނ&si��1��X8��~]k{�hh8��n/��`��,��{�[	�^p"��~� �ށ�v�VC���"�u�{���G�;�m�t}D׌s,Ow*˽K���L)�|�G�_K�	��i\����r��ޣ��|�~���N���ǩ���K�5�f�p����qh�,��e��gv>��m��8�'GGGW5�� 9��\�7��7�dj��L;)oOݻ~�Qh ��������y~.o:�N0����r���z�/��hi��3lT�V@��}����(����8�U�u�����Ӗ�ֿ>y�@ڤ:���,��yWD�@��Vx���/�R����{�L�a��i�n�>��,� �@����*X���eT �ɨ��l���5$����0��8�e�<D>�/���4^f}��a���^3UD�ǐ����	��Y5W�];�E�Qz���HWEg������V�;����C��'|�[QB���� �e���f�_*l�:}|��>`�8a��w�
��a3�
��Y��0�C�<���W����0�;: Wu�d�Ŕ`�$��SLÑ ����C{��$�IG&�M�̂�
��������4J^��&*:�FB'RRMG1 l\���5Ϝ���R�n�����K����5��ӍYM����z����k��c�lѿ�����7E�� �egc�������2"Cq�7l��D�8�B�uW�i�|)���[
=��J}h�����Vsy���J��khzz�{�|^O��ʊ�atola�Ic�����K��-���\��o�!XE��8��<Bc�_�(!�<ԋa�����������P�Ƥ��Ԅj�p�]|x�|���{�:1SE���TK[�������f����~�����?�UJ�0�hGݚt�����N�a]�Ng���UY��`����?�3��50�0�P�.O��8LCX����%ټ���Zy����� �4J�_�h����#��[�H{5��������Y�>��k��Bk����%�^�,���2ؽ���m���2E��B���UGR:B$~^ �� Z�^�ȑO�V�k̯ǡ���r�%�<Z����p\l?�Tl)�<����.��� *��!�;��U�I��lo!-Ymq���YjR}he�����l+v�@a���o�5��,��.�Xg��M�ܵ��^���I~��[ _4�y���o�f�׈ȐH>e4�*����/�Ҝ������^K�h��{�>䏛⤊�*I�UP�σ�-���,�.z�6���3fh��ڠO�ަH�4;��y�9R�Z�����C��t��iQb(gf!(�1-��4��s�G�N`�� >���_���)���7ǹ���9M�o�����U(�P�wA��V�[��PP�F��Y�L!�5��Ld̖c����!��7�=�f��a:^�}O�����T"���%���h�'�����G�s���M��(,I,���I���@op_N���c��-)��8���\�36^�%���w�a��ш��v@���kK��7��2GЫ�4p��\n���򭭧�ON�D&P�K<�d�(�+DL|P%e"å5����LnE~���Vs�ģHH[� }"��3_�n��?y�E���f�֝�oܕT�.TsX��e@��2s�3���wZ>��s���-�f���U�&C�
_ΞT����Hc������{)&�:cH���:esq�ۥ2F�<��"�>Xa�;�hQ�P�8P�4�1���'�W�Z�*�g�xE��M�w|��c��g����0s�\<� 1�?D�Lcs�D�x��9���S��.�<Ċ�g!���Y~�G�|/�uX��8ؑ�����kF0{��祪o��u���.�J-*M�v�MM�p�S��R�no��&�Ԓ��S�!9Ck��y�-M���bH�Fr�ڝ�P�a�׶U5a�z��q��0�.a�w`���ܻ����A���І�d+p�M��`���o�C5�k��	��)�6�XѠ��8�L��]��Tv�o(|z1�z��p���9⍆5�*A"ey��O, ��Q�?4�0�oh2L����&e��u��'������R��G+���J_A�Fצ�E��.��󦾓a��F)�|��`r�%�����6`���]}3�^��f6;N(1�ְ2ZE`*�pA����6~�R��pϘ��|}�h� ���d�Y}����F��֋��*B��+Blfz4�a-ي
r�^%�{sM���^J��F�a�U�����[҄��̀�yإP���Uآ�jj��pn��@2��9����q!��o�l<�;n?u�̏Wc�j@�
Qw�;�#:�j����r�_����/��������rW�A�,X���gC�R ��1�����UeU;�}үa�>>4����q�6Ta��� I����W7����8�V^(�(v�=�WIup���$�Y�3�b"�N@t���}���u�ͨŜ*�#p	y�"s�-m<|���yy2,�'�M<�L��,�F.÷l<j\®6,i9]#s)Օ(��(�.$�P��� ��l\�ƥ>�����w���"�xH)�MWp�c�-��^����M���C��77�h�
*,x�Lz�(�N��dG7G�/h@��GXW�?��,�o$�b���I0V�T@��[043�f���w3��_)l:��g�_iU�
ϫ�U�w���X�	r�@X��RqC㫔l2�|����k$㽺����dl��Cc�i�~�p���jN�*N��Ď_����k8�s�������@a�L�L�.�7��鑘Gi(>��N�gE�0lu�x-�.:�G�ò!,
��Ñ�Ru2��fl�n�qS		]�kq�s���)�Gs��(�Ix�d�B׺������ w���������t�=�Tܸ�f����ݑ�C�\$v'U�Z�OԕQy	A���B|0�9G�9�͒XN6���/��;���?�8x֟u��r-;p�dd`[?
{"W�F:M�jz��a�l �M�(A����b�݋"0��q��`���
�-~�Y⡣�1�/������zXz:T<ؓ�S����;^:�߱�v^+��eLg���H�P��5ֲ�4���=�ki��?�z����9j�·���nA�<=i��
�Z�(���7>7K{�H�sM��EQ,ݪ3��ЭtW-z���'0�F:����8��6�6�Љ�u� ��4}� ��N�{����,,C"�"�� R⫎�����D�Kώ��Y^��WR��^T�Z�?,f{��0�pq0�1��vͭ�jt�~ڝ� ���
�0�^��Ȋ���X�x`��$j���1��Nfy��3�g�رz�듆U��=��E�"��v�n[^h�j[f�d�]�h�̑��)�UVW�}�b�m�I:�e��J��B�x�1��7MWt\��4���-��D�ca�c��u��E�{�.�+�K@���"�� ��Z��xV�]���̘���w>g�f�[���[�_��F�Gm��?^P���x0:��N߂��*x<�4nh�Bw�m�[�1�Y����C4.�Q��}�H����'K�7�+"�8�r��W	X���#�œ�Y���=ɛ�4W�
(Kf�)��+�E�񵂣���{��!���x-��}��~�d+W������<;��n�uR3x1��VTt�Y�J��������_x��ɏ�N��ة:�I7���T���v��f��7�y"SrR���̚Xt������vKa����K6����eK1ob��<�F,+�k:��l�q=|J��l�bi�\~ѯ��!�ى�HsO�w��M�]�)iB���";Ylq~��r8�G�p*����<S��� �tGx�20�0�S�Sy��G����>*��%��pf ���{��j?�)��: �ly�(�D�=R�A��/Z;�EgQ�[�]bv��|נ�u�?�"�ǽN�#��={H9�������ǰ�$}��U�V4�]5ˢ_�'S���q�L�����c�֯���Փ��X�ɭL��U���J�3���uj*�k�����lk���n�z��*��q�l�l�E� =Z�ڤ�_�j���g�)WR�q�����2d>�o���K,��ތ"�K���SpE�(��ޅ�dHN�,^��5�B��0ē�.�����+"�9|yk8r�q�]�Lנg<�/��b������@ɀryM���=�Z��7�p�+���Y��Ր�@�o��2�N��=��nf͊xq��7�lF��`ZƆ�(�����2āi�!ƫ��A��p��
�X?�e�X�����D��%s��~�ƇXg{,���	��y��zk��|�w&�~e��[ ��ձ8�C�7��R)/��\�)���*��GҰ5�T�����St�^�Zhd&�͇$񫯢�/��.��ߴx��W.��d #IҊ���7�������X��ֻ�v)a�E�sih;�A<�3�U���빡�NI��$n^��V��¨@Rb��sK��� ��\E'ם��UL��L���O���;���6�I ������{Fx�Cȷ57h�a8����{�C��Fl�	O�.`G1Zz��oE9"�v�si�m@����O(��a��d.t��A��1�E��w/�3$�G���@�k}��"�ieH+5֙��
a��=ؠ�oX�R)�����5D�y�3{������#���e�*��$����a7�/�k��k��C.cƸҥ%
v��N�^����鵴w��_���S\V��]#R��	4����Ѥ0�p�\؇�ߐ�0u�e�m0��qy�pO�Dv_�l��YWކ`��ӽ����۷5����$<����q04P���N�d�v��{��v���0�~!y5�1���Q$�U�V�"�X8{'cT�1�d� �zu@��Wtk�O������bo_	BE������p{��_:~= `�hJ��a���]�'�ĝ�������d?n��T̖�·
=��|ڔo\ۨ�"�J����w�wv�*FKP���C��3[�2�(��?�_�,��R�T�\�^}T�p؍��\�4)Xr=Пu�BF��UDM���)�z��mj�n��� ɐ�V�5�"N���\��ֲ{���r6���v���l��K��vя* �}h�4u��/b�m��W*0��,��mvB�.�VZ�E`�4�Jd�S(eXɖ^�o�R�O������
��l`r=V��Tp���y (٧���.{Q�^U�N����b��z�W���t��E��>p)v��<`���4�3��vd�W�5l�b���:t,�J�Mw�L�H�Pg��Y�r�{�7R"_�δ����4�~UBӼ��#b%
���u �����1k���9�в*V5G�[�C���9�L�\Z�g3ϐ��ď����GS��pϻ�N�D��L���GQ�I��>X�BcU�o�:`�s��"p<,�r�|�Α��@>+�i�I�;�����R��.���q/ڊX��RΘ��ם�x
+/�\N�q0#�OE�{Od����h]b݄�f���{>q��H'��!�=�Em�}������%˙�U�̠�G?!	(���a����)�u��ڮ��p穥ōp7&�Q/�Jøz��!wTl�;�x\P���ף3��&ܙ��ƵOz����A��ӛ�Ze
bJҸ�*���s����xˀ����;!wiq���P��E�CqB��-^(^���Iq�w��
��s��}�{�aɗ=�֬�w͚���Ʒ����#"?�i�hHݢ��R_��9.�bؿ�\I�7������yb�<��<��h��뼍p��	�aS����n���y`����q�(I�_\C����[�(IZ�J-,f¿��Kܵ8d[��2��mo��ʽ[m&��|5�1]�����}�O��Y���i+ A"Q[^�E5�yl����RȐ]V�7� �A9�fn�%e�z痞�Y��h0B���EĆ�t����� ����A�_3_w2���+�S�L���te"+�����rl��]��bj/�i�c~���B��5
�j�m�!y0�lA�z&~�����'}�8O�^8wk/�s���	��f|�Q�xw��s&8T/��j��x���~\���q��ܑn�X���\�C�{��;��%��m��)��D��$O�N�C��/����xFˠ+��ǆ�{;�܇�̞�����b3[�u�߯hh��b�+j7��ޔ�~0ꯏL9&���҃W�z�|��Q��i�z-V��6����؂uST���?r��n�u�`�uvη��=���p�i��	�}����~o�+���	.&{gGV}���o��ơA����P�<���#E�9Ė�^�(b����W����ɲh��C^�?|{����q0��e�>������������ې��S휚��C9krJv���HY���X������X��g4��>)�I��>;�߿���Q���t�v7���7��!��&vɞɀ�>��M�����������N"������2�\�V�M�pY��ɑ�<==N���u당N�]��*%C�j4�CBFRX�d��-�=�K�U�-g�e�vr@XTt�I���f��aĦ�Խ»��%���`���&cU�e�j���sr4�)��~ oØݏL2�t����l�LI&��j 6c�+$�avc!���%�C��cw��τq��q!RkJ?�V�!��yԞ��$�`��W=ܽ=��
�^�4Oy�
/n��7�[k)��԰�̼��Kqq�}֑�8֗'UfeV?l�x��J3��?C���Ac�<��6������7���!	|'�']��uV�����t�2g��溁�f,�ոH�����>��}�s��lL�ꓲ6�]��B���-��L�����ad� ��z\vj�K� ;Sg��@�9/2W ���]I���{��56�
G���� Ά�!x�y~����ք���~m:��%W��O��3;�,�ʽ�U{N5��z>W�g��j��;�wf	��?z�"A��6������#��SDN�D�ø���z��nάq�݇�/L��i�At
�b5�U~����a�,?�ⷻ��-$�#>��f��8�Bu��y�I��"�����v[uEC��&�u;]i���#!���8�[|X/�NOx���_�պ��jئ�2�2�a�&Ӌi���bO��#�e��#�ҫ��!�,2{OR�B[���V� r�ي��IϖwU�@zs.�I�C1��" ��c�%�:!O�`&�I�����q!
�`05M"�"��/���Khw^Ph����MoS��$��(�%$z�4�$���_�z��필�b��v8,Rw����NS�I\�<+?LÄ�@{�����x3]�|V��`�0_bV���'��
�}36@*fd��c��`F��;|E�T����H��|;����i@�1I ���*�g\ɢ�'v��xY���V 
M��`��S A�U����w�9|�$ru1��/��j�ޝ&��M�|�	
Jѽ1�ӷ�᜿ M<���Ny�a�"�b_)���y���G��GSI�ZΎpa��/�Ȱ�>��r�z��.U�<����$�� �cX�>����f����1� ŷ��;4_V~���z�z��	���{�󩙌 ��j5�L�e�u�lS#1�X5�
��/d�ih�$�k�Ze7��?�BlWt�Mߺ��"8�'3k~��-����vu���{�n�}�s�9E�V�h�'4h�rw^89:Rg�=��ؐs
1���6z�T[���pX���o��lݞOEtA��j���HS��-5o�	琟t�*�*Fu�Ot��kr2�����cL��t���Ս��7�g~@�҉�Z����"���n�"�B�k�MoD�r�R��I�O/~��X>�V�"ۘ��'�����#��'�)O8Q�W^��!�h��CO�G�����J.��i��߂��T��g�n��&[����x8~�Wg��� �>�D�H�A�_�UJ��Um.&��g�� Tl@���wU*��G������̌��[ZG~cn�/��bt4���q#�*E,*�Z�g'3��������D����~a����Q�Y�8w��Ӱ����m,x�/��d�k�RV���@d��q� �����;�$�,���#��@Bg�s���S%x�T->�7c\���ИZk�J��ί�h̤�Ov��}8HDS=�3�l�I�q6}�uz{������t�3�F�Џ��<=NvD��:��ٹ��Z{��5)��ZE�>�w؉Ǚ�+2�S\ct��
D�(�j��l�YD#�����okD?r	��E���	��&2��ՁW��oV�mz��~ŧ�b�G����@�)=9�4Kh��	�����|���:{\�$;�M��V�{�#ҿ�x�g]�K��z���vFK�),|�0�1W���;?�v3��ֵkև>����/�o1�j�c�4�#۟�(VclG%܆ۂ��3�Ê��L?C|j��c�h$�A� 
ǲ�8���ϫ:�t� ��x�1�h켺�`@��Y�T ��u}��+^����&޻��ݗ/j'b��p�M��55mM{� vv`�.LFtRz��&��wj�c�x^v����W��}(�N$����Z>�>�pK1J|n�=C����W��H_c� H/�޽?�9�ڛgxk�QXY��D'p��Y�.`���mp+]���I1�IY5�49�|
b�߿퇽c
��Ri�����c� ��eDI�5Iqz>j�`/ݵ��c�6o��7���O����x7�v��_ ��c�(蟯u�~4�!�=�Ә�!��@�r��Y0�E@M@�w�٤{�����i�Sq[�%3R�{	�ޣ�w��H'U2>��䜃�t��7��J(�E�=ݍP'U��K�}��/{Y��ޑeA����|6\L�y�r�8^�'}R�V�<�n,�uY� �ȭ��a�S֦�^��|����ס �Y*���E9:�޶
3�#)W�r�N�Tť�;W�Ӱ�Ƞ,��XPe�9V���xqS�nD=%��%�?1�m�e��u�n��?6����K��7�<�i?j��%)C�����Q�2����W�;���|7,$Q����˕�-�Z��D��9�6�[���e�m<�z4�SQ,4�5V�vy���d�"͵?$��a�ġ�L[E�(�,R�������[�c5�U;�� �#��ry��
;�gm�@N��I){D���'z�Mo��������o�(Bb�yb��R�^#���L�nE����)�Ul��Mu�u�h"C�ix����y��n�᧿;U;XX��LL��d�,��N#�fQn&|	AY�#U���� �'M�O�Ϳ�z��%�a�bBM)�o��t�-~X�_mf�+J��A�q<��� �c��c��z�4
�e3���G�T�yC1I�X��ԧk�ś���cz�k�HI��k
F��lHm�-�=y�;)�O�)����
]�A��M�3�7���N��zz�UTͧ��
�/d�:��U�~4�%E���	.w*
KM��wb��k�B�</Z3$1ŗ��~w�Q<���NPzȑJ���f��qQ�2�z��=M����۳�?�a?�c,A}{�6l��Q�?g �-�|��v�/n<��3�8�)�"y������@D�pZ��N��b����q�_MOޥ��#	P��5����WU08XJI!ykT�/�q��{������ك_�Uˑܝ�� �YИB벙����F���Qڑ�O-k���BX��79����Jʊ�e�γ,�\�� iUG�@쇯�YT�	w��Q������O_p)ڦ����"I���ƾ��lN���k�HR�吋�v��+�ʹ��Hʉ�k�:�JQ2�~�|��:x+6�lo_�:������J��@��&��G"�n�'��u��ȋ�GE��V��x�z�bY$^T�1?��~SsF����~�=F*&� 
ls�Q����>��g�p�s~D��ʃb����Pv7�g̿gS9I�ї���Bς�0�L��F���?���E�I�'�iZ_
(����������eW\ �w+Կ�F�7��;����N~��0����E�������΂�ˆ W' N�a�V�Å܅�k��G�k��a��ݒ���§ʠ���ҟv�F?��ߢ�<�r̿�!۟����'f�4�[�����w��:=����b|��2ڀҔx|��Uh��l�Þ���=_("J����;�����������F��п^ �i&n�z���s��E=ʘ}�^�f�m��lg"u�J�w��H��q�Y��}6��eE!d���xjFg�`ֹ������#E�5��ð�Zq}dJ%�:�x�.)�
��m���L���Ǧ����zv����$%d���Oj��ϫ>�:=/V��OW��̡�,�L��*����wH��{����vn�dP�V��\�W1c(y$ZR�F,�[�#0O�M�����
)k�yqñ��?ô�:w:�:��R�i��� ��1�};��L���������ʵ�⥲�Y8�g/���4*~�G����4�Ύ8V%kʘZ=kU[M2\�GP�B�u�*�����F�F��G�?��h�P{Z�c�[/�D�����CG�I8�47���I6[��|b��H��BAU�)d�q�6FZ%�L@��M�萋��{.m�~�N�>��z5NHH�a��	D���C.¥͒�W?�vq���ɄU�u���y���H�[.#�5z�ݟ��xfD̷�Ae9�a�?���v8����*�EP�]"����yK��U��)j�� � �$ �$:{ ��X$�]/�5C�>��J�vq��B<�+�?���̞��Vn</ax,�{_�.�<���W��Jb�܀�ޣ98#D4Jf�`�L���H���5�T��/ڭ`�2�*8<HB�R���b��;<)i���	�7\>�^�Þ�{�����6�5f�<��'�u���W��Z���=��ȼ���b�)�i�0���!�Hd�>B��8Q:xJ��B�`�`_�؉u9��f���wF.�p�?��O*�#��4Z���}`U�{_k_z�0Y4"����Qc��䐨���O8���=�y9��I�6����fօ�^(I��4G��F�T�{|�¯*m��k��v���p�h+W:�)�唀��Љ�u.m���K�͜;E�[�Z��*&��g1>^
��Ey��RF���䨒C����%�>n�oQ8��,[��l<�I��bɎ����oX�v=���T�p��Y���.�4M�P e1ׄ��@X���Z��/��ө�����"z����K2%����ki�#�ZI<���:D�-/�g������H��b���a-�S��p����&��9�A>�sNiEEw����t�s�k
-�����-�P\\�U�l�?[��M����oڍ�йR(o�{폗�9�:�L|�&is���N;q�n�z�ţ�EA��I�P�.N"M}���u���B̶r�}5�RtUD�^�f����a��0��0�'�������4{�=�g�9M �!X�X��A�x��r�}��V�*ԕ�%䑖��=LB��������WZ��ȕ�lo��5��#�ـ��[�JSF;����jԉPAE�o����q��u�]>�EL�����޷䬿�𛀯/�MM�w��Ƥz��L"�1�="}Z���Q?�	ռ�v�m�9v{o����Y�c�+tC�������q��c/.~=Iv���R
�ګ p��P��6$h�T!����*�Ѵxvk�jN��8N��}>��=�B������f�t�Q�\��=�N`�zDX���/�}�Q�T�.�)�_�7,�$�_�f��Y-PBt��A�ߟ\ǩ�Y��Q':#%#�[���jmɼP��<~�������o�/�׽k��/�+�}5�������}�2�;�!��@�o�**C<?E��U�I�x��
�
��M��ssd=}r?+�H���tB�o�-�;@s͟Y�{.�Ϋ�֭M�4������<�N\T�u���g��4:o�w+���Q��fi��=?���]ќ�S�_��e�$d>#T92P$���ȿ�9ҍ�ir_;�Z�)���ְq�!}��pn9X�'ȼ��4��U޼|��!-��w�z�������c�D���ĵ�<�:ÿ���uv=Z�}>��?�u��)Ǣ��	�"I$�)x�����wi /.�i�Hz� �Ȓ�v��*��P�n��+j����y����2Օ���D��~+��7ᤊ�ު���fx�Z)F����ʧK��<�����k4���g�'���8�>
�	��Jڦ��D���n��x�B�θ�)bXʩ�d�=�Y����v����`�-A� 8�)���(z9W`̩Z��~�l@�"KD��ɥ��	n`�3ka�em�$���\L��~l��(y8��r���f����l����C�J�n��Lt�)iW_m2�<����24'gj?�C���)��l���+w�����^��ޛ��w�/�x|C]	�.}Zt>����!��|�����M�}����$��ßtvy�f�편|���5��s; �����6�V�������N�y��ڧ�Ō�hK��)�n���+���y�E�o*K1_Jp�����<�������h9vK6V�~��/Y�͕u#�Gr�g�͔W^�D{9���3�SF!VS,�w�_?h%(�X ��� 3W�Q��;'+|)��J{u�����o�\��!Y�����n�դ��eד]� d��� |���=2�4%��=�Ռ�K�P�/߽t��D�E��p�R�I��jdK�_�>��i�Kf�n-�s/�[�|:���.��vO*���0�܌]�����)���@c��U�Օ}����CbU? ���W:
�&�x�g��?V`��­i$����#ϱ����s;
<3�8��pwi��{Q@�v�0�ꮌy�QG���C����C�"������Yۊ9��"u
�3ф����д���(釖���L��?����_%E���|B�a��R��t^���r�s>�h�sD���Ai��5����i���"@*�B�C�1�p��j�b�W"��23;k֟E굱l�Q�#��|[{:S��-% 6e�P�G =|�ڑ��&�tlϥ�6�1����fm~�����2��N6фʅ-�`Ր7]ޖCm�~E7BL�j!O������Tk��e`��
��;L��,�Cۂ7�[N�˺˟��*_ɠîs����)��k����ζ�)����
�(^μ�*�V�ZB@�x��Te�AF�Е��7|���U��o:,��Xؾ��#Q�����]���)>U�t�׎����V�������e��uƠ�� #t�8�wOߕ�F2�n9����?�:?���9�"��|�&�=.�P$�/����!�S	F�,��i��X���NG�:��AF�(g}���tM�{<l�s�m��U�XeS1�
����}��wH�=�Ʋ�%K�OY��߶[��f��O��p��x_�
�$�����:��cs�LLx]P}�� �#/~�C6���)!��p�r�)=܂�2��c�l�:{��	KZ�J�t���X;����~��K����x�G&ɇ�gTbf��7�#��H8�G��o.(���ey"��y>$]�o�i?�#��U�����n���� ��>�#4$��T~'�dWxC�W�s���;On.f��S4_�����j��[u��sԡ���
�Kv~�Ngr�����Vk�Eu�>ڿ=�
����#��)����1����F^���7ABp���^��V�?�Ѕ,��3���Ob R����M��F4
Z#/w��vj4�Ee�_���<���I�ZG���z8FX����#3_��,R��\1BoU�v(�[+]z�
���$�~��Xs���U^�@��5�VL;K#�;J��@7Z�5�<p����K�4���M���彠�X5�8���#�������*}��uУ�cjI����~�����-m�N�n����{&�Q7e��^��09<�A8��q�0���3B�O��Rr~��&z7믎�	�=T^%�U������j�.���.��??��c��#h����H�wk�?���#����lx�.�q2�( ����<2���9e}��>�#@e�JR0�K�3��;5�ùP�uJED�أVM��-Ǉ��'��F�(DTޫ5ͮՋ��N3������W�\p��M�a)9�Ab0'��^f^(&�S ����>�\�P7T�0���`��jr�jO�d�̔���z�N�o����zO���L�,P��{��A������jqI(�����
����~�T�E�0-�dI����F-�BɎgƷ����E0����6�I�w���S�`��?כړ�..ђ�����W,_�*�7�T'�c51g�9w�@r�O��7=��ܯ�=D�u'����w���/k&Ó�H��~�2[�⶗����&Z恹{�j[�����~�������N�q�\��CE�����pO������]�	Wi�;GA�.B�^ID?��kգ _O@*���V�!���Q�q�^H��S���P剻��p���{}��dx�2��^G��N�~I�P�V���x�8�Y������eHͷ+5`��\�QP��뿫G"����3����6^�g:l8�L1fB�ƽux�x�
���0r�-��<�K ��PΑǖROMM?J���wzf�]>�<���yM^	��`bYk+F�w�b]�l�k/��c&�ر�I0r���JO3��X����?��'��5m
����p�`��))�v�$q�7�-�_�SG�^�Fr�؏}g�w��|T)���� 8�Sm�q8�>z��K�|6fG�C!ފFJ��+Hԧ���ʇ��.�������8���<����\����SSQ95������.����S���)Ȝ8Y��Aٵ�༿�G:��.M�n���\]֓���K��c��KL��]���sQ0E2�{U��h4췌j�1S�b=��{�R�cw�s���<jq�P��X�y�dj�w�Y�|��{>�����^��S�����v}:�l�:@�#�WТ�ִ#�4�a@=g���ֹ��qȝ�����q�E���jL��|��V6fZ��x���"e����~.�7���n7��>Y����1���W� oÚU�)���J�(u���e�G�ϼz��in���K0iߤu�WU���}��?9�7�T��g����e�zVyOve״�����U	m�G�I�q�1�x8��^��úWQ?�<̌�e�D�gdj=��*���f+Ycrm��7�)YǄ�����'z����N2�ZO+�$z�g�3W���h�C�j�B����8��rc�J�mf-��'�E����8�.���B̿Q.8���3�$QN�恽��DO�8S���&=�B,���Z� "�x��������,c�ǒ�I^��i���~�lؼ��ΑQ��*��L��D�/�j�Z�}F�4��T�h��ǐ3o[��pMN(2�G/�&�d�"�x�ј���n����Bc�%>5���/\�@'J����LV|�Ϳ�+��u��j���'O���5�!���/���-�ȶ3�j!�w��Z�d���� ���X�`x��Y��w���%�Z}�k"��4�6J;�Tٗ�1�?�?�5����5�`�@��\�FV�8]͋^SArE�ц�h��*�t��(O�	B@Ic�>�1�E�F�������0��i�S*����[� z')��	�F���������JR������G���ג�^@O5�G�h�G!���öF~��ߊ>�Bh�><x���ׂ�8z������M��&s/3�>��gn���B���Fc�h�I�ٓCX�x���7�S�5������︓�ȸj�Y���^�Q�g@O�O��D�7RǍi�4}O�=���	�d�}�#1�'�`EVUr��a�[sN���`^��?�̓"���j�9+9ޔHyֳn�Y r�.`am^�i�y��%P�Thi�)�:!xɛ*�bAl�0	1��NV�B4YM�jD�ke1�x��O����J����JK{RO
�/��:�֤��}�PM�"�&m�����̵�N��p�T�� ��6�Z��ed9���r�ls�\�7\0�4����_�덩����}J��`I�����8�{���k�"�bd$KZX~O������b3�������|�1>��f�ms诃)�6�-S��O���c4�v�H�Em������L"�@������0˥X�~B���K�1U	C@)TyD�V?����7��e����Y��«�w���Th�`�Ir���X�h���;�?��̒o��������y�)��
�Zq�!vYn9�I�ܬl�wx�Ocb�m����"!چ�QVl4�C��l9��`=�>$��Ǣ�N�`KA�`w*eD��)VA-Adm�C�r��D�:�K��*Ƞ�'�v0�J�~2hp�T���F�H�~~,��(0���CM#cW%�NU{Ei�����	��?�m�C+�ޡ��������Z�Jb������t��S��^��+�W����?gLPL���%n�^��x��>�./.��N�m���DQm����8��0�[y����;�B��N��_}0X�(����&�ʞU�]�N�� f����N��8�əD0�t�D�U�|���!��ɹdO�Z�������:����j��X<[<��q�C�i�i�/�<Kb������b��d�(y-x6n���X!��Oy���%��YL�kD�}���Y��{���/�T&�Pt
�w=;�)�2�F��1:�c7E{����V����=-�O�OZp �|�RLS���R6��ւZ3D�EP*$gb�:������K�	{7X=	ps!;%k�z���i�	�3Yǎ]�0��lWIYds��� 7���KD�t��9�A%���dT��l��w������@�/����l��G���;!�9��q"l��g�����3�wa��/ɂ���QW�н%?h
����F$M��@}��8b7�A�Uh4h�5տ��:�v��f	t��{#�3�^xل���q����!��I�-C�r[i��/kCy�zd�g�<�'Fs�������1�d�h#���.,$��0h��ፊ��%�pN�F�4T�Օ�q�4���[���q�[�g>�x����<pI�?Qj2�C��DB��Q����\����3�ЊX2����x�ߢ(��B�=��u������j�ɜ�P�E'(���	}�.a�Ő�i� .Ji`������� ѽ|�+��P�!��q��ؒ�-d�OgZ���Mbyx�b�;�L���s̜��N�;BR�lI|� �wϖ{�=:]����K��d�m�"շ��X�C
K�UY�d˼r<�^SL�����W�y%(��;o��Wڭq��7ß�"{��i/ҚQG6�\�l�0���nP|�0jx�DS*r�]_8~��]=�"���:b�|�ø�e�6�	!�u2�8��it�K�y)��b�B�`���@<I]���X����ߪ.6�Wm�q���Ѽ{�I~c�5Z�{)�����K	ö��hKwY/cH�3�V��u�N�a~i�<1K��r�C�_������ɕ!f�X�hK����"՘��7w�ǌ]?y�v����(�t�!�gQ�'��Ʊ?9M��f�}��l�wE�mŻ�����S�1�E���Ͷ���r4�9�a��t��lM��o�B�ʮ��K1!% �A;���I��V�-ۄjܚ}[�����2J�ꦠs�~k��-H���	��*��
��	���:m�[����6��J���&���+0���$�n�v|�	���a��[Rcyl�#��T� ��߄oUړ�8k�ڝ�/�+D�9EBa��A������DMb	w���k��v�X �8?��740�(�
Sށ)�(��|�,��s SY�lr���_���伀���҂��@�&i�z�~ylGl���n�s�{�1��l��Y���O>9�"n�C/�P� �&��ܞh=��.ʹ.��~[	��?����^΂=D�&��U[C�5�Mf�����)9���z��O�1$����թyRuhow����J�<�<#gc���?��l�O���&��� N�bW(���fH����W��@�m?��Vڅ������]~'[����-cr!p��~ϖKm?�{|�7��)ߎ�������%���'{����`���G=F�ЗU��aZ�Q���%2��k�[�L��ަ.��|\���8!lp���^�wn.����+O�o���	�Q��� �����>3����޲��Б$)����w6�=��5��(~�䉜>�l�pv��:��[��5+��v�H�eyۺ�r/��;�[�ByO�NT���G�{^�8q�
����톯�g��R�+=�gw���+Η_g��b'�h�v2u�����n�<��B�8�'�X"��kF|;�,���\Zs�3�2�N�j	g���d'L�Bߺr5�c�8��A���ӭ'-���F&�\�%Nio�������J4��k�</�����d����Yk�d�ҹU��ܞy�jˤ}�Rj.�*a�A�V�Pn��	+��f�d�Ԟǒe3<�6�X��.��4Ee�*�qS��	l�4��@ͱ�3E:�y`�1&�:af���;�E��'�-2�+���'R'�����Ҷ���4eF&&�fȟ��	(]N �T���A��2Xs��]�5�ݽ������N�{!
C΄O&f�����s~�1��a����U~4;�+�?D��Q]Pvx7�F35�[�2*�ۚ���v���h,�ȴ�b���B�
���|sVi^�V��zn��	h|>u�ܟy�f��_��ul���͏ߔ],��u+su��S�Fx����}Ez����G�H[71�g�&~7�Ў+�|yޏLn�Q���!2���C�~Q
����!��C��.��šAe�.=�N����R9D޾r��Rr�WX-.�������ԧR���p�1�㠹�����_�8C��-u�~��c5B�#�����.e\Z���ؘ�K���p�K�k_�f^V-�}��A�f���j��N���Ji��IRx��Xp ���	��\L��ڢ���_���L���YM�UAڶ���~�|W\����n�BZV-����S���8	՞�w��~4�P9������H�F����+���%�ˍ431L�
cf�-�/�rPz���(�m��U&�r9���Q�!e�#��c�8�M�Se�B6�z>�~䙷i�����{�TR-|�Bu�O�_E��\����(W�@h��@XN� ��Yٲ�"�.{���D�ԫ�l\��t1�.p�uK����+����p<�ꞿ��n	������v��z���`[�'b�h+�r��S�~o���3?蟤./;��Vtg��A���N�k��Խf��V���2����,�:3 ;�h֌�����Nf��Y r�y�Z��g�;�Zn������I�	ZHuA�t{��|p��KX���,�y7�Z�T��ν��]��LSpo�̛C\��?2��i\�,ҡ�A��.�����Ѭ��)G�4m(��,׶,1H:tq��Vwh���M�s����s�7~��[�S!A=C+������V}wP+x�­H퇒�jfz1V؏d{H^����$�p�Z���ʊ���/�)j�Ǻ@F�.�X@7w�i�L�췖���t4�D�Q�2�-��z��"ʚh�J�9>+�8i�|@n6>��G�4�^?�J��C3t�K�Y�D���[O�wӽtn<�ֻ����n�T+*(:5	`�ʃ<Z���SzA$��<�z����B�6>�ほ<W��:_DB�[9�UZ��/�M��*v���\�|�ѭ������)����^Dp*m�F*�/������04s�������th��^x���P����0"D�"�:O4X91YLЖ)D��D��P���gK��+x7�s7���5l�3��)�cf;���3��Fx���}K�͏5kѭ�x�R��u;��._o�坛!�	����YY$�UB�]71L����]-�FJR�:҂����;]]�OI}�'���\Y�d��Qk��l�&LV�$T�fޏ��J'q�U���L�_�AsK��Q��H�Z7�7 �ش����Z�S�]�G-�#Z^,�N�Z��B��%g�H�
%������U��l��e�Xd�On�E*�KK�WH�S]N�Z7�I�@35Uѯ9����<��|@�����*���WB���,u�ܔR����?R��v�w�KI�xSJ�KX�c��� aۭZ]z�2��S�kږ����ۇf�<�o����Ï����w~"�vη����p~VZ^}Sͼ�
�G��2>�zF)1ށ��ƽe�=��6z&�!��%���󵽄�+�f�޴H6�-W�Ґ��I��ٷ[zd�Y�{)���f�~z0Y�Ӵ;�;߻-�lv����b{0��A	-����3sj��g�-�\����,Sٿ�.���_^�l��ֿ�ŷ�(4����l���>��P������w��K�8�7��"���s�R�l]w�F��4����j��S�O��5˽b�0����Ʊ�. m'j^�q��7{'y;�O�R9�Ju�X�Ȱx[3L߆�4+]ݢP}�"8��c̓��ϝ�y��)���+�TT�jm-�� ���#۱�7g�w����}����;׾6f��:V�=]�='Q�����<)uI~ڒ�-~�JP�����w/]��)�((����<!̶G^����&*�zЗ�ʍh�6n}} �\X[&��"���ؕKt�KT����+CK�����������Q��U�Sƕ��3D�#ƙg�j/�Fk]�D��'467X�8��Fth�W����1Ix��JL�i�٪2�|
��d�bs"��͏ҟ��~�J�v�+�>�r��'����[�O>4��$���_��е��4q��~�\��ݛ�@R_�-޺��T�쩎�;l{�\B?
5!���E(����>S�xϵ2ۑ����k��'u��ų��(_�dgteK�.��2�7e�B�9��W�vf�oW�}�/ZW��(�S8J�_o�>H�������C7���}0~�w�%2*.���|��W¾wf
�P{Q�����ʠ[����٧\�5�TC�$�u��EHo^����4�W�P��盾s7kۖ��`�N�;��}=	8�F��
�|?� (��]��z7�nf	^����wt�/N��XA�|�xoK�doP�ACQs�#�ez@�B��`���,�g��q_m����޻��:Y���9�`ltb�4��g����z��2��x��mh*��U�B���چ~\^�M	�����	!��}6r#��"��6��F$�4ֿ�_;���%���T����c�e�@�|�����@>��˹푀R�[J�4]-~_[�2�v���8��qg�-�qg%6��\Г�1�B����U�ͤ��h_i��$g�]eؒ߰ɏ'1�\B��w�R�|2�/m��[q����\�������]1'+5m���=S������ӗ���:�� ��V�d�E $sH�p��U?kn������S�r��RQE�<}7�?����Z�#���c�u��F��Nv���L�j��K'�����cVE�6+2 ��(��t}�~�@}3���t������{��7�� �{�[��8k!l�!P�K�c���+�C�����7s^+��)��}�f��<=4���3���h~ӡS�N��r����1��d��?�E(���"=��=���a2��S�'JB��A�,1}>�V�#^&��v˯Q5;��P9E��N�ns��-̐gO�E�����N�,5��`���1ϫi��ٹ�Sٹ�_�haV��������W�7n��Ej�WU�	iM�2�]����\F�i�Ѕ�r-Qp/gdb4߶��������=6���~��NLGꉚK�}�|��ʥ H�p~�.|���)��+
Q)�!�4?5k���1���K���&2g,���f�t��}@�TR�!" �5BD�R�A����-L�;%���1J�ƀ/�����׎c����{��{��K\�H�eTţư�׾��I���RiDkp��u�ו�D��u�탧���B��F��0���_�5�Q(:.H�iu�5}L�Y���[k"�r�&}}u@M�G���O�Z���F�<�B&h�0��!��R�u�CS��ɽdz^���<�\ 
p$U�j���ڽ�K3�z��K�z[6D�h=ɪ��������o�MU�|+�Pf/���6l��9�+3�t?{;�n�suK��C�N�Ktkv;_<J��״���΀��|�@�fm1a�]/��)OC֊��7��������dq�u�@F ��~�u���4�:�@��!�\Ji�7����U=�W�����S����̝��� ƛ����ԦI�泒G}R'��KI�VmD�N/ӾVy���^X��#/w�q�n�S-�?a{No�F4*/1׿�\��QA��b�[����YC��=]��L�+���'l��*eT���m��a�~�۱[~���,Y���!m 9|����Rw35���(+�/^]�`4@6�����9��#:�R�A�kL��cg��[���d��Q��LuSn]pWy3_��SH�{:U� ��$'�~Ȇ/�@(^yQ���w����'ź6s��<L9����(qcB�(���A�&��-��,���N�bnU���j���岟�x��0�d�z�ر��r�������Bc��g�2�=0�)~Y /]X&��(��G=Է��:�L��J�=H	��13�Uk�oA~BP,�r��"%P�8�_H����*�� �Nߒ՘�t�}@�A"������(*�9EМk@�g]|�>+��U΢r�Q�� [H"'x�О��>����&��Q!a��4�AwN��G�_��ծ�c$�R1��,@��`�+d�~c��\��+?C/5}.7�t�,�6��-�u��h@���x��'Aϫז~�����3�:t1G[k�_�3J���K"D~����ܝ)YZq�Փv�&�T��v�/��y��ڜ�tD�lϡ���Wq�����C���W=/i�Ǌ��*8�i��cBfέ9)�k$���ɱ�0^w���I�peV���eG?�뎖3G��#�V�/;}�V��n�,G��.'g�X�.cX�ʦ��d���>[�BUG$����r_zN��]����[�_�˭8�^���є(� �X��R�)�rtzQ�}V5���?��Z�3|p9J���1������ys5W�,��{�%,��J�oE�FK�A�V�C�.�2���/�$x(���@��������L~ɵ�R5��"���M	B� Q�~<L�f������39��|���_�@kd�Y��$�q�EESƢs}3(�s鿗�˹�f�&�%�XYZKLF7�a��J��{��*�?+Ŧ���rܙ[��ٟ�q��y$�_�</K�W�V�xv��aP��W�����'���ü~�~��/_��������BT���w��4�i�9T6m�8�Ĺ-%��s0�6��Z{l޻�~��3&i�p��Rޠ���x���L �\^^�H�t��y�
⇜�`����Hb�b����A��r]3��c��;3���t�����?;��]G?V��?a1G�@+�gqT	r�����*Ri�^(c�L�8��Z�HK�vx�amzoX�^޻t)\�R_F�R<(Oϐ�F���2�{Z�HRh�ϪE��ޅ�r~���ET��4<�3��f������>d4�xO(H��o����ӭ>^�lV�k� :����jW�/����+��Qi�[b����l'LQ�KEp�n���L���,��{~"'T=�J�w��\��	��`���K��T�'!_0)���l���� f5�� �$��x%�b�:�Sy���G���sy^,VH��NRms�lY��+Y����{uk��k[CGN���cX���`��?�-ߙ���G,����V�2d������,�%�m|��f�Z�>��tR2�-/�(-��r&>���A>�>p�X?����8���R_��w��1L?��7 �$`Y	�5���!�+�Z�[�x��N^]?��q�/����VUM+���3������U��8�=�[�;u駟�����.)�51�}���`�@&�
]Lc�h+���)����bu��"h�2f�-�{k�"KzǷ���݂J��.k�`nB��~��K�1�z������Sb����T�_��^CO�gc�4������[�(�C�^�/׊8��(D�=�Q̈́M�Q%�;�Mlܪ��yH��x���u��xmii�k�w�c��I��A�n(�]-�)_Ⱦ�Y�<EAn��Q���1�r�Τi��o�!�7��W�l|@�On�CH�W�(]�<�}�����>�wm�߷K�tUb������ ����5K��31�4�xd�/�G�w�|��&R@�>XU��T��⦸�������9����׫���Q��uo'V{�R&Xu��_�������j�OOkŲ��kZL�2|$а�l#X|J�nf����R�@�C��?Z�d�!�Ӄ�V��P7�lo�I��E�/���g�(���g��kݳ?G�\\=d�=�������?:�����#����H治��ߩl�&����j6�Բ߷z<��wd(c�$�_�"�����8 �WK��\�}�ׂ�䱱 �D�����;�ep����^/W�����jc{r-[%��"͐l^��������r�Z�u��-��Z�!�ݲ�h���,����^�H��3װr�c�K �ᡶz�>@�/ӛ�9�}#�z1��Q��G���^Ä�J"��)��/f��*��� z",<��u2��@���z�,��IӶV�Y�������ΥHU,ʾ��J�ǃSq�j�E�j.��/Ɇ���D2��U�~xn�g�pꮮdT89��y��E��`S�:?��Y{[����#l�����������u����D��m�0w��#�ߗ3a�e���p�Kq6�(06/�x�,Ş;��Xs\66%x�QEl�fȲK�X�=����c6
��+�w~�hu����+��[+���*�MnW�0+YHL��5 O�s��tx��B��A60��HQ*�I)�%�&�EI�]_�>A�_��>-��ѝҪ����/ۢS� ��pi��&��|�&{|B����v�Z�����0'��_�{�|)��h/�B��}/�1(�@׹��$�U�7諛Ľ��R�^��z�J�%���nTr����h�]�'�;�sW��o7��@��ko����7d�� �۔�/>df����� ������8�
QF�5������ϋ5!=Q2�g~H���y��f1�q�c��d���FU�5�-MiD��h!�4T�+j���[�Pu>Q���{λ����k�De��8KI=#}hA��Z�ʎ���S��:���1
߬�8��N�y�]3�'��$I�(,�����N�O�k�I#�g�LfvF�kY�IE�Uï�E��K�2��JK7��Z"�oU�n�m(�R��",��s�jm�cl�|GY*�x~_���S9 4� K��V�"�b�Mw��C��KuN�Lj)~ ��]˿�Z<擬��&��_1��z�RQhvl�n��V���UG�)RX�y��/*�Y����4#gR�����hT�|I��F��v���k�Q!�)6�[��~h~Q�Cւ�
�ߝ48�yT�ꐀ��������2D��U��':J�YX�.�y���*bF�����k�9(�����t����k�o���tf��Լe�)��`�LR&):v� �L��d��b~h���d;���ak��9���*�P��ㆾ?G(Dq�ZQ��ʎy�*��t���Z_j�fx�������}��"!+��Gc�Wķ je��,�ݚ�����Y_�ݧu8M��9�Vڦ k@�_��� ��UCb���y^�e�ǀ]��`�7�pD��*���8;��t:�qb�$�A��~F�P�u�W��}��]`u���|��ː�_�*`M�9��i��=[���m���L>VpS��f�u"�f���k��R����:�������G��t��޷Ϟ={g�i�\
D�w���c���w���<�%�^�]g@c���;o�����4�h��$�"��ޔ�^!a7���=L�b��2��D�"���~��9#��k�&���"�-=
��@u���2��!#fW��q����u\_|g�Q���I1�j|�e�a��[^U/�ee���F�ga�����Y*��/�$��0UO����x_��0����l�i^Y�/�khj���W�G�L�`�qG\>���kE{�Rl&�r"�;�\�U�RCVb�{	�s�L�M��%���u����"���.B�w��"�������y�Q'ü�A���GE�����h��:h7�ǫ�јȋM,*�
�ĊM�.R׋��M�L�b���q�M��k��o����}V��$��WU�6ѯ���(������-��c��t��M8{��g�����r8�G4� ���kb{�<��$b��X��K��^���:���7������M�|Oe.l�D��]��g>Ј���ט�W���0ב#���J Dx�O�������T����kk���pl��7!�'oI��X�G ��3���}'pJ��,��GM̲�I�[��1����RD��0�v��S�%8SaS���N��A���4��/,O�n.ν�P=���7����A���G��K\���^x��ͺ8ԋo��1�;�Vq�ZEeke����B��B;���C�V����R�Y���s�*#�0'�_�n"NK4�6	^}s~����X�>��?۰�%�}]~L�V����d��:��f[��P����(�;�D<���P��Ŝzu�.��_C���_�4A��b���*�O7�˓��U�:~�n�h�n��_�4��({K�i���~�~9}��-Z� ���o$��А;�u��:L=R-Dg��RpŹ����_8O���$�gk~�=K�B=� �{W���}3���xn"i��^�r��i`60~�ґ�D��,����_�y
����tb
�x���	�H��;�4��&�}/��]�c�?��g4�nG�p���+E.H��Q���̣8��Q�B����%~���5�V��	(�捇�5�<�8�A-���`��`��s���cI� `���O�%�Gh��\R��"��~��߄�a;����2���D��� )"�ՠ $Ժw�M]��������޽�TT�!��L�G=�"�Ev�p[��K������XDS9�*<J����r����mM��!~��Ȅ\E���qt�	����<-�F��#Q7����]�%�/;�v����Jã�VߔOφ�u�Iء�Cd���5��;��t���\�m`5�j��P �_�=q_kZ�RW�V�l�(�Ny���x��:0���ܫ"���	6���w�����;�QBb��u�*g���Pp��b�[�L-ʼc,��w�̱)�g��a�d�Ą��fD���v�5i��@c�s�`�#*�������G?���m9$'NЌ����K��%�<��>5"�����h��s���AM�6��
�U�1�?x�I��T�t��@\���K��i֊��FhF����o�]�tZh�7���q��l{��~d;+�#*�z��:d��A�)\�$PP/T�=��حc�z�b�t�	q�yjs;%z�/{�_��YZ�h���H4-�)x�Z�԰��J_f�=V�����-�`�m�Q�5�h���?������˴�7X�9�G��x#C�ͷ�]?#�v�j��dsyh��1~5Y�rr�H�_�>�߻�*2^��4���C�J���?,���1����O��	�܍ܾ}�ε�u!��h��y�7�9��	s`�ښ�
|���N��NU�@nn[�U��U���F���[MfE���o:�,�R ��߿�o\63���D��mҷuo�F�?4L?{�A���W>k4Dn^�~hK��#�x���Vٹ`~d2�;�+6:�a,��o
�܂z��޽,ޟ�����N_S3��o�7������d���X�4��_�N�;��F8D��$����JI���ك�(9/;�O'�O�r�̦�k�+|۩{�ɖ} �q#�]��PG[�VZ�X\rn=9���U��c�a��`Q��6A9�~(���UE�fv�g�V�ʻ��Z�J�N	ފ�H��n�r�q���1��]��HL�-�&�p��e �K��Q��91s��Ĉy�'�XS�X����+䵞����WQ�0�s�#�ձ�����-��	E_�0��)r�������Q�MX1{�����������mJ?�] ��]��9oN�2;�e�ϯ�
�V�[Z4��S�)n���(�zة�g�ތp���qΥ����c�T�H�_��XuI������ց�r����߆�O�q�Qq� y�:�f��@�a�����.�T��:�2���t��z��ϴ��,>O/���הW����zl�-2��}�v9r��z�2Ƌ��֕w���ƽF�����2i���iDZ�׶���g��gk+�7��n��g5��WQZ@��j-s�Sc�o�S���}w�o�?��N���"�<� ���7)z/�_5B�{����
Wt�W�yת�#,��������v:�U�����yo����R�D��D��b� t~On��]�p�� JԩЖ�ؙ��N�Dm;s��ү���bF,����(5�&j�$w�-���R��|������#/񮰁2����Y�PJ����^Z)̟������ez(J@n�
�njw�rDcF�R)����U?���G*�-6��M!�<9����#	�;k��}�f�lk�ytu�GF32<����/Q3��o�$J5}7����b�t�����L��΅H�xk�L]?Tu�x��JϝU�H�]s�C�駽���Z	6G]ŗv;��j�k&�!y8���~z�c�V,��GN��W�@���V\�6 t����j)�����7�d��ع'?����e"%*�d.2�4/�Z��	��пa�ڧ?�6��
�>,��c�X��x^��SDۀ�������GОK?�O-�;����G�#_\z�++ػց���螾�����B��������j���@n��u����B���3Z�Y��]z;_g�MG�X�?�
/���Ǧ�TI��'F�;��iZu��f���A~�pl���o0!��*���რ�ʹ�=���Ѝ�: ړO��r���Hzk>�+/��9c~x�
)��HN�Q����}<����$G�qƈe��r��rx_�O��MF^��-�\��Nv��z��I�Ӟ�ҩ�������6�p�֫��an�Q��=���Js���F�� 8���e�28�Qڃ2V ʔ>jk�>�0�S߰���/��R-��y�#�Yk/��������k	��Y�J��Q+c~ܥ�P��Fׅ��x@rd�j�k�5�Z(X�����]�G��b}�ū�L����S߽oݑ�����GiJ�=��[���VC�LIK欇�c����\���"�����c��@zK-�]��VƧ�\Ծ�!|��g�������}�%Uc��bR&q�@�[O��Ym��~(�eb<��:�>� 8?���rzV��7ǆ�;����j\�|����g�݄)�����I�ٸ7Q��^1���SX��Cv����<��V�_a��Wn5��]�`e)�*a�a:�7�
�Oߗ�>'�%�ٶ�Q���Q�2�� ���H�.i%X��gg�>^~he�W�e{�:_h��gk����}����OG��'�HdlO��D�M諾��_���,}��3lF`~6��|$�5�K�JHۼ�,�W���c�STI51�8AƇs���T�Zq�^�Y���#l�����L�l�8]�;���Z��?��ͱy�����s�]�����({fm����q��B�{�4c�b��!�Xgd��WJ����~E'�滚��Q
d���`�Я��c�NB,'� ��i@\76:��6Q4e�?.�L:�����h�A�h�gkj���M�˭�Ϊ����nP��yڍ@M5~R�u��"i�hV�w�Q��>I{�\z�� 2�/7뮿�w8�+I�0�R'��2�~�3�'���DC�D�s��4pVֺ��Y�zv�u�D�޽/�.s#l�q�U��A���7'B.���y�#\��Ay�
�>pEofW�}�Z�'$<#���!֤��l��:Mda� ��e%�����<b��Y��e�:&���L?�w �W|�?�Z�89ë�{`���l��[�&���2s�S�*/$H�մ��xUOtx�H�l��P����}N�;���[W�������/�˗¿��O�������>���������}�C��N�w����n����W���~]�'1wF(�Aև��x���Ϩ�Bi7���ϑXŏ�KȽ���%4`x�K��O�>���w�T���u'O��s�w�^���4
2TV"�����JH��F�n�*��8��kFJ�~<�����s��q��A��>�`z���Է��dE��ʘ�;p-5��ׁ���*�ⅶa���&f<�4�YW�Y����{z3�hF�`������l���-_0I-�S&����Z!�Y|���n�c =��f��<��ի�o|�&��\����V߱�U�e��k-R9��RxG�v�W�3T	On;k.�4��)wnJ���G:i�:$���s�G~6�p��v�>V�TAXn����*[��z���aH{��#�|Go�Wo�橅2��׽�:��	�{E�W�����S;�{&�i� �N�>��8��)^�݃O�����C��~��hs�U<�,����U'��7n���su���_��E�F{:7�i41��t�a���'�;72C��rKGU��O�4��Y�g��K�����G�ޛ��d�W1�����Bs<��|�w.o�T��e~ʈ����b!�-�f�'�7�^�'�tk��V9�RD��5�窅�|q+&x�&�:���BV�@ P���M������px�HlOAj�ٗ�U������968�/2�����T�f�+����Try-AL�"�B���y�f|�Q:GMS�m�G=����{���O�n]�! �!�D>���6�וy��r��H�鯧�s0$��*��s&�Wb��R\�IJ|�}�v4�cz��S�d=��,n}iq)�I����3�?�Z����S�K@.
��L��z���a>yeL���S���K�TaL^��$��{e�g�8��7�/�:ұ�л��vϠ�,�fҢ!�����Yݸp��cև�b��̒�]��'hyT�-��:���x�W��yzk��8g�Vw_J�i{�e'��mӊ_�w�-�m#�>\8΃^ƌFAש���u�~ �l��=ʮ� ���w����CT�ϖ��������5f���%�b���=��	S$�����}�X,��X9��+#|c2� (��>y��G*�7o�?���i>��ru���s��v�@��\×����t��Ȇ�Z�=�xq��rz��n�4����j��ro�3��S�6M�B��<��#�I��L����I9��?dyE8�lZ�Ƌ�4y������ͤ��~�i��<+��=�ݩG�����S�gs'31�mdG��Ġ%{tk�HEYϛ|{�"y+G��U��i��_����e"5TZ33�+��z��?���t08�n>�3?z+��P�m��4�d糣�j�;��[�Ҹ\������<�e�a��L�L�/C��,���`i#��ݛh�r�r4v� 'Y���Y
#B�yM������U��ܼ`�R��ׁ�ڠ�n��~z�\�^!�5�/�|`V�<[`	(.?�͌�@n��Uo�j� G%������
�g:��e�k�t����7�����Y^��Y��˛H>�o��pWT�����L���@��m�� c=�y��f����7�?ݟ��Rp���ߨM���)�빅؂�Ь
���O��� �
^���*	��zh&�o|��C�k�-�4���d�H^�i�w\���� \����-�7�S����pЅQ�e�Ќ���
@.�X���沰]�2N��~�T]y�џ���{U6����-f��)���#�^�W�ڑP
��0� vcP9H��_��5���i�2=a���)nׇ�{H�a�n?�{O��k">�O�����9H_�5�7�H~����HE�N.!�j���B.��9����ku�kaM�������4��fg��;Oh�cpu�>��w�����Ɠ=� /!���ȿUS���� ��m���{���93�w{.jaC�А����3�bf�m��9�o�|cN�׵���[�o�9�t�Vo����k=s�����"kC��
�ax�*�C����0�qs`Vs]���A�J�W���Θ�1���y�Ij}�ٔX��� �?��\��Q"�딡!���Kŧo�Z���ٓ
��F^XdGRg.�2C�}O2�����D�ۦ�8�%�n4�CB"��,.����U˱{��e�M����K�u�\Qs����(�s8�Z]7�����h��9A��IQ�^a��å�eǡ� �fҖ+��Mi��&쫠��.N�!��q��o+�j��@�KC�?T�d�*�����d(���v{Xs���"��#���N�Qo���i3�rP���ϒ�땵�\SnFx�?�D��#^�L��9+�m��=����kuMcT���ӟmi=������@F�o=_0#>c���{��֎K�砕��{�B��Bn�9�Uǋ�g�ˀ�{ˇ���Q��P�����/=���N"� �y���
m\�t�#�?�U�j˺��<���0؎���M�ՑT��ĈT8�Q8���jnN4�V�X69��D�#�-��^�!Pk��>㥏�Y���S�Ae�FkR&G��3�+��C '+o��O9E����9,����+z*��GE��p��*L}`�n�.��.;��ͯ�r��)�#w��Y�d&���Ŵ
b6����mƽ\�|]����C�{,&�E-�������Cb��RTNw������܀��.�زU�|�7o�# �S;ˀ|\d�	���I�ߜz�-4�0��y�^kO�t��-F�)(�~}��Q%������`��F�>��	�`�L��F9kSX�R<��~Mc1�M>[/�R�l��NL�1l��tD�Qa����l��h�{�E0���&�a�7U¤#���_r�}����F�Z�ǚc(�K,^�.�Ut15�rK�����u�,����.b����;{n�����V�V4�rLM�Y�E�߼v�t���w)Z{Js����r$o'�в�j�\F�4�L�ZRנ�,�<�g�s�r�"��Hъ��N[���*�T��8��m6��m��*4���5=�C[$C�����
��`���)ju���x^�f�w~�����#���[�
�[�[늜�Ó�gj�ꦹtM�(Ukl���2�5%���"���`H�c��� ��Lt���B#'�ۼ����Ć޻C�FnC�63��Y��,�|Y-͝A��ڲ�.���sW����&%~�,�.���=n���t���3��g�},O`u��)=�u �����h��鮁���\����t3�&���$���eq��NLs��>|)�*�/@�LT��z�+����zO�:�*ɸ�� ��-�c��q�����3���)x��}3��zΰmM�)sL��@��:�$��s�k>�]WoŔ+c�?�ֹ��#��l�_�mc�cF�$r�v$�������K��Ň�����3�cf���_�B7�*F��Oz�T�aUO�l\:%�"{[��*�<�͂@���t(�W.`��C���"�n�=�����V��UC;c������Õ8�i*vb2�@�C7sZ��\�wt����\Y���8AI�n�����e9jQ�u���ǯ��gh�v�q֎����0�׎��8���JƆ�V&�	�:���]�������hׂ��v�;�ΫSA?�O?� ��Kj4�UA�_�(\?�ko���G���֏�SA_�a�n��U�&Q!��"�������A
���;�P�LfvǊ.�j5�^�29�����"'�0�^	��3�ۦ�"͌��
����z��'7�cnP�\�*��-M|e6wvn�['���o6�}��64��wgk�d�L��m��r/�.�� �d����t#D.�s�@�w�n.��M*^��I�^Z�%���E,�pz��Yv�*������88K��B��k�����x���=�o���C(�"���=	R��ܯ ߛ�A�G�_0p;�9�xNz�t����l<���׉t������B�ـ�w��9�Eξ��^?��ön��A篱����YZ�Z}�ZW|B?>aԥ���Y�er_$�n(��Gu�<c���;�=�q��\8��l8��?6*蛕�x�d�;m.t{(���淡R'�#���Rc�����-��}��+K�t&�E���=�9�@�Z��N�h��f�M�̪ޮJ���{���sˀ!F�Muu7]�8�!���C,�+�m-j(E~����+��9�	8{a �?�߈5�����Mo=>B=��^�&9&o-㍐o�h��v��mTW�[!�Y��J��Z�S�И�-S�z�zM}"�mGA�"��S�|�U0��`�'�V`*R�&Y�ZTZ�ʶ�Ki����,G$ZG�ϔk���1������X`�;���	<g�<�u�U������.��Ž�>��Zt.Í~���v���^�����fg=9
nwe�ʖy<�wo}Ѿ���uW�W��l*�S�*0�����z��@���L�tH�p�}�V%��䩍z���0�z�D��]�W�86 N� ,�T��(�?�� ��Dz*II��c����`�#Y���
(�de���(��8�U#+]�L���K��)���B]��BTZ����l�E������L�]9��^�r�wޙ����'j��c��v?��$Uf��N�#)u˟rBt��XX	�j�0����c!���&�R�\��F�9�sb����b�P�W>�Cf��tF�� ��A~�tL� �
�lS[�Y%��3�bN?Wvߢ���1O��#�����+�S��Ϯ�E?��N�^����5�Cy���i����H�Q���\�M�(ejϸ��X.-�qЃ�L5��~����a����n(�[��]��H�;�7���+�0��_�����Ë�����b���$ yIN�0]v����_��R����RC�z���	�U�l��G8eF#I��g��_%ꋮYD�Lʽ�]�Τ�|O�	5֯5ddf����Ȁ�G�-��l��Vl�BM���]}�r<<��)�<�Ϻ��Z�\�_�H9Ʒ�~��=_ëk��P����oBd�[+R=�@	��_)��#,�҃������c�\7�;͇Z�%�<ZRa>D���\�(�)KI�8�8S���>��U�h�(�s�ޛ�?a�5���W	�cD�U-<}c��Fm䤑�jv~8��L/�%?T|���tQ�s��E-�S�`8��\g�s5<8��;��O�-�1����ޥ;F�Y�dȠ,s�p.+>B�]}�f�S�nY�=�ߡ���3���=�n�������W��������v���+��?Gl%�_K�fy������nZzRW[qW󮪕�����O�;7^ap�Ɔ�Ez+�9ܱ�̋Pm���b5�:5�h�lV�Mj���� ��~��7]�DE����_Ҭx�Fm��3��6���8f��z�`����.2+c��n�_e�h����X:=q<K|��f���B^��y�	'G�	��e2k"�j�~�7��ȉ�&��}ސ	!�2��|fw}u#:��K�^b��`t��2~��X��0�m��5�$��f�#׍wF�6X2_)�)��5��ݒnBx�ԅ���"���rZ&g> ן\���[�]���@\�xZ!iˬ�4կԨY2_��,7�e��tn�N�_&;+�T?�l-��g��Lu�Gމ¨���r9���{���#1K�g� �W���U?�Ẋ�x���N�Ɨ��2Y��'�����̇�����e����r��
�l�aX�����"�@�N(9o�
徇��Q�$�^�V�Y7��j���9���6�녏65 r'҉@�lqő�l�i���=���zM�r�)���u�Hި�޿q��&LS�'��%�t�c�b�H6��U��%!b6c���$�A���������#�n"4o���h
�s�����C�ǣ
�A�V�-}��)ꚰ;3r����T�p�t�oO���!{����b�{MH4�g��}�iE:<��n��Bz��f�G��[���<�c�<"���L�Ƀ��._1ug�%|h� �7���,���V��
sGc�5���D�W�MW3�KY4��ϊ�ω�/��5DU���i�	�x�R�~�El�A���X�K v�ݡ��\c64�J��#BϪɻ�͑�[�a�9gS�Y�j�5'�_i��%T�j_0����;���]�|	\�F��1m`<<Q��>#lA��/s��M��w��D�U��'܂�݌{ɳ������3�ue���?B�`r�=��(�,��M�N}���m��E�vr�39�[`�鋿��iX�(xb&�۴9t��ʃ�dZY9HT)7�Fd�D�	^~h��^�2O�Y�W"7�P�=�x���CP�h30U�1���D! A��x��&���D�VPsmAq�!\��9YG�: ���J3M2���]�γ<ZwZ����Q�a6LG]�����j�^F��{��W��g11T)i�B�Zu&x�������k+��B�$��✧v%n�q�+�Ag���}�}kh�J�޹l���eMb�<ڀ�gp���{0�7�p�!Xۏ��u��y��@�az?�/&t�	�R�zS3G���@�`��8f\��BAVs��=w�lDk)��=���b��!�[�	�.���:����B�!���g7BM�keLK��ʟ�.�Q
r����g�|.]�?����kJ�G4EX�J-�u�x;>����V�=�����ş�/�m�n��⧭_���jF�s����I��- �%��Z�a$}x"�$>DB+c%��
5�b�<����9<����Pɤ�.��{S�m<Y���OP��8Q�}�g�"?Ν���8�鰤�"�W�.B���R>��A��2uo��q�aU�:�~�=�O�_c�F.�;?R����(�e*�l��cmַ6'��aA���]s�5��ܴc�&���[��r�����9����]N�`���|�ʍ>v�BM{CE���Hu_�D��q+Vw���(��^e��l`'^�&�Ά�/�E�s�F�]Ѽ�ӽe;�b�9$��x�m�>�8�D�`�U�ɩ%�Π����\��|��\���{_�ap�,����W�p�������jf���U�{@�_�R�S��2��$��Ֆ��L�Ƣ�)R)(iDDh.�hN��(%�ru�Uͣ�<�/N����\���8o|��gHjv�:�.���� F�$��k�L�
�g!]���h��Gp}��li�f���B�{@�ً{�%7|K�Wn��q�=�\�k����w��Pc]��j? ���q4�V��r��CGZe�f]l��۾�[/��a��|O��k1?Iނ//�9�%��#��wF"��Y���ތ�\��d6#2~
�}������E��������ɑ��9���緹H�W^!�Q�#F��Y�ȧ���>Sy��×hW��c�s��&�8�iG���B���K�����a���$���e�֬zA	7�%q<E��-��������e��e��5�yg�F���gp���ƽo���:�l�d�������ׂ�+�1�z��2&�#^edMU��98<$!X������k
��%�@����!���*��ʎ��5� �M ��[�m�e?^���w=R�c���u�R�gt��
c�b{K9;Xy�%�[�:����33Ӥ�S���]]D��Ybj��Ůl눨gm,��~��:ɟ?�q洟��<h��|��W��|��lb�6 �Y�������=����F�D�� �DV��K�ؘ�
�F��/֒$�" -v��L;ԡ0f�L>8����72v�]�~+N��"L;���T�&YF�O?z�;��$s{ׂ�1c�9?\��|��e������fi)�������������������da?(���m<��ss֤ab��5;�X�׉�MBj�MoTj����q�w	�ZJ�V"�sS	ѧq�9L�E8����;@�U�A�k.���Ry�֚�A�6��
��w����.���Ը��\�k�.a�E>��?��c�-EBi׻�����ݳ�g8��'*��&�=�cv]�<T�h�E���:Ts�ϗt����U�ܷɶΚ��Lrʎ8�Km���S���G�[�E�F4R�t#�R"�t�t7��-%�C���PCJ�0H� g�����ι�����yb�{��^���tY�?�[7�'-W�lK��d;߾U�od����N8�����5#�������0k�߾k�D2�=:�-��@�\�ݧ%������z2����4X����{}��x���=�O���
�^��ē�����T���OL:tk������_��ȋb�?��Jz��� �v�� ֐���xݙkC�(!v��0�;8qu��7���ۍf_C�s=6s]����6�۵��%�@OFe����m��A|2Y��\�`�����k�����q�?�j��/0�:�y �������d5F�1^�*��%���r>��>�ڴ m�i[]�~'P���}1����o�8t��ʘXݖ�}�
���w�.�̌�y��X��>�nB�>y�k����
���il4Q�ܮc��]�@)�b�Ob.UOr�~}#-�Zn��9����LFd1�G|����� �X�L0�	�<d���5{���V���0��,���,�]+D-�\u4>墢�;�^}Z��`�K����~,�SA��f2{K_���$��X��J:���l�֓�o�N�(F8��8^�_P6W�C`�ZeF��9o�&򮁤mз[���jKX߉R �)����FJu�M�6<{E���N�<G'����Jͤ|r��X�KI�����ĺ�����bd\���GOǔ`9�f!8�^���2�S�-�n�0��(4�:���v%3A�ͯ��XL9x��N���f@|��T6B�?�����a7ɐ�}{�� �������|ƺYz�K�W�ND�;�c�s��eQ�k�g*��o:��44V**[��^a?^�`�W��f����F�l����d���,��θ�o�y5un^�Rw�f�k�1����5��ix�������q�E�\�G���
����@��s�0G���*�H�4!!�,i��i-�1P�R{t�����Qv�M�6Z�s�@�%���,봲�W�#x�g���Wt��J�'�A�`(es��M��<��>��\?��[�ݢW8z���Z�����xc�%�7*���ʨ^�Yz��KGa��5L�G��T������O�,
�'2X�'J�|~�a��k�p���^��"E��R��Lz�d.� ����c�䢸q1ԊA���h]�?~���-�5w�̩��N�v.@��2_݃� Z_��`K�������@Q��I�}�:t�/f}�f�,�h"�.�c`��k�n����V�LF}{���MȱJPUE'�Yܶ�Y�QDe'��ͧu�@�8Y����5OE�ZjfyuY��`r�����}��a0p�r/y��Ɣ3L��?�T�p�XʤH�m7������o�?q�o�������cb A�Z�Z5T7	L�(auB%�2ջ�q�E	����%.�:Q�1j���K��tJ
���qh�ֈo�/���+�$�}�����W���I`��a�M�g��:G-�%�O?=�]:R��?�jE-<�r��4�����u�r��J�'�	��7��]���)����(;R�o��Q���.�w�]��c����u���*E�߉0������L�U~�j�tg�{����j''���Tœ3}��@#�Gph�e{v�[_챛�@�����N�a��~�Y�Qt�ܙ�?�N�����*���@�$,�]+��J:�������sԫ��'�R�����o~a\.�Û��� 1ɠ����C9� ��b�3f�!�~�L�?��˖rny�1<˖�N��N��@'�]v�	��bB��5�n!�̶�Ȧ/��a� ���de��vbk��Jz����x\.y������vPPr�̆W�7:�)դ�	���NJ~u�j)�HY��0B'���_l�������7|=������^�Vk������B|�x�Qmt���K�A���uf�{3>Ѥ��7<2���x��妓u�������f��>�K`�,G��x�P�\��\2��8��]s��Pב�$�I5J@s��ܲ.{�
mlN����ʐ:�EW(�&����$�A��JG/�&lxF��
ΠCZ-Er�.��H��]�0�ELӴ(Є0'7\��Պ�{;� ��$ԋ˫0���4嗝�vla�q��p��ּxw�ծ������peP핋-d�	���ב��CCV���礽9k�k�fK�{	|4�>���nς�?��0ґ5��Z�$�:A�`���?Y��Ș���6��V��G��#O�ƾ6������\�y��>�8�d4���4�"A0:�,��u�����cLm=˝�.�Hs�E����1.� �8�3��B�U�c�B��?d9fܙ��P��C	K��Vմ9�	�n��b�Q/��bu9{u�$�q�E��κM/l�%�昑���8L�q#S^�?
!$�m0K��ɿ��$a}�j3�]��	�
,�>B�J����:Y� iwUS �t�Z�u[�-���S�Y#�~�!;/�z���.�eI�4(l��G�;�>�W�����4�[}	n}�;%��O$}h�f���v=�F_�o��"��o��3��.��,�K�lW}�J����_# ��nQ�83	3�����":io;�d�,Ҍ�c?� K��	?Uޘ�)�����w����5o �dh���Ϙ�ZA/�r.M����f������a�KQaݟ���U&�V�0�����ʠ�^�t�-Q���Z�bnk��4�w��OI���$n���]s/T�l�ۦ���>^eP�K�_Dyn���rD���.�˴�G���ݭ��?�!b!馎���x�k�'G9�䚚b}k6f�r�
&;.R
�����z7�oyӗ�~k0Gs����@����B��>R���)�OJZ9�їw�"�"�m�g�s��?���p����|B�T�j�Uo��?�R&m��'o>��0\��a�R@F��t�c�==�L]>Se���f��?9<a�+&dV�ҬTE��A����'�>�iĶd-o͌=
�㫖���~��v�b��c�;ݨ��ʹ��k4S����*v�9�J�;���3g�]�f�<'s	�5�2���V��CM��S3�Yj�6��:;�S��y�B��c/��n��l�ڶ/��g���#'�}���Oz��GdG�y���^��C�pw$��!����-	�݅�,���+A�=�񲯮>`�uR����ol����0����*��� c��?nӲl���oKs?ƨ'�A�N\�y�N�楯��ڢ?K8\�/������\ν�a'���p��D���c��
�t"��������DD�CW����_f�V䊠�7�ɻ��yGu&���/࢛�v���ڐw�B��Dǡ�r\!�.�S�;�8U11�'�Qn������1�ڴ���������0��%�]���6��Y0tP����$�U1v�/�|k�t�y���l��;_�����YaA�B�B�s������46�ިT�Ԗ�Kԩ5����;"�Q��4�ގ�	�����`�S{���\�Z(H_6kа��~]Y�޵T>�~�a�~���CLZĀ���ք�,f�K(
<[���[��}R.�9$ݔ:Ag(������"�]D�-E2����+��u���Q�DE#Q�T"�xզ�E��o�D������Լk^�\���ͧ�OO(�hnWpܢMtI��py�D��#����� 2I��T�?i���T)P3">���J���k��;� "�LfW982��/㧹
*�M�^	�j�!P.p�N�2k�gQ�˛ +C�}]�E�2z����=ȉ�w�Kr��U�e�8��4��4j^�#d�1�Zc,�=[���˻�����P�`�_$�Fo��N����Q>M�"�<�����1��?]U�M/<�H�M��[b�6��4���n�
�\b���L�5�����]�29�9�Z�O!����}�q�_�D���mn��{v����Q�W�Z�%��l\{ηд�s6w��5�,ۤ˖��4渭ʳ� ډ�]�c/J+u�� �h�	m��00���쎘E�b�xF�s��� R�#<J/h��_'�GN�e x<R��%�C���je�R�3o����;�B�Spe�׮�2�<xh�$�	ʡ��
r۴G��L�����z��uJu4a]v�Êv&i�[�$�wL�2'%'ۮr$e\����ٱ�0$百�V��>��˼�0��tZ��3�����~w�f�s�L� R�7�%`���-�Kv�O�8��8J8�/ũ<Z������U��>�;*������U�����<�ϱ�������{ٿC\�Ez;�}�t�J�M��<�$�²��< ft�����Q�F�o$�W��BF��Ve�ҝᬡA�y^�^S�y3Q�rc�Y��g���$2+�������:��5��@�NL�[�Cg��<�[��ˌ��(=�r���E��iM��{^��A���aw9�^���㩇C�����?l�"��I�,�p_yP�k�λ2V�{�m,��G���G�Y��Ῑ���w��X��ʄn��*m���\�����G��\��7zխ�5���f�����vӫ���b���m�
����Hx��}W$w�:0�=��q�'��/P�n�F}����57�Tn����c������^M��>]^��l�c��9j��e�/@%Jhr�$�Qm�=�8�ۙ�}w� 29m$ rKE��a~�W��8��Y'㵜��h�����_6�T�K�!^rr�(sQ��|o'm�[y�o�۾3�䒗�&>oG9M(*҂����9;��v\:��E��p�߇uOo��,�i��X!&}m�~W��y"��+�����@�9G֥۝����8`D�_���h���5�+*bp����䒕��܁⺘μ�hUt|q�r5PV�'19X�7b�FA����:|3נ�l�l{�D�&
�JD�Zw2QW�:ѫ�����L��̿�a�8|k��g��������H_����oQ��W�Wm\�r��UP��hCC�/�T 'P�y�7�}�ϲ�CN�-	U�Z�`�V����l���t���M���L-k~�v�5b��B�(���=+�z`��|+I��[��rB�r��.y�_�#u�֒a\��r����ǠJ��c|�z��X2����r�^�nsړ\����Z��/��fɵ{�{Q6300�B�:�z�y4_�=vZ�����ߧ�꺃�_���,��ʹ	��.�JJI��� ����4I������u�r:JY��{;�
/�=����x����A�����"��؟y��s�u?F��u�ݘP�������a����aׅ�����d�`U�?~�SDh`pW\��z�D��_���S']������s�J�5���Fw⺸�����&,�]d�W�E����=��	�㤖����hs����vlҸB�o�Y�V��޳���C�!�H�������=��� ���6��f+�z�K��ӄ�L��}>p��d�sU��+�0h�����gڳ�`��@�_��X����"~������eVx8�(���v�ɏP�|?m&��7�pB�ɬD���q ��T�hXN|�MZ��oo�{S�I-0�uf��YhtNt�
�5͂f�|�������輟
�=���v��[�:�)�j��ï_"e~wX� ��q�S�z������2��i�)�8�R-K@�㰔�3�����@h�ڸ���{Rb�w~/�.m��J���b�t���8&֔��e�T$S��X��a,������1������ِ��b#UZ�	�o������PW��!mkxM���(�i#�9�V6�T�+B����o�ւ:)d
 ��q2�CFʾR��u����.��zy�?�`�{ĴN�<��p�3?6	zȎ�d���0U��,"�wzF�����fL�e4L��	������0��hz���k�'�pL�䒍,�M_!�Pb�)� �i��y�J��5�%�ȐJ�p��=_��f�)�s�ƹ�^r�顷R�A������6�`���',�>���
�ol�������Uh_���Ю��G��>��-��I�����u�zS���Y����l�r�U�*Iq�ݲML%<��b|:O^f���0��	�O
�W�?����]G}�5���|ׇg�%�9�^_�z�+�(�a�8_��t�����捐�u�R�Ǩ�_�dha�=CDK�I�zƣֹ������ƻ��x����{�Gc!���i��]L��B��<���d��2q����ɰ*3��ܛ��7��{Z̈t��pp�@Mhe��z�6p,b>��tb
������H¶�K��L��qo�;M?�l�QP���!�뛣g�x�d����S\�q���t��K����V��'��q�ƫ��ٴ�SS��VM�`d@�UY?\P��K4���llHo�Ã/'�	z5����SyZY�'Rƿ�n��X�:�m�_o��M���
���'�21����۲̧q}�P��g`,�Ź�&���ȚT��Π�|��Pz��"}�~"S�.a���<z8�2,��z���y�D�7�|�������W��<佰s�g� ڧghJH>-�����7D���G�{����*Mzߌ��Rj߀3x�)bbT�Ҥ�?<Vpc���bn	�o}s�S�~�By����5�>w���N�� ��V'u�y3]_w"��S�{v\m��}���W��|�8���v��V0���$��V诂�6��nӧu�|�TzR���+���þ��3`��X�\�][Suw�°�u�*b��$� ��j���&4[e&!)1�iw�FAK��2�@ݟ������WY�
����Q#��`��
���o�ȑ���"V�֬b��f�h��3���jp�oNbl2���P��f�Hd}���9,���X~�VH�vQ�*�p��dI�[�14�E�
\|���̀A^�~$b
]F��9�ӄ��;:�z�{$�Z������/�>�%��f�~T�v�.pk�s����������;Ru�t��� �H�D
r��bM�'`�X���j�a�b3�H�������H`�Ԁ�f֛�]�m�'AG�	�ܪƎ;R\��&8��	mK�"dR�}�Fi�9��l��9hhY����x��$����eصgȸ���ֲH7z�Y %)���/���2��MV_��4.�1IR�n��݇��c���r�1a��T|z�b���?����e�p�b��8p��dƙ��~%u�J�d{�^~M�\��i�[�O�X����&Mc��݆���s��6�̀��Z��;��[�	_|�����k-W��J{7�ـ=z�v/F�c
xb6��÷՝9,?��螞�i���,ͅ��f@>HI�{��QA�����#8�q�˾�A�v^�����X"����V�^�;|��J��Y���������R%ܕ_����]�m�I[���X��{t��W3���4�����;:�k�}�m��޵W^~��~B�6��CT�^�݄A
p��`ߵ�;m�(�Ҿ� �|�����.� ��Tll�k��w����0I�!d�;!raY�`/ }��  +p �qv/Q�U����������a;�4�J?Z�P|��w��Z��h��7wZ�D�EVj�^���7�XW��PE2��	�.�+��5��E��n�s�l���z�f��w���gX��X._،��*�gy��������x��i�
�N�q�}4V>�L��àlM�T^�ӓ,=S���&a7i�U4k�O}�sF�qi:Ŗ>w@G4��`ߧ����&s�g�����
@����
�G�v�4o�dᇮ�$� )H��5-t�>�{@_`��ECG\�w��z|�.kR�2���!B2�}�S��c��T�V͈@G���ܹ�3P���"�^�E)^r��h�5�h�^���`�n*kq���D�)�x�^���rS��i���^DH�DLN>��՛Q{�6،������'Å��w߁��~�/���=��pP*K`\��Ԏ��G�=h���Sy���s}�ۆX���߂Ƚ"J�#�ڗ(�P�_u��c�@ᵼWW�G	�_�z������%����;B�%8��q	�&�Q���E�`i;=妣ثgA7�����yW%��!Y��ll��Yog�5�Z��.�A�]��u���8<��Dt����;����/��O(�;~�ߦ�&H9>��q�2h�>S�vw�{����j`�Ɉ2�e��h�8.un=
/��b�dG7��I�74E#E��o�5�GTh��h��w�g��'mxZ)�:�o-�V�d���_����ktV}��e{Q�U�Ȓ�mcB��[�AS�q'M�}���43,Q���"S@C/��C��C1	�ɴ��E�KZU��h�["ģ�����ؙ��h���G=Qb�l�VkWD�/C��S�Zj����DN��:�.^'rB�dGr�PVEq"審c�fج�(a9[_����4U ����I�L�`�ک�`�'_B���oEr���V4@��[�Bl�E�����k�x
�g՘njq��U5�lA�s1��J>������I��˶f���f��`i��p�=��os��r����ٚ�B��שY���Kݏ�J/n��%��O�cn����*�VG�̍o������q&~�N^��k���L����љ�=�4bђ�~q^l���1~цu�1w,!�c H�R	A��)X�AYƽf_��ċU�(ϼ����^A�{JH�.k��m��N�:��ʀ�q�{����s�G�~�ڻ@�lĮB+0��l����ez��K�����B�&�Gq���Uf��"���e��'��q��d����.TQ�\Dg�a�b澎�n�2�����e����ww��e%��f۵+-^a����c{z��ʷ��+�M�9Fbjw�[pNkp����
�z"�K2��W�1׻����������j��L[o����.?�}D��flBi����F(P����oh-,�,�� ���\l6eY �'��$�3"�����E]h�bt��ʊu���O�l�Q��H��u�_{����gR���mc�:lH�7�RQ}�5{�^Ɵ�
z��o'�|��T��9Z�L��V5D��6�����U1��J���mp�Ủ�v��Qi��ŧ�� 7�ҷ5�z�����M�����MN���"�/��A�)?g9Or�v7U_z~��ށ�L~ɼE��A M1v:ϑ-��T	k�����T��r���+�,5;��@�"���:�>ͺeޘi�\�����ǵ�$k��a0�;�	]y_�Ch�/󸧵�>������������0��k]�O�l�Q
�i^H��;�ߒN�
5U��V*�kt+y�	�����Ч�쐍<ӗ�|ԁ,ݖ7�0�j��e:�hy�
G�޲w�VUݕ�Pq����h���2.A��Q�d\-�H	�%�s5.��� �~� �<n�˾Z&�> >7�<#JU��+�3��R�!BЮ�$8V1����<+���;����fx][����d�[�|q�YK+�	�c� 2�wNu��il��E��N[k����8��v�7��L1���tc���2*h:��UR�W�O�lg��h"2h�D�G�3WT!�w&����M��iV�2Y��'�g<��dNa�T��˦��-6������b���]X�<�s��o����HT?t�k�\�S\�x6Et�;N�����W���록ڪ�^c$޻.��BvG�W�Sk���r��ݔ��Enx<^W.��y�3o�H3�<SL������ -�h�0�ΐz�/�GU���?��lx��1�Vf.ϥЙD]E�O�J��ܵۓ̞��˄�f�������%����o���Z{�W�;�h!���d�[�����z�Z;�#	l7T���D�	���y�H .�:�L��}V804aܡ�Νe��x�mI��ӼꉙI��,����s�O�s/�FS�q��T �G�&(���Zs?��l��Vv�g=M��|(��b+.@r�S��ۣ�����`B0_.n#4��{;��޻�tB�����&�nwg�t�X3YZ!��=m4Ua m�ҁ,��ơ�)sQ	�5;IG�	8��1:�������m��޾��HcȬ'0�[Y\ޏ�����˗�T�q�����Q3��=f�5n��� O���ӟ~������A1<���+B/騒�빉�2b*z� �YQյK�@_��$���K)��`�p�_���;�>~����(\'���ZF��;Cq���|w��)ۗV�l���e��s]���M�o�,h�� 1�$�v��2`[Y�s�l���JMx�"�?��f�s��D��b"gsN%�=N���{pۻ_�-Ww��N��"�kH�Lcd�T�-�W�Æy��O�Z�P�."�9��1��,6~��߽`�h h%t�WWk	Ri�t������0K��4�
�caҒ[#\��s?������nς<0���@�ѲBKX�҂)
���Ѩ�bPM����U�b�3�������x�I�:g�g1��c38H�> �o����]O�����tzY��FˊT����?rM�)���ڭ�4��:r�u������!ͮ����g�~NB��c�wrE���^?y�,Ӄ��.o����#���y�Q��� m��hG?�Y�7�� H��ddy�x@���DX_kB�+�i��Ջ���&�*���C�sD���ז��o<��Z*�ڳ�O>D��[�%�)� %��'��?$W�CFK���n�_�]$���8����G�R�1϶{-�lxkm  y�}6�8e��Utc2"��ٗYC�da�yGs���@�ɋ������t�m����s`��ho����6�k�^u�r%�յ~G�@���vIO�ygo���9�IA?��)+T�{�l�mt��b�B�B߹ +"�t�:�[�Lm7��07��[�f���i��揭�Y��"z(B�O'�~�
�#H:�G;��n��ȸ:�@팡�m���K�;6�+�nS��w���6�!�6���n��q'���/Տ���lS1)��jߧ��qC�Y�mGd�O7ҥe�� E��T۾}/�tm,�W�I���x�.7L���
��<��v�B����^�~�ׯ�ᨚԌeh����W����x�ygՏ�'���!�5;sf���|x���N�~�wy>T�(Ty���v��{6��c�'�����P��jJ�T�������_�n��x+5苑GL���$W�I�����Q�ˇ�KG��D����l��LtO�<t�Qgw{�1�}���<���*�_��8�+G���%yL[����B������_�Ť�9Q������,�1Ş�b�
(F�J���e����l�<m�ņ!&Я���.v���no���qɆ�"ZQU$�t�D}#�Q��bk%p��n<�}���z۝@=�&�<��&Vc�_#�N�"G�^a8O����,[|g.�ӧ;M�JsZ����RpE���4�}��A ��$��(�%�or=�'�bA�v�/�'fӼÖ%6�m����.�yE�}U`�zT�����nPL(�s�Vf;<k�!�V�}Q�P<p��1�U��5V$�D�	?@��'l��|g��;MR �v�C���������^��smb�\�9��ؘ�������R�z΍��dC�c�c�E:)�h_���.iE��7R'-Wx6�c"	?p��A����#$* ��9��+�zLhKu��%���=C��Lj�)6�o0�ElnDgeS+��p��ZS���]�u���4����Q�Yb�������D=�)����HD��Y4�F�]�Kv4L�Es5�!����5���W�^	償��/l7�U7]�O]�u݄�b����P��3�4OK8�z`N
B�9���\�}&��	���&=�GX�T��%�͒&�J�A�A�N�:�В ��p��K��!��H=,�BmVʇ���Ӛ�ɚo�+
'\<�͆���r��͠�k�>�ם՛'$c}î���[kю6h��Y덄U�.�{�Ba&ӝ���C��@�q�����]�K�4�}��|C�@����<*��F`Op�;���ʕ� ˍK�nc;s�I̒d���*L��?�l���?Jw~�KF�h�ux�ұ�F�k�WFӀa|*=���YU�?�u�4b��ec�J���q���V����j�E\�r�i�|��3�ފ�j�i 0�Es��[�~z��r������P6��Y�,"�m���Ǫ�'�O���`V6#��6�t��O��4��{�s�*"�YCH�m/|�����U��o��'�s��ۚ�K(�F+]\3�}�.���q�Z�����0l_iӜ����Ϳ��;\_�R�?^Dj�C7�Xͣ����nΒ��D��� DS�l\p���h���r�W"�}���+�I#SGj�b��lP�A�7�1$H�] -ߺ8�:�Zŭ�� t�H��P:?Y`��_�����HJb�=�1���D�W��A9��RP9�&��-u#g2�Mι��U��mM�~ߑ;
�}�X5���{Qe:��}4f����d���Ǝ5�M�e6������OQvDn'�
�${�<�#�&m�ݘ��c��Û�q/{��v�$�}1�=΍>j[�IB6�p�#ls׊����/SJ<�ڨ��W�|r\iL���;��yN�`2qq�f�>+���ei\=�����~���ټ6iD#Z�D-]a9�I������^GsD;R.F�Yʼv���?7
��:i��c];9�#G�9[���%z3�v��	��^2�B����b�����@=�z-��X�>����*�7B�<���֩]������J�?mw���3�h�D�y���b�=���v������^ !j��C�LX����L�3h���e�
� �KD��C��EO�G��P��4؅�
�K��b�jr�V���mP��r�k����rG����U�+����ާF���Y����e3��LH߰�b��p׻*U��f��}�W�E�b�OI�!�vɴ�.�H��*��n	�
�[��DM�lv��ʾE��T�����3��.�j���	b��/G�Ѵ�U�����h��Fg�ſ���/V��p�@�7B���G��3�57�"C�ϜG���o
����>��k�Z(j�iw�ޯ� ��=$%�eXY����]���,�����O�}��_��B[��g��5xˋ��g<�/a?ٮ�����2B��6��L+����ԉ9���$�'���jzd���2�^�o��7�Hv�������PN8�2����O;�<_4�s���ˣ�^Y��fZh�oVO�>��~�}�Y؋3��m�r�c#�߾�g����C�G��5�nI0G�i!���<�[�>��O�e��~z��!��wŊ�Fzp�=|�.��#��@@&���:a�̦��/%��gg���R܇� ��2 ߧ:�����Y��>��[N��q�Q��xU���g��t� �-Gow���L(��j:@��r��ͺ��@X�#��%p�/ 'Wn%ߞ%�9�ڜH��:���$t��bZ/�Y"�~�Tsoi� N�Gzk�	�Sz��x۹,*n`N�R����9�����?7��<�"��dZ��W�ur���uj?���Ozu���Pgu�67�����X��#{M�����]�,H�����s����-�9ּe���_<��Km+f� ���\B���蘏Jy-�3�=o��m�n+<\xυț���x�L*ws�C&�E9����	�y6}�X����%��4޽G�D��fn�p2������II��k:'�nĔ,.q�ޅ�5�>��i0�W��\�i���C�St��g}K>���X--	�Kƍ�4�F�ϭ~�i�u�H��b��Đ���p���M<�d��(w��T�*���
������'�`펍?��b��g��K�g���u�ʹ�g��px�VD��4��sw8c>��E�ȏ��i/�_<˷�-*���oLL��Pn�5��������"&tJ(~��Z�&'��Y�)�
�5i�m�[ks���3A�����f����(��ͣ��O\����9������ˌ�D5dE"UC(U��o�K�'�/�3�;E�!���G�З@I�!`6%8�˟M{�j�?�~���yݯ}v*���|�P= �^BUAᲈ�jl����i��٠�pl��67���K9v�E�z��=�_s&��o�Hn+���*��0X������I_��9�Il<k���Z�+̣��r��*;��:��[D�yU]88G$Ҝ-�̟<v���|(e�t!�����k���h(и�3^��t�A��;�������3<tW�{1��_�-���3+���3"Í�v+�Qi}1W)fq�ԕ�jH������<4W�����X �Ho�����.���Y���|Ion����+�W���[�c�ǁ���o�n�vR��:Y�-&O- 8P�/^м�G�X�d}NT���1}�l����l�,�dC��X(%�w1oEI҇�^��R;�9��;K�)�d�3�Ox��y��o�\�u/�rO�ڌiDmk���RA�G�n�t�����>�>>_���lR��:�y��Jխ��0�&������ӟ�[��g��v�7��56�e�>W�'�;T��ƶڤ���;�:9����͑Թ��8[L}�#�p�ź2F��� ����6���y��N�������:Z��L���篐�kN�i���$օ�1�t~�^>|��J��y��B���JZ~;�7)���֯n�����k5��^�sx�"!�}���l�B��XM e�b���k�cB���%4��D������2����;݂	,{�b3����,oq����?,�<k�[`�2�Z�8��^�������Ô��0j@���o���nc�q}�i1|��&Bh��$�6��?���r������[S���P#�?!���%L�^=<��?3�^:t˒@�M;>)1�.}�,x�� ��(
ڂ�&��Bڲr$v3%x\���J�z>���l�Q8k!��i�8��Ѿ#0�S�ѿ�M4N;4�,�t�p�h�E�OuNpҢS�O���N����r#�v��nܿočS��!;~��
dJ����"Z���=�4!D�ż}�#���UN��M�T�(�^:��<�e]�JN�6���^ܑ�O[�n�4�L`�1�)��c1N�����BQ[K��:�E��l7�[�C�^��B�{�*/�\8�~u-��������S���v��k���3s��x��`ށN�ىb��1��J/\��I��E	�3�����K=b�y8�Y]����
�����T��?���U�����'࡯�A����ck��u����`�ں�af��C`o�lG�%�P +��@/�#L;mUol-S;�Ĝ��i4�8�&g���@��U�V"�=���,⛠oĎ�B� ��pʦ76콈͢0R����b�E�9���6�Lk�z����A��(��~F�ӓ��Zh�.�����wtr����%r!%#����4~�G%�d5OMe\�;���R9C�W~o�?�JqI�{�O�z��e� 9�}��'����	�<�m���p9e_x6�RM7�3|�5acR�ְۢgK�Y�ybAD�r� �t��Ϗ�Qf����L��@�����<H���ߧ�PM��j�V���9��@K��D$�n��'��ô�f�M��*D1�0u򜧶z�o�.L���b�	կ}m*~�ynw3�ͦ�?�%k���7mץ��cL�_��_��w]�:NT8��v&��-�^OaSA�ܢ�z�P����C��1��U¥�֊_�J� u�����Sq]��f����S�7 �죹�~�Oz����ʚ/&��R ��q?�η=��i��ᙅ�fZ"���Ltx���)�K�`)�D�Ɨ��WT�g�ç'7������}R��r,o�����8�p����%��{��R7�w=���Z�i����Fv�F�ِ�r�i0zU7�To|F��������s'��$�yi��O�������5x��T���[��f)��_�T>mn�[��6�%���x�IPɁ��^��F8OM�'�L/�#��B�����a����2��yk��x�|0��YKR;��a��S����GC��}.�@hp��:���G��A�g�w�_�0|f6>c��	ѯK�g\�.��K�d�I8[V��}q�����^���`m��B�f.4�}�Ƞ�E�s
�2�1~W��i�?k׀L�KC��7���`CLF���t����n�ͧ�mv�K�>��o�ړ ����q�l�Q��T�'�-^�����܊�D�m-6Q'�9��U��q�:�8�g3����l/��E�9M=�n����oL7���Z絽��"�Dt?Im?��d@ܷ�$�`�7�l�T%�p�q��sz����p���VmK-~��/u�uS�|��E9�����7N�ߏ��R�(�.__I~���{��Wߘ�r��h*uK�<K�y�d]E�P�Rf�z����U�X�9����1^�[�����H*'��{@�}�u�+��5+���?���[�z6.|��z�&��xA7ҍ ))�J�(�"  0�{�H�HIH3�����0:G���{�g����}�s>q�X����L_M�yq����}r����:���M�&������[O�I�!_����K`)j�s�^�?\�O3����g[��7��ۈ6b�zA�t��83vS�%&�F���>1O¥?�b��M*�UC��A�m�9ci��g�x��!7�-0(�PJ�UD��l}����l*A2{=w=E��B�s�����NQ�)�7���v�I�9>���<I�^�`��ՒX���d��"X�<%��>����u?�N
5�Z��ϵ��s�k[�A� *���2|�i�La����ݥz������TRÓ��9�kǎEpe��N#��z�oٗ���[�lH��<�7�|_�	�k�9�����'�%\�*V��"1�'��Ac,�"�3�Z,&�e�'3�K·ؐM3	�ɹ@ܕ��:����UU��O�w	C�I�\��Y�D���]�_��Za��A���g��Ox6��;q4擣W����Z\}�q�{^f��������C��\���FU��ـ�>[��!�x �F���&���0��V��(�]��I��7�*�x����\)��7v���GD�>N!��m���N(�5�R�_���8�5�G|j�C�x��k����!?�w��\bM�g����>u�lk�������B`�q�<�߃U��fwk~���<ÒZ�҆ X�`	׉H>���QE9�W�nٝ�R�7<�����u���ŗ�~=���,��^8���� ��w��g�+������������k�R������T|�X����<�/�K5*T��$n+��ҵy��
�<��Qʯ�����P��g�A��y�,izhH�����ߥ����<��"N�	�M6O^6yi��cb�թoQ��S,���M-�D�@&_�\QB�=�#n�x"�|�-O1�.3�ҫ!}���寫�(w0������'�T7��?��qw~�7��yy�m6�����l�֜�3%�绯BQ�����_&�q��9�O��`F���O�yk���~�n���^�֥��h�ˏ��E���A�B��7��kS{�Ò;�M�⑽?Szfw�{_��QK��voT�KGF�&����>��LU�ea�V���p�B�q�k�ڀ����2H�+Q�L���c�S:�P����_�$7���O�s��[����������������1���g�����wx;�Ko�i��D�itC�rꧽveI����{]���8[�t��q��wX�]c�\�%X��C|&,��VقƱ��q�U;�ٶX�J�U�=��i���.A�ϧ ������
��.j����ܤT�ڗ�[[ޙM\]y8ۮ��`v�]�ڦ�А�F��3~���8kD�:_���ɆЧ\?����;�*�beH9l�\�����6_=�|<~�ǭ[��MΆ���������2�$��l�z����5.%S�^|�_��c��9���#A���}���T}���5@� b���K�{�%ۏ�l�/T�-�G�5�L���4�����Rt�z\93���u�iz,��\h���M�Ie��C4\�)�򇋖S�ef�j��a��p!��L�L��L�o��йs��ᙇ��plI�@�͗3I�Hܛ�~��s$&�N�ߕr{�)�r5��Zb������*V�b����}"jA������﹞�h��ƕpO1kЫ�3� �#��ɹ��re=�!W�$O���:�3�v�xE��b�Ch��C��#�>�
J||!����Y
3E��gE�d�����x5�f�q�,�����3ĺι�c�\�-Ŕ��l��y����j��f�1,���y�Č���L��L�Z�7N�Aɝ N�����GTdt뗾I%�,gm���)�7Mf y��ܒB��KF��%p i�\���-,�x���-�����y�3��@���Ot��䌀�i�Hsm��7λ߃�v��ل�,	��7���"U:+�Xhvʈ�?ṗ�Uտ�����E��$��4s���_��Y:��7͆,�D:�9��6��]9���D3x$��[gUVBL}F:��<6��璯�������pK���Y~���E��s����4<bcA�܂���p
x�>���Lk�H�1�Y�I��[�mp`t�`��$�����M�M��Ֆi��<��e��ă�̛O�j1�J�#�ō[VK�"�&���Z���/
�
S��S($
����6�w" �*L���H�`࿷f
 i��NO�mi�0,軿/�ͭ`C�������o&̦<$�e�	�^"����o����7I�@��c����W��;<�������W�����.�e��L`jEN�=���қ-��~�ҹ��Jݖ*��"D��8?25�&Z�C��g}�ː�����?|ʳ��-�$����7'��ΦL���'���Y~**zJ�����, I�;��""�>,dl�ehu|�WHx+Q+�v���&ZTP`9{	�i4僦ܓ�.�<��N�"��Y�3%`)���h�y:4H2�̰��Q���=�Cs����7G��́���R9�͉���ʥ���6�O�S��1�l��d᭥<!�Ok�e,x�Q����}[���0g��m�k�%.o��?��z^k���:��ϻZ��핹�P�g�_&��p.���	F�|��Fqaǳ{&O���eX�z7�20��@�\B����߱,��H�܊֑��>eV�J��rdds�A��cSJ��Vȇ��ڹ�'��}nD���o���7C�{���Ɂ)M@� ��]̍Y\��<r�j)J�-P��5km8Q�|�>+����;�Zu"=�S��#w@��!�im^2�"�������� ����DǨ�&c�Up�줍����T����"�< �5�u��m�K���7�9#N�е���y�����U�މ����>�@����jH��H+�v����"6��nM�#U�6�r%[�iP���=� ����?��?ӥ��q�^owt���h^w�a^�=�/N��P���"�sjz���y�9΢��g��e�j���U�w`M�C�oƥ��z����I=^���Y����64\^v�sʖd�<�����\/�H�o|������?� m ay�a���υ����c������G�������D�͚CE@	�zֶ��]Q!SĲ+c,��b��o���ו8Xz-�9r}�ֲ��}�}����.C�q����z�g2؈3���yH��l�&�g5�m>9�D
�yG��Nk�S�2�mn�i����.��͒~&:��Zҽj�m�h:�$�\��B;.���B���me�����f�o�+%ռ�/b��:Cr)�JB�����j,�*@'�v
�.�;��a|tm����т�P�l��3�� ���r��81��0���u��k����*�6&��e����+Ÿm
5]{I˞�U���jW�,���<0��D5���X��-R��v<+�<��G�G�)լ�����i��:J��p��0�ļ����������j�Nw����q]��K!#i�X�c�_p���V�2��|�;������|�.�-|�u�=%hpt� ���C��ݐL�ŕ�7&%��r��,���l������C�|KY(h������ntV�Yʱ�vqW�0�uE��{��.��E�5�nr���O�j/l[@��'����|]��m��DD���z�c������XL�|���`$��o����+��}�A"B�hm:�k>�{M����ڦ:����=}��i2	��K�Q��d��2#�Y�0�9��.�U1F����7������`�q�A"&��x�kb�:�=��T�'(�	�ƀ<1Y>�؉�R��~��}���zqw��cO�׵�/V�E�ꇠI��dr1�<𧺯q�1�� �g2�J���x�sW�y(���g7*����w_�m��]��e֛���� ^����M�\��c,�6yf�X<p�λV�����Rb��n���ʢ$�[Ye� �x�w��	:U�s���3J��#��%d]3s�\�M뭭ؤ�|�|��M-���A��Z?��~�O���LP)7��i�]��my$�[}̛E��������o�����U�OV�Er��bٮ�erqV�6����/Y�J?��g�p���-o��)�'ڎ����޷S���66X�.�XU�i�<��74��8|d��[y0Ԉ�� �*�����i�ժۜ��:������$t>p���0��~�ߥ_�����q���`���z�q������G價�Ɛ���_�m�V�@n�:�8��D��F�C(A��a��@�d��!~���F?gi"F��,Z�r���{n���#U������ۥ��ۡ����P��D�w��	6j��L���G���/ʼ9L���>̪�m����7A��Q��G"��G�qb�R�٨�[��E�\NIh&���A2]xx�;k�H�Zo�����GN�*����G8'��N&Y�D�08��t��BNT2y�+�xv��h�53���QF�WVy 3��'+ڴeOq�^�ˌ�MS:HL=���$>�͕c�Ѻ{��[o=Jh����tS��6@=���P`�p���hߟ⧟��} ��e�Wq��F���͆Y��o�X�C�W-���}6�^]�#~mɻ���``�CD�!��Wjv�K~�ej�i����TiF�1+2�ÀUL��ѹq�j,Ft�F��ڽLr���
�q�s��3K[����T���O Ij4�}ߧ�%��Jq�^ڒk�$��kС\���L2�/5�:�j�z���(����>��i
��WܠK�WA� Ÿ�,�Y2�z�Y�r��.=ot�Gx���Vb��d �q� ������Rث�˰�G���[�8��ƖV���A���]Y��O0­�"B��+f�W�hsgN���q��{v���1FA�h����}�I�RQ�0���E/��&G|�?vk�����!�1}�hv�7�M�My	�f��Q ��}��4��,i
3e{�M�ryD�������P$s�Zr�Aѥf��4�����ܛǺx�M�Y�D�t;��\n���
Pg���%�%�řK5]|3�+��D`�>��*�W�nzbat�`����~���'�n��T�o�[�̍�^ל�u��:r"��א�Q��_�nلx������'A�y�AI�r��N���fZ���1�l������}����链g�f���f�̵^�^a"�|�za~��mn��i�������H��婷��X2�;"ř����z��P۝���
���~|ݭJ��Z1�ߧ_�_��xYm� o4_�p�Aͩ�3���9/1�r*�_��r7;��׆U�Wd�y�>�9o׃y�Cy��r�<�9���r�ą���N:%��㑅�e��^�*����՘�j������� ��"��˷�kB�X;� "�H_�\��up�︑YG7H�}ǖ��=(e���_��
MZ��R
�˴uBܴ�}�^�A�n&hJgM:�F�֬��;���.�.5��M�YC��W�Y���AZZ���$ѳ��אU{�O��>~�v�XƁ��U��A�d��,�}��a��˞�H�O�%y�ɗ��##�:���uũzO��s4R��؍m�V\x\��nMFZ5,C$�=���м��FQGŎ�3�C��~�T�/<Iw2�k#����� �2������6Fl{��@��>h-np��tݼ6�����8�c��b�B�N�_Џ�E*ȹ]|����u�4R����\n��U/���pa|P�!=� ����[UJ]��Z������Ƚk�'�
��n"'����	��k�QKֲL�����'#7����P��}�o<���%�=<'7�T���$�zK�����ɐ��h�S��h�2hs������_��<��#�v�j�9��37��ܗ�|T;��5l�#�7L	T���l"�Ȱ
«J7�:wk4�v�]�R�G��4�f�;�=��;���t��y5p�ΌI�ߐ�6I��C�	���ظ�ْ����\�e"�eNGp��b��M4�9��޸���/��-u��-b��U�\J�~#���[X���gݼ%�|s4)^u�x����<���;�֩� [d�9F���kj����Ca�-��&8ǐ�ڪ�)����em=��h=���c�C]'Y:��}E{�ܱ��}��A`1'���Y̱�:��$<Ƿ�D���n��ߞ����������|Fօ�Uw�D�B��˗�3-��D���9��<�|>w%ϠT���x��e)*�P����g���܌�-��)3�������B��/S��Ci�H���p[4m��~h�7�A�Pc�[��h�Ni��%I1,�ɤ8-*Z�N��28ˢ`��Ȼ<swi�!���r��R>k�@�3�!P�S�#Ҳ��X=�����Ij<#�\D��|�c�~��q`g�q�Ŝb��ߺ��U��a��K t�+��L &K1��29������{B��}ɂ�s�8�p/*�(�X�Жm�j�No�1�1i����QS��Z0.ٺԱ@�ᖶn~ݾ	x��`kǱkg}�faR.S����.��*�D�By3ο����E��E�)�|�Iw`~y���S�B��d;�`�0M]M���`�*t�Ŷ+�'X��X������"2��G��.��-?��
VB|�=��+S΋�Wpa~�'2��A2c�5G����%��PU�@^��wE��G��|��3X�j�أ���ۦ���]��Ph��TD�wơ���6�������Ec`~Vj�� �"��n�er��۝N�M:Z�4���E�!��,�r1F�KP��%�I'�|}��:����י�{lR��>#������ź�wg͝3�^3�Q�5�:$�]t�ֿ#��73˵͉�}
jݺ�@r�����ߦcĆ�"�\�[�<���岲T���.IZ}���#@Ĕ>���志.V�7�^l�uk�G[7F��!�;�7�d"=E|����VG*�>R�h��������ψ�w��z�����*rD�W�Ȩ.MuT��I�0~����� lؠuc��@%����"��%���S��'� �;�wR���0��L`�O�a�<�ɛ����_,�$�}�'��A ���z�
 d��4ZEZ�������8,���R��*=<9!�\�)�[�Yg
�#�ޫ x�?��qY�'����t��PJK R����bjK �0�*e���V�+��g�L�`�Hp�ok���HYkv?�	#��a6�[�"�3�I+�oXi��=v��۵{��6�C�X�WF>­�O��6�Leo��+�ƋI����{g�Ư?YY�u���x����O����B�O��H��_>�8|4����Td<���f���ʁ���Ȼ�B������u��2j�^��^g�c��X�"Q���p�?���:��)��n�,�tl�vc��)�����c̟��[��[H��+';=�>!����c�H����y�m�[3e��]�I�;��,x$����\�8��q8��W�w����{f��O0�r�O��pH ����,-�r)*,C_��D�8��a�a��Ѥ���w[9��7E��~ ��)��J��nT��l�6B��c�'=,�D�*����
� Ʒz���Q����W�
|<Ҹk�w��p=��3��oːƒ*��ץ�h~����5�4y��U0��<�
��\�L��g�߮�>Oe��j�k������`I��KN��*��fL�k����=� �_	��.�oj?�� r���"�~��|ǓȯG�!m^��J	��l��"_�9,�L�<:�)�m���[M�!�Dd	>�����N�k��ߺa󾐩k�����Ԧ�>F8�����S��ŋw�6���b+�p�DC���o`h��͓i��Ҝbd��?����ڇ�=='K
�����.|���*[I��!<�S�"+���ɦ4���r�`�p��s��=���z��?� iY���t�Dw{wYp/º=�O���:n����A�N.66�PUy��j�g�H���	���70)�ؗv����$��5�w �����..`L,�$[��]6�oÑv&��EAD��pVY��-��1�o��"&/��đ���A�xQ9�>�%��n9=3��\m�ݷj��_�{IT��/�|���Rw.�����&&��k].��5.7$oC���ǇJV]^%K���|�@u����6�>� �4�s��+�y`��K���c�G�Li9�FgXg�`��g�;UJ�{�8J�=:��Uj�dOX��"��L,�W�Fe�p�Ǯ�����.D����O�D} ¤&�5"#<�%/���g��6����������tl�G*���M��*y�i���8���5�D8X�Fc6�_)�'~�Y�L�ل(y7��"���S��<���@&l�m�
M��r���Yl�;d?��F�����/L�.S��� �T�g�;�$��wX��o���O�w��[/!�u�� �������/����Ut㠭:5RP6D>;�k<NUH�Jł�|�$ZiY��T|1�-,�WR��vܧ��Za��
Z<�����[�c�����{Z���~(����-��k�*���2�_��̌Eч����O9X�o��@�v~��5Z0�J�o|�I%7����'J�#�b-�_�֋븑(����2x�W_�<'���$�t�ZU����]r.[�]���?�Y=��[W��>�8r���Dׯ����g�I�.�H.�!zPAx��,�K��aO��T���x�&Z���MO�� ��4�k�Q�g���2��/rv_�No�3�
2�܊�]���n�ֆ*�+m�`0^MSm���o͸>ݤ9yP�/�����
.��Y�$��/�2�f��a�qZ%y�5Yd�m������2�%m!�A���K2��x����CA�s�����������'U�l<���k)>�NM��[�5�U�a��y�:�[(\I4���1Ћ%���l[�4a��;�Xn���
�:V�z\�,R>��D��P<U;�,I��A�9������i��y�=t�G;�-�&1+���;���2��
������=}���+�lh������R6��Ƴ�|y��ދ��jin{�*�-�:\�P���Pnv�3����;�%�m�f���k�\&��*�P0�9��7�(;� ��x�*�,���Jd�5�߰�N�=~�Ok^�����@]�'���C��w�;}.�ͥg�/a2�zN��{搘���e��б$�����N9�~:`����n�q��͘�{�^�ɥ��aRR�N��i�:VM���He�=tzA��V�ȫ�.�)nL�?���Ù��b$�L����m mY����+�(R�}W��ʛ���*`J6cn�--$O	���~�oW�~��e㦧a��ՓJ9�a��e���!�%�y|"�5L	�^���+CO#�$o�����\�Qw� �	�*D����䶜�{Sd^�;��70
���{9�p���܍i��$^�\J.�74��Y��n�Cb鸭D��3JC��Y��9�0Bh��&�����2&��m��ևY�������
���B�(��K����������'
���V��wI$��<�����T'�����\�*1�������_vRM R�vRLkD�:q�S7��h2	t�}� �G�D�?3�U��f(�0��-Q��e�!x��y�.��y\��ZX
^4�2�o�4��������\�1�=�s�pg@|{�������Th�	�r��(,mJl9��f��%)t�ߛK�K�n
�c_'��zE�
#�Ŵ���=V{X�~(6/)�F�de�fk>��}5�{J;!������O��f�V-�XN�D,b�C`53r_LW�c1x����dk~�as!�[���%r��{�� ��&x�Z���z*'/$ُ;++�p��Hf�x�p\1K��7)�Ω��U���{�|_��i������E�����ɺ�����M^W`�N��>�re`c
9�h�'�ANM�Jn��+�a!��7�G��J�^��^r�3A���ه���=`!�gy��	t��˔X�v�5����O]<�=��u3��?4"I��+� ��,������:q/�0r"���L��\2ӆ����~�瑝x�����X�����!K��Ӓ�.:,�MI�Ij`���\�~�e��e���|���
�����M�SVF����~=��̧ΐ��&� fv9�t���r�,?�hdޡ��h�n���b�۬I��Ÿ䬔8�����rAP�~��;�aʼ���&�YXQ������k�H6ex9֏{gk��W|x�V�01�U�/��)2O�/r�ر��Τ	7eX2�m��z��S/�K�$��S�X��$�q��P�}Ε�x�q�A��m�/�s��d���=Y7X��q������ӼBil�>��LK�J��G U~\<����Ih�,�&���q)�M�uu�M,�&��]j�-:Ԭ��6H5�9<l����wS�D�H����7����j�R�����6_P��*g'c����`l[s���'�M�����l��Tz�\Q�s���H�6���B2+�Ɵ�?�#q���Ï�R�Y6�4�����}s%��SèڑٛHg�����-Fߦe�#�G��R_q�A��ʔc��Ј��k�LsF�MqY�� �*:^\��|�Q����e�x���O�$�(J	9��3�h��5�2���<"oҩ&���~��t�+O�T]���0"�a�;�*1�R�ٿR�r��r��G����P{P$�N�T�����|u4����߱[�ر,_ӵ?/_c�|uҀX��1Z��3�:��byՌv�i�%#������P�N������&�"�/bk��ah��qGi�B���G��[���P����LJ������)��@���ͲP�_ǝ	�ePHL����GU��I���s�����b��8�[w�r� ;F�<���'��������<^��?��3���%#�Ht=bk��b��.�
P�˷�x����OF7�rN=�����w��"ǛX����W��!2upd�dk7�?Z#�~ï�@�{?�e�"��8��Q`s	���ʝ��b~v�A֔�,g�f����B;��c���T�&W ��ߪ�(�^3��M�97;?*hmU��.n�[��	���h�߆�B��O�e�����|��D��	�^�qJ���\<�⟫�m����ױ�қ�2K_׼[3��I���_�&{	,SY@�n�K��g� �.��,���u@Q�wwA.������}`�Q�ݔr����˓�m�Q;�LN���9~����� ��vl��GD�@S���C�زK����G�\n{�� Ʊ��T\�I�-���˓m,|�7�Sm0�%�F�К�!𸜝�����T�d��%���-A�B��2�O�j�/�M�ϔ�,���c�[Q��7QmV�����o�Զ.� ��$�w��݆���X�G"4)ǟq�R�c��Qy|	U����j6X��Wk��͙1N�r�H�,�4��D�R�[n�{��B�r��<ZH���|��2 _o}�����%=wS~;*�����rYpZ�b�)�4�$�p3��<�:&�{O�D�A�vڟ�_a]�����`���_"=	���oϒ3�Ź�-f i�O����!�Do�H#4��%���:�� ���E�u.��ۣ7`�b��zJ���,=9!:C5�n�c/Zg�/��G�,[gF?�~֧#��(�"c�����[1y0B�F�-���Nb��=��Hɨ9e�&���w%A�v)�1YC{>�,�x;��L����G%��F{4��-/r���������C�b��������5nȜ���NY5���0����Ty'�٨��Ui*ϱ�%{�S
��n?i`$�:�y/������cdjgfE���HڟW�Z�� ��%�K6ZA��d�0M�y�ar����$�pV�Lö��.Ϸ�J�rW�({ȥ
W{��i*�{����eB���㹿�V=�m��}8��xw-p�>�`� .<�*�
ڭ�6;T|n�O�� ,�i
����C���_���3��ೊ��،���Q.H����F�=2�䏞��J��+R˿@�-%1\�Br1p�K��K��?r�/"�D��/O�8� p�K'R�x����!�HP}�ߕ�~�o?�z{��r��k(4�$/�d3��R�7N_u�d׮�n�<?�|:+m��6 �7�2���v�%��+���J��M%�;�$4�_:�r'�����EL�9	-�����˄��]jsa�{d"&���:Y 
!64�*�#��B�%UF�p5�2���M��~K������цkC�/
���#fC+�
"�(���Q5KRm��3�?J*
�
%��و��RD]�rd�+&�`H
I}�hɎ�#6�$/I�N�]>�om!O=�µ*�/y�p
���c������+�]`�'�nF��¥GF�k R66��jF�)$���"$8���X�M��=X�@,�B[���u8/�$��%�^9��Jj	 >Y�>��|�*���2��+��QywzY���ډ��'M(��Cԭd��)�cԢ�J.�jk��Ѧw�C��l3�ua�&}�	q��o\�J��:z�U�ը��|+F��&�0��OT>�\��*��m^A���En@���&����`�|�df��:'r����nB��ҭt�ۗ�������	�1����j��?������U�,�<1���]_O������G��$����{��>��0S7aܵ���z!�����Ok:�����/��7L1�]X;s�����'�C*t��.��f�x*z�Q�F�$���ϲ湫����W�9�'���R��0�ï�
s�#����s���p��˻%y���;M�`ԟ�$�w��n���zS[�&�Sf�.Ā渨��*�z���ts�ޒ��O�����BI&n���^5hq�x#�J�{i�
�T����Ģ��0b��B _W���էaW�S����i)���Pb���
U��+V.��\G	���ܭIOS0�V���TR2��:D�R���A ׮�u�v�rާ�QH�e6�K藠P�飯����7�M��d^e���ۼ����cxp��w�����Z�b\�o����
P����L�\Ee�ް�_���o�<Rs���&��G�E.}׌���V彴p͗��k�P�nˑx�&?��нo���lQ�Kj6aGO��i��q�,m$�^��\9>*)YYd �?牪Y3{%Z���̐��ꆳ���]r:���@�v��w���x��Q9jC��
�ۖ3\٦r풖m��3��jT-��G���t/78p���׽��X'���ͺ�_���ͫ�^ײs��zC?ĭ��]�@�)Xf�d�����s��!һ�%�8
TU�@�<�v]���7�[���-�.,>w3��`d�����6G<��k
�-��e�䲦�8���EP�O�-���"�`��ײ��H���ן�,�&��v �N�)�m4�ff��ߧ��Z�d{D�7l��s2�1
�k���e}y��X�>"��X�>rs�6�X�	`R�+%㐻V,��`�u�ʻ�mg�PJ�MX�1�5���Pn-�u����Ό�{زYȭb��3J���*������(̀�TO��1�O�/�3bi���9z-����yv�S���*�{��̖��e#���b���-����b�X���/p]���H-�/^� S�16���m�]d���ޓ��H�v
�L	��N_����6ټ��	\��Kh/���z����bqz;��c{U�\T�﵊m;9$)1V��(��w��M\z�/����-��gq��Z.dό���@��vU�L�*����I7�8��� ��p�o��07�1�(]�FQ��P8��= G����.�Mi{��e��� ���{��]��+���x�6B9������em��~I�@��{��%��r���$=RVꖖ}r�.���q�=����+d�;���ֲ�!S�]�>���y�㳂V�r��]��P6��'d�L`�4~���6�g�Vs�í���:{]\��g�,'Т�;���ʇh@Eߘ�9Z<�&��JU�qT�\E*7!`�S>�{Ȣ#�5�@����w���9J��N7��Ed��L���i����P�/9��:XG�	�N�g�s���=�1&���A���H��+�Y��%[�a{�A`�E2x#�d�p���bj�o���W�4�b���˝��H�,?��v״٤ڮFż�t�k�V6�KN�p�����y�6���'Dત<����M t�cѓh;$R�z���2���+�Z�aH�Ҝ�_�V�遘�تt_Xw�4.�th���Z�\��I�uS�ʃ00m>^N�[j������D&�G�ف���]���6f3�؞����[x��ɧ*��{�o�g	��Ѽw9m~��Ц+;�D���(��D���S��|�:�\o���������KN���ҙvf_	�5�"�||�xXЫV�Os�
��$7']�<w'��1�H�+�IIz�ve�y>����S��X(�1�Siw{#�����)���C��6��eU��t���
����c�%3۲P<��T��qAr�J�k��gd�|nE;8�:��㽗R�Ue�J񭀈n�e)1,�=�[�gz4d�AlI���7i@�Ǡ���5�|�|[Q��Q�v����?p�b7O�L�U~����*��P��ÜlA��I"�VHrG�
 G$�B	�` �!����f�8��1�,:��_�+��>�	n;щ{ȇk��8��A�����!Jbr%�e��{0�����F��2D2��1�8�Ni1Ü��VW��[25��Dg?��;E��;�*@��Z4�
O�n������Z7�Q-fg3/��ɶ��J���ul	�&AM�b�n��v�X�~��T)1PCS��+�ڋ�1Q.�/�c�����9+�v��:���_@�Q�7w�R�'�ީ;z$��pT���P���~��H���7|�H�>�tLO���`�=��]�B׼�r�ˤ���G��]�C�a��Ė@H�&�u�Ot@-�.�\L�P�QbP�V�B/,����������6r�"*?Lԍ���*���%���Ȭ�k&c �C���R�z�~�i�~Xƌ�7?h^ݱ��iasL~�/�o-�G*m�w�������ќx�,�"���o��r�A�y�ߘ��u-����o�\.>T
���Xs/�?�텔�t��I!�Q���!V�k�����G4^�^��]IfЦ�#��4�ڢg_�q!�]n���_�~�� 6*�'�L�Ɓ_wfr�*.���
� �ݧ(�LIscۅ�$����*r�F�N�38-2��:i��E��U���+�q���[���Ȧ�q��yK@_ߔt����Dd@Q_t@�>n�(�![�0R>޿?Fz���V��85�X�K��V2;:w )�X�����d�a5ٷ��L����v�|�~��>�2�P��pc?�R7��7�c��@xW�&#ݶ���丟��JQ���\����A0�/��d��S��B�x��m]W��J�b��t�5v��8�Z��uI-�;�#a�c��<ٷ�ɀ*)��D5�$Ԛ:{ �؈:~�$�D�d2�3o�����-��چ��}!�OB_M�Gk�+Z���,����
x]X%#	2?�r�U!��_+�}1�&_{�E������t�P�RGF���2��i��o���NΦ5
���x�����5��ə���I�k�ez�r�og�6��w�3vxT��ǰj&�]'�����&����P�$g*�����8Z%�XRX����ސ��5��QS �7���l�7�n�J����ʜ �@�	�_�;hU��3� ��&��Ա��O����B����V��k}��>�0I慚(��Ч�e��/��=	q>>����Q�k֞�r�x�$���������I<�'�CO ���;���\�a�ɦ'Yt$���C�@��D��+�#�3�c3������2]2�]/����.%P�n�Xtl��K�������H��\�E��'m뽡��d��QR �Q�m�C	&�xT�(�/�9�74�5԰T1&��5k�8}/w�\s	���\D���9c|��� ������o$����S�	f�O��G{��v�dMXgҾx���G�2��D��<�7�
u��n��'V�U՗�5 ����]������꜕��gǶ���^1�{9Ĉ���=�3;1� ��ؘ��N��FT9;�*D���WbƐB{�q�M�u�i��pՂO�1�O�n�3ڼLrC#GN�W���� ��s|ԗ�4?��t�4��4�i��_��߰/wd�A��q�|>ye��'è:��U�:���%ٛj���/�o5r�x�h�\��EH�=�O�!�m�/���H����@���X\X2�KE`�.��S���:O�

��|ȝONnA9����w�7a�q*������|����PMm[�T)JQ@����� �I-TE�-�nCA��&��PC�K�%�J@Zh�?x�����{g�19��ךkι��|���R(ԑ��WL�8��Rr4��yi{��l��a}��Sc]�I /����$��栮<��{���Y�oLs�:��k��p�m�����A�V�.�^^j�e|u{Zފ8����Z���ʳ�����3�dh 껼��^'K
�\���?C�FM�����۷m�z�Dބe=w�P���:U*��8jqR������j������Nԝ��?GZ�Y`*���.��_ʡ��%�ی���xJݾ8�2�������E��s7$������.�S�w�vv��h�o��f,���4�F�If �^�47t����ӓ}�a@1���7�hE�ܩx�<D����cT��ˊ��F蒜A�H��4����g֗�q?��Vt���ۉ((�t���3<J�5�T�Ay���+�WD���i��W��������/�)%��E�I���^������o�7��B������W�qG�#
Fx|h��[�l�ʠN�`��W����:]z�ynJ3钽�	Ѡ��.�oߤ�g����2�^��"���"j~�b��Jd$�.U'�>�2�u���vv���?��(f1��
g�?q���C�CK����]B@v��0H��BD�\y��x�^��jc�5�%<�� ����J�H F7N@��ۿ��>��㐯E�Fo���{,j�����课�O������,� $��t�8>xq������R��C�G�����}�5��ž��I׿�S\f��1%X���p�Rp���me�'>�&�|��(�����h�{*c�Y~pO��JK�w{��(��c�TlFi�YS�	�ˆ
�F�fM��u�)z���{FG^���[M���l4b����+�6��C8���J�Ji�I�e��jg]����K|ictku�h��^�_��ʙh
:0<�HQ�J+q-�		��� ��R�b3�i���-m@&uyi���W�C?�=�=T����,�
whxp�DDX\��*�mjQ�d�����HՍ�F�$Q��������z��G_dvP ��q~~���@|ŝ&��U���.8`$j�xNb����_����gҐ�پ���YH�_֔��C7��KE��S���J1���������g�C��|Oʚ��{�˓�P7����Y/+4�k2R���p�v�P�wU(Ų�R�q�ypMgw�	N����i���m�9̹o��_+���Z#ך^!���5��1x�̹z:>^�����	����ǯLTD��Y�Gv�nNP���G1��+x������Sv�>�Vn`%Z�"T66�G���t\�	���E��K����p���J%�?Ow����o�k�1��BIs���|�g�"�.	��k>�s��>=���|��h��u���T�>u%��8a>�m��$Gy��o�oi�����g]����ק�	���S��9E7�݊ "�D�+���hi~��/����������١����?���m��gx5
@�Bڛ���.�B&��&ץ��~c��d.y����,Ä�߽��{1�}�K0����a�B��1�\���ڳ�4���.{}�>��#��a1M���v�N��s>��%���:W�Q�1��O�䞋���VM�9X����n ᛴ�f�)yC}r���i�O�),���g%�A%�Ɉ�*9�We��Z�is���y���\�O%����=��Q(�g�9�r2�9�?~�n(�R�%7�����B:G y�z�v{L��ˇ��<��I�u�-�&�z+��������ײ��_y���E{gF��Z����9k�7m�eU]�ؿ-6����\~߷5��Ha���'x��`�����̇��>2��_�
���t��&��Cn�,;��Ǥl�g����O��ƨ3��[8.Y$�<&����7������Y�%�:�������Ȏ�?Q�ɷ�٥�����*6f��޷�(��i�ﺗJ�$K2�ܙ�r��U�o/E�*^�i�|/<"ޛ�3��C3l/�Ft�Y�Jo�L�>�`���_+ y�Y���g��h�%$��Z��3M�щw��$_P{� |��#�4����}J�|~��ȥ*[P&������4��_%)��Y�:�Ȭ�C�0G.x�Z,x�Mx���ͼ�+�G��dR��K�({j�G��C�g�ʛ1����@-��� k����T��+OB�>���̷x�d���eVj�j��ky��s�<��vi��y�E5���+�%t9��(K���_J ~q{�~�2%�d�K� uׄ;gS"����
xd&��&�pzsT]�Oڪ"�zug���6$~$�"W�?�թ��ȏ�u=�{L*\�N��?w��s���^��g6� ��d�!���7f8[�;"��}5<�6�o�E7a|���9�zԣ��5�OlZ9�q��fz�(u��Um?�x����i}��f��ßW�2Es?!N�D{���^ɴuq���!��a�s����}Tl��vb���Kf����<�W*���	��~�@�Fʶ���54��*!��Zu��w���xxޢ����ᭋ�1Y`g�;a�R3��	�i	G�52&�����<yb4�!@ĖCW/�����d��Q!Sm%�!��g[�����������{*�Lg���ĸ��K�<�}v�c2xHF}p!�z����#�Qx���R)p��!/U3�|}��3��f���i��;�����~r�hEĳ�Z���U[�3}����2u��d���e�Ҭ#��9*���3�Y�*������Ωf�&��/�_)���E��8q�����͛��1q��L��2�ΐ����s�<���!����>�M�T��?���'g�Cm�q��������Y�{��я������+e�.�1��E��W?���L�Em+���si>T��kW�Y�$ ڣF�`�o����U�=���l�+޾G�g��R=��k	��J1�3v�kd�J�v4<�Aě��QpJ����Q	ٝ����9�����Cye�/����gϤ��PT���֓ݝL��l�aK5���V���߂�T�T�|j�����0��|E>�Z͡w.'e�}��|_C�Լ��Ϧ�&����$�a$��T���E�<�_��צ�𓶨p$��u��t���<�_�k% �!S#za�<n͓Σ;6�Vm`�bڹL$��U����g�g�{/-�W�:��ۊT�S.n]�6�wn��+��F��i�;��(Y?�.��u�\߸Bz����=�DanU�
�v�-���M�R��Y�V!;������|��g�aUy�иKS�x��wvtjN�k�"��6L]�X�<�O.ʽrC�7�� �J� �o$�\��p�$ۂ��1�������x�,]g����t呣������/��۽��ۉ�\�kN���sw���,[��j���2�ܥT����.�R�d�;oWK�MR��~����x�6&��֔�_���7����Z���#��c���7��H93oo[a7�����P���L�uEi����PO%^����h+�q��<�L"zά}g��%D����3w���HҤ��9�L�Ui���țb.�Ԇ&�T����P�l���U{GG̱x�)��9��s̪�5�S�\�5̐�5��/Q�{ϐ�Na�kiH����=+U��:�O�4�n����>&R,iW��(�mhl�6Ԕ&�5���?gC�ۼȦ\x�l4�l3f�%�#֭����Hl3z�����4.>w#��߇Y�ntQ\
%��ĐJ�N�����v�E�!��[�[Bh����Y��a�-��W��WR���d���	�}_���zW���W7�XW ��:�J�Lr~T��m��oҳ�l5G54k|�ƹ�s�6���H��I�]!������-���1�0w�ڽ0�Ai���B��F�G�4=>NW���?wy�j�Gv�uă�sӗ�E�m���~�`I�����[�u�[L�ݘ+��
������<�BzB�i�U��[�@bq��5~�{�G)l�"/�,���y_��̹�Hv_�YhVZ����&ĮO^Q��c��������L3�rx�%��5�,��[�a��c�6Y�g�4���i�7/�y���z�dVf��5���mM9]%�l-P�v1�f�aae
����F�Ñ���-:����1N�����b�/;�߻5m}$-ݘ'��1y>h���L��{���8���4;}�$�ʹ�~ ��#2�dia	 �V�Ot�{�_�b������H�Gk=�g�LùE_,�h7��0�Z�_�x(����3�*#`=��q�S�g�q_�s�'�~��N5���0v7U8)�t��ٓ��9�����<�y�ȳ��x��!��xoX�յ@����.�&����yb�mO����pXu�6џ��9�y�u�7���B�-�<{ߑCM*����N��O���S��L�Y�4&�P����ֹ_�BZ���?nF+�M瞎�mp��V�����n��tL<g��|O_Vv���%���]o�8�p��p��21z7�i/�k{�Z|Y��W~d�,0?�t��'WH�����O�[ lb�iU���v�e8��_$���4����S��V�&��0X���gx�*uqt�A`���@����$��Z^~OA�ā��x���]5/@����K1�b�gz�k_��ήD���&_%����Ɇ(�=����������;\,(:l��@1�D\s�<or��۔>��L2����NcP|�^Jq[���7������2����.!lDm܆|e؟�XGz��#��u�!��A�N�ԗ���#~e�����fj���M.uq��̿+b�\O0rT�}*<韌����9��i��FP�?���0;���}lU���҇�%-/,at=�uNj=Tp���@e��@i��W=�<(�ߣΘ���㒷t:�c��%E�@�%�՟���L��(�g���Z�/C���|��5(�����Ru�x2�:�{��\lq���L'��˿�D����0i�8h�ER�UƵgc��?c�#��TM�{r�6�䬊�o��j}�,}�]�b��PJ�rw��N%L I�������?wy0Z�H[y���OZ;-'4"�(}I"��9�|�U�ك���jb�3�_=�ʛ�/9�>o�0�M��J������M�ț5���D�+k��b+��_�Tѥ�8�=��]����g���(��*����]��/��}y��d��7��%�q��bޜ�Rk��ɀ2�Jk��K [4��me����y6>6�O҇|L��]�nM��yH�-oWgi�(���b~���E��.���S��Qy�wʼ���o�?;W��0�>�n��v�zQ�?Ejw�pƢ�r�?(9�kVh�r�)��_�Q�s>�h߂7�%e�#�U#ܜ�5�Z�k~������V^��7���	���|�9$�,��7Մ	z�ԅM��Y�y)g%��8���Ն�P���� J�A@1�cW����CP@�Q�K����}ʂ�--LQ��U$�����/��	5���U"ǻI-(�Fvj$����*����s�F�ծIԳI����.�V:mʱʔ˾�+���x.Kt��vg�{5��N�"���A��5y'�;ט�:�����Fdz�����8p�ݗ�52c�h�z�G��
��4k~�_��Z�kX�h8�,xe�~��o���S ����F��F*[��L<�_�k�ְ>��J��W��k[F��j<��^`C�����6�@��~�K�҈��py�&uuPk��l��R���G ,Kn���?���[��1Sm4�*��m�Fׇa�r�ua<����WCZ��vj��6��Yi�3wҨ/�Z�<U!�63��% �?��;�~_���4�@X)ni�}f<R�H�2��`4���dgf"�!3��/OJ+��۝#���ܙu�H�Xt�c�"����Dz2�M�-�5+��+JYp���%Qh��x�pr��fJ�H��]0��x=��BN���<o0W���1�
��Q��H���)�?��\б��,�<	4�^�d�Q�����ɖ	:d�Y�Zg@���e����S�������*s'W�����C�G�,>���G^~�	�������5C��em�◪�����L��nGEk���G���Qʲ���ݾ�йc-;��,D�@��Y�x����~���iގA���B[Ŝy��x�8U��.B�/Q��A���}�h�c��"� �f�Cw}|7��/�f�h��`��a݈�I���j�Ș���H������u��3��6�Υ(��r��#���q��������%����k��j<��;�F;�S�Ǆ5�{�xL�lDH��9�2�Cڝ����q��	\���w�}g) y'���K��	���.�f$�+ݥ�ұ?8����ȏ�l��o�"�2����$T�^J͒7��E�kμ&'�>Ĥ�Uŝ�H���>͆u�y�
Oa/�v�ZZ��v�3�Q3���˂��t��+f�Ч+�M�;è�bV��j	���:������5��_��opOĞ���py!��oޠ��b��}�_���ύ�>�{��@�}��,����?�D��߮j::5l)�\/;�P�)+���ϫB�w"��~���~��N`+�D.T�K�I�_%E�w���/8��p����em:��g�T9��ϴAA�Arn�YH}ï��t�ic�3O�W���iL�����ޘ��Q����fh���Z��ʄ?�(`l�2,@�M�6-���p�zH���p��M�s�!}O(����'	\f'bK�+��pa�����)A�|���>��qעU�d��������]K/O�ۛ7(�����8�V-��S�FX�J9���o^ �u�J�A�ڲ�_��c/��`8\2���$aX	�gbb�=���9r�z���)��8�Zx4���Jo�L"����O�F\��K෋���>C�̨���3�V�xx���	�Īy�ʒ�qY@�$\wqyL_A����R��~`R��S3i�Mar�.G?�x���$�?'����(4"��ӧ������Y:�Ag܄ La�¯�2���؏�a�=�paG/>؆[��'�~~M&�,�j��_di.β^O���O�4�Ms�6Mq�CWY�$�e[� M��	�oG	� ���EԶ����8uy4�i���\'%�1꿐���ywÊ�=��c���S�OA��R��ok#n��o�ᄟ��h����Dgb��0���U��*�]�n����Λ=�P�5d�1"�g��"�X�w莆]wy�,��+k�����n�kd$v��c���5z�3��8;�^�E�B~,S_���ϋ3~��'S���zp�KV6vV��K�ޢ�xm̒�S%��1��^�������{���k�Up�PQKɣvͯE~��R�e�3�����6�w�l{a1���$��?I�"èD��?=�i�:��~T�=�h^|�׋-
��F<���1	��ܩ�MRe����s��}N��3����Qt��)�NO�B~Ѿ �%���D�"�[k#��~4�8�c��*S�^b��.�%����
��=�5��sk+��$���y��
[�p濗�����u���
�F
��D�;����������m�A�Ecid�-�>:3 9W�/�N52��'��/�R_S*��G>�������1���¿y?�[{����7�F��/$,�mO�kC&��G��tM*�gP�XPy��ˋ���d_�~1У��ȧ0��bw�JkO�����J�ee���VZb^t���h��Y��Q���7���K���v�z�𵮵�m� I�k����/��z'4f�"���L	��&ċ���$�WB¤�,�O�?_�]sa�a�z�Ɛ�>�i���-7��@'�~N�����N�hT�9�.���mĚ�Rڅ�c��J|r>��=����2|]�R�b��� �`�h\�
H �Fn��z̾M����gG�l����P;~=D���P(�W���dCQ#��������\>�������޺.������r`m�7���T����g��e��56&K���/>kE�ðA�u)m�Nub@��	ݘ�gG[\�eĳ�����"��L�������]{j�)�ms�[P�"tm*�[ $ָC�t�K�{�35�Z>3���`m�a���ɺy�����tG�߲Jn�[Ӻ(]`�bJ�1��?MF��n�+�`"H�8�}��34��tG[cX����G}�ؖ��z��@P!�R�A�:烱�/���˗����OLB�)9��6�?#��Y�N������o��5CT� �0�4����G�c�#�_��m�����~[D���B��]\ō���F���P��g���tR���sy%I�"v�$�Y��X��~0�k���1�m�˹{�5h�pԝ|E���CX�G+��6GNK�j�Y�j8g��xC�x�W�FH�B�O���忠��+��c榏���Wg�	��Q.����a��4A�}��"�B��C��C��{�IOU��x�ޅ%oU���R�w%�^��H�G�'�Ey�[�II�/A�X��S@5���&��[c'�a�_^!���za��gZN�6OƁ��9�-j�NG�v�	e�Jz7i~�/��&�x�/��V��Ba���K?qZ�U�7��79�����T�N��}PIӞi(YZ���E�Ԓ/s�'5��Y���l��L��|��&�:�<�Jx�o*�6�����v~T�j&ni_��&@է������-�}�TY���k}Z�����p+�!����� *V����f���75���m�5*�L�W�6	����O�����%�������Z�Ձj�?������=�c����jh�ԡU��Xq�5���U�9��|O�=�[�$���E�z�eq2�7�!w�����y�0e5�I`��݂��+������=Z�5C���=��{������C���q��
k��aB�m7��`�9�	n^-ν�'R��N{Z�`W�t4u�����p��bAj��%t���C�۵	��1�����SG�I.��GzJ7�<�#,�{`�7����Β󟛶K���=�{�k�$G�u�^
��Z����{o�8���'�2�z� mV/	G�0�d�Ȣ dU05�0�"tA�q�	�W�Ը�
�8�݉��x8�KR'��f���RJ�T/��9���R{6i���$�0)�,Sb1T��r�4���MV�����*� �7�R�9@�o�N�"��Nh�kuǀ�-?��o��:�PGDT`\����D�o��
T�|�>��.B[�̸(���₦2����Ad����׿/��F��n����ǀ�.�4=fJ�N �)����>��^���>	h`Cv_��#^����-�]��k���Q��N�Ͷ9��Z��|#�48;����^��2�ݘ#�,I,�`jR�~g����\���E���z�@Y�Q^����̿@D"�}F(к",-�Re���R!Մ�Žj��T,W��%D�\�+����7o`4FyX6��.d(�@��198�ꓨ�A�zL���[L �' '_@�|�f�"�jPG�I���p_��O��A���f�����3M�;���2����ݩ����J�a=�����q1��rW��`7�.M�(m�_�SR�|1ډQ_/�ZWL��Zzq�`Z�p�Oi�=�0v�1u��v�S������?�9��P�wAN�1�Cwa�}���n��.ѭ�gw�؎.<�J3�����'垨:=���>��p�)kE�����	+�a�)��ԳG�R�`[Y����e�j��:��5�r)�`��E��.�Ĭ��4۵.g'���Ύ.{�!�0��~������h��|w�0���[4���b�!I,� z����@�K��Hӿ�G�U�<���m[=���;�5��'ގUA%�$/lu�(a�G5P��k�N��N�w�K��'0@^0�������f������g�i9Ӫө�4TؐM,�W�.���)���/��~�;,�7���D/��/f��L����]��a��B�<Lۂ7N� �E��B���%���J�<����(O����p�k>0i$�ܫ������Ӆ� �G����Fk��J���Ρ�I֠�O�~K���V%���oZ]K���&��/p]�7��՗����	l��.�Y��N�<��û�=�Q�f��@�����񩡣�wы�p�Oo^|����@�j�Bm�P�JTyCJ�>�B�se�%�ĺ�Dc�k���t����+��43*U���v9��\{m5�iH^oo�cQB�����B���^���9s������q�nA�ԣ�F1�M�YP��pg^h��&������|�Y#]�g>�����ط.��ؗx#L��觲��6���X���{��JSXv����{��
�𪇪p�XM�L��n��5{p㧞��֎��<�BQ3��"��F�}J�p���U�>P*v9���n�<���yD�ը��~�ZW��9p�fˣ�h��GC'�X,��X2+�8-�N	����|%�c�����UG�����B�KՀm���p3nA�5��vY����
�
��;��G���w��^����:tC�T���f�vIO���S+SJ_r�;cq��Ό�����k�����SW�3pF�CƼCY�*5	#Yv����OQ�	5�=1G�kE�7e��#+z�^>����aߟ\��e�r���j����[��{�+���[B�;�7��I�@dk/ͤ@C�S�u1�O�����9���Ϯ��y��i�H�Hǈ^b���$�P9T~*�&GK��O|��O��ݮ>Z-�="��u�X ���4��9�����ݼ=��)eQ�>o�rzx�@X�/6-80��5<*=�j���|v��K�uc�!�46E�;�*FA(>�U:�%�"�r��O��CRA��y�aw��X"WH�I`P:�Fm��|��0~�l>�/U�SV�������	5�^�F��Y�cդ�DOdr�*p¤m��<�e
0���rH���Z���ĝU�MMnuRM]5Ս��IS.�c�i,���{sw�]/����g*jJ�H���ի}�K]�����bFL�����j�S{��W��x�T���lJ5v@4i.�~@k�g��&��/�?�j&����*]��:Vk�-.4�ϙt�F�Vp�z8TO=�޵��zJ?��s���`�� �7��-�TV�~N����%����-�
��%�+<����c	2]D��hR(��P��2!�*�eܺ��K�#O�[-�g��A�|Bh.�l��rއ�:b%�Y<��UU��BFC��c�
���尺&5��V�~۔k<R�˝@2��@<�<l��n��NK��ES�:�[�^��	������8:�;����ι�^�tDC}v�;�恈��ح�(��G�I:�g�+���w�9���x;�L����$ !�n1�8Ts�����%*���3���q.�s�v�����N�A��Ԫ5�ԃRɟ�*3%�3�.=����ӻ8�ח{��]P���� �	�����ǹ�B�ȚӤ����t��4�3K��o=0.�D�d����ŷ�ni�Ud7KK��	w>Iw�$`��N���]���s�C%"�T��>1�1�s������K�A4o�m�k��f-�e�R����ШX�F2�H��2��3Ջ�Dp�y�NB�pC�QFMWɝר�|�#��O�E-~���=����^�|��.U�QP�]��&���҇�����=�OH7����  `������2��� F�Zc!��ߎa�Z�NsKJ-CkX������xP憵��VM��{��}��Q�q��R�3PܻYj�|C�9�P�g��ؼ��8��-XTQ^������9�
י�{�NY��p}�lӱ�r��>3�N���@��E���BV)�ퟹh�8�'��&���P0���ݒM�Pl����V��8r��^13�*y�3GCh���D�������KL��A<��
��uү�e�nmE�� �Kӎc���Ő�g��q�2���l��:�@Cma�J�c�fa��:-~h6�N�iF�j�O"u���\��qw��Jx�9�!U�`�j7�<�Q�<�<��YL�-�;��$)L�����\����_�}����\����ܱ�<�(3R���!E�Ӵ1� ]뫣��3!��;�f�ϙ����2�`�~$�'6���u�[9���
iWL�"όa��_�t#�>�,E�8&��&��';� ��P�x�+r7�T/RR��'Y�^D�u�D�@%T8�a�$
��d�U��!���c[[����ꃣ�a}��ZQ�X�T7wC�cK�Y�e�]�a�o.��b#R�G�8�c�r�;��|c��/���a�l#@�J�M�r��J�0+�O�	�q��~�כ��)�*�	����� nɂ��jj�?�*�vu\|brB������a�ǜ�f�B���^R脻�ʣ��|���fO�Q��h>���l��W���0KY��'kL����n*5�NR�a����<_�W��T�ݜ�i���*p~��j�1M�b�,����`���ݤ��o�B��Sv��Z��iqA����Q���c����4���yQ	�i6Kv)�t�����B�`\�$�f>�tW�Ƈ� �W�����!85�VW�CHP��@/j�2<r�#�T��r�_��Ъ�і�F�;vq
�"ࠐ ��~���P����c��F�o�U9���>(������E:MJP��X���|(b��NL��4�TB>؃ۓ7K�P^ukk<F!��}�a�uS8��	�����z��!��tKlrf�W�7ڋ.a��c]��<�]ǜ�M�N}����������]�L
(]��z��4}��^K��	h��-P���L�����Mܛ��@z����N��"Q�[������j��\3��[��T���+� HUg0є�]Z�^��U0?�ל!�4��p�6�l� \���$Zb�uf�8��@e��w�Ftr"�Eg��`�&&��s¼+��x  M�H<�X�K��$u�����5�X&��i0a�f&�4Q�NwB�1���)�� /��,�
�~�٬�m��k��T�!�Z���siܔ9�𧲯>�1�l��8L[,���g�LH��k#�sv���ׂ�;�l��E.	h�4��i�9���3]�+]nmV��a��Ѝ��٘7��I*=3����zMؕ�.�)�F�q����b�./�LFCx5EK����&@cX'M�f���{|����h+0`jn@�ş8��<p��!}�g��n����,�G�b�  ʐ���ƺ��]ߡ�s��EӅ��B_c<��蒠�ۇJG^�"�6$������@�n1���h�k���-�<�����}�����>.�?�
[3�#yj4��W���鞚_�0a��������3�����,u�W�(�@Ӡ����x,�,~l��:8R��z7���4��s�v��{��m|j5L�8�dP=
��]FJ�Ew_��ͤ�����l���ꤧ3�/�4���z��f�B���oȌ���"!��/u|˻B�S��p���M2#��x�δp���n�g���<��ζ�n�1l{T������Q;���ٓ���z��n��r�<	,��G�R��h��r��܁��)��̀)��(��E`�(UK�T��f�Q�wM���Q�,~pw?��6�w<	$-R*�G2�ӳ�m��Nc���<��a�fd#(�Z����'�.ܗ\�9������x2B�T�r���dVN�I�!�qg(``n*�8I����H��AOn�MA|^ژ("��`o�����6��;򢿰w�^h��E�$�	\!du��}�5��b,���� �C���||�R�|ˆ��� c�5g�wl��[e	���.y�4m2�Y�Ì��7"e�ivM�������E��V4Y�k8|���Û��;ʆ*C7�����s��O���*�@F%d͘:���?�-��}F��N%�e���� Z5�����;og�N��'�o��M&c0��� �w�>2�2T9���|Z�X�������|d�q��� ����Kw��j��*�3.:N���x��(mR޼8p��b�M!f+��S\��V�z��~3;�KDt�¤��3��i\�l��u�O�N��[M}�gZ���ʇrS-f�O��*G^;��4g@*#�HPcw��+����c����r�)� ��(�q��*c2{�[�����f�g�5�KI!I�,J}�u�S4����L}C&�zH��T5Y�'�G����Y�Ŕ1��d}�/�����R|��\b�H��ޥ��Of��q��z���9���ú�7��~�c�n£ܫ��[�@)�NǀvD����I�0�
��k��!	�,�w�i�D�0tH���dR�C�zg?��3���{eH�CN�@�4��lu�g�S0@f�B�,4�*�Q(o�u�#bܠ���w�qhp ��dA�{�И�Ң��叇/���U��	O<���y1:��%&Q��\;
�Lr۲�c�n,��"���p��S�H���ձ8���<:��P� V�����^ٯ㻊r7��J��"��(�y����0+��21�Z�^[k�.��?w/�Jnuvܘ}������87��Rz�hiX��6[�_I���p��s�f)IS2#W�o��g�T=����*U1f�'��wYv����n����	zWKлmgc0��YFh�>�_9��  _�5Eo�r���h��J~��f�����4�~*�Ŀb�8 X�/k��e����1_��x���7�?�Mq�;�b�N����["�0]WO����H��`KM\���r���K�bK��J/��������ԉFN&����!Q0���G ��dQ�N�@"x�?��z3�	ϭ��!��b�1`��'ʚ�xňu�������T]`��T���z��ec��p�p�3B�][QL�|���2��ِ�h/�"��P�}�"Lw6�fϑ��Ǎ%�<<L�Y=38�R���R���|��s��8r���{���@�e��x�g�؎/�X�<.��WFL&��F�fوuo')4!e�h� OW��k���ܟ�B �J�lNǉ}�~47@{6Z�tmR�e����D6�����T"S�$x��v�D���B��Y �}Y�E_o�D�G(2���})��f׌�|�I��|1N����ڡ����7�+jVT�[�hR�jY��x}�\�$�0-R������/�E�b_T95!piF\E2�b�Q�0�`���L���%0��KG�f�/`>S����|��$Fc�J+]�C�	��A��g�23�ŋ\L�WM��пN�㲛�-�$�h7�23:Q3���{XN�L'��6{��JN�d$?X3�:j,��0����ZJjιL��R�Zg���p�4�]�i3V���
rr�����U�L�J�G�yE�ql�����o+/�s>�S��6/�T��z�+�h��{]@����[PF�j=��*(=��.im��x��r0�2T������p�ݴ�0Z�����l�p�m��S;v����t�x��{�辵�$�|I2y>d#�<!lO��.����s�o�����$�*t��J2|4I����ϨDҒ��m
�Ҩ���a�^b�>�&���W������<\�Ѡx�E�ޣӌ勺�8���h�^�0{l�/�%�Y�9c++g{�o�l\QܬF&�kĈ�y1ź�A�L� �*��RnU=����� R<�s(߯�mS?�}Z7\���n�5VG|[z0#T0S�U�a?T̟�[Tg7�&��'�Tn5E��eID��{7l���Ʋ�K��K��t ��|�r��K�s��,us�0j�i�1��J���M43$� z�)�<
�B��`̊N6��i��o|3E,#��@|�_�9x(8ͨ��"��7D%�ٚ��6Ժ�6};;q>>mj�"�e�&����H����m��Av.x�Ko�����$P��5cQ��`@o*m�s}�ߕ}���E��u�-%M�Ww��*��e��iv����Y
c�2�n;P�����*�<�a��~�F�:���s���DD%��=D��@J}�e}�y������j,�������Eh$8��"��Ҩ�[���:�HQ!�ఞ�^�a��9��+NN&E��>U.� ]�+�U��i����º�W���
� �J2�UKï ��Eɢ�:.�ҧj_�;7�ƭ� ����k:����T�,@4h��q�j�&*�L�>.���ve��o�j�� �N��~�����Y!�Z�Qu���G�4 +#-����B�5sݠ(�<�͜��dȋ�G�n	�Y���v�*��Y\�ں��.��N"��F�����bƌ���fTwO���j[�liVW��!Xd���y���uY�������K�p�x����\x�Hcg�����#������MI�u�X��ߚW������6=�Y�l�K��h�)��ūfԚex}C� ��T��ǝ!M�ǀ��ڊ�Fa���|����b���Ypl{�k�X���6�x�9(]1�^�o�RrO����(���x7 մr	W��2mP�5k�tB}T�y������ZA-���ui��&g$��O��-����C����-
̜Y��|�/W����[m���C>t.�>E�2:�s�/H1��v�A[V�Y/aG�Ή��(���%|�C�g��;^���Є��6���e�Ȗ�E�\c�7���v�>]��▟�n�+0pqIG&�Fo��4�z�O��TǢ8�N!���yrK!�`�T�J�ފ�*��t�P���6���y/�z^������;�����x�����jS��Y�kW�U�F�Vk���{Q����m��;�U�����1� �/}����������\��9��K�f��s2���-��H	)U�6(͚�x�g0���O��N|k).S��*g������{�dЍYư���%��큄.�# ��%R��egM�<�����ki�s�[�ƌ��_�f�}d�����ƿ� ��}_�Z�燚֌^m>�nvW��%Y��rh�$Si+�(��T�{�)V��x��쟞!uX�-��х�:L�R�[���]�uw�Z?z�L�]_��%����i�l�`����wMq�6?�uGfM���*ʆ�/�ڷ�6n�<4��T��w�����~������ַ��1F�[tL㧥�YY�-�3W�oѝ,[�i��i����3��=�dW�����uE��fӏ���+'~O>L;��;h�1�5G�!�5�i�:Ƌ��cI^:���n�+7i+C���}l�G�/�x�L[�]�M^_U��3,"p�����}rIe'���v�,#����:඙0ֱ�=ͺ��6��t��sܚ��������a��L��O�p>[1�H����L�+��NuG]���u�&�oi�1��t:�=&^𛶂}�F,颼���,3m��m�6j�u�iB��V)a{U�Ռ�AgҠ��8'5A�TF�RA�Y�A嵇��R�8q2*��d�/��1<�n��GL�Q�̌ �D�L��}X5�k�n�u����ӣ��}R~ɹ�<�[�|
yJ�*� %�?�F���~϶��q�������8���+���j�V:IP�/�(k�۱��0�'��Z-_cA��mc9V""�E< m+�c���R�0��d�=
Wa[W鶀���*�*���#t���c[4z�`���o�Mʠ�����f�&�)3tB]�?�+V ˰>��x�⡟F�vR_���)���l,�y=ә���.�4u���n� �L��z�i��ѽ�bjYU�7˶�f��� BӖ���p����r��8甩�B�X�^�����$Q'fE�r!U�����>xЗ��-w��xu�g��}y�p�8oF��<-d��I�rA*���ॾy���|�v8��^[�;JR��ӵ�v�Qo���,��e�V�����nV�����̠!�@WH����R]�
)�A�5�>�q��
�����z?R#K3L�]<�p� �^J8�|��t�,J�f�����t.��]�4�*fx-�+�s������A�ɂM�-綴���'�-�2�GyJ��������kJm.LZ9:�t���x��y���)�Y�%�~K��W�[�� �3�O�;�U�c�EU�[؎�{�j�ݥ̬�
D--�T���*]�\Z����}���z�xz۽��IVh�n�aX<���/?,2�����%yw�D�ǰ�rP��k�M7�o�K��7Aj���V\�̲�����lK
�r��������M��5+�;f�3ݏC͸�;��g{��>��w�y�����腪�U�wf� ӱ��4��0�1?Q1��r-�3���W845�I��K�X��<�-��x�hYu�q/Lܚpy�.�:?��i�-�!^��T�br���g_�b���PI��1w�lPj�D�Д9Q��p���;��������p�a�A�x����co�W�r**�2��1U�	��}�9�ɳc�B�P`=\�<����ٺ�/�y����%Ng����d5�φ�8�H�ތ���7`�U����|�k0���p�k��{���3��x.Q[�sﶩQ���tf�����0Q�|�Y�3]9W�w�q���㿱�o��t�/�>�
~�ka����Zp]'����j�
b��TN_Q��ޅ_��T�F���0ιHk�'M������Aw�2�B�N/s[��{�e8zS�u,N��kFyU0�;-�}�����w�������<V%����k1���U(5O9��dl���P������P%�x�M�U��m(
iɀ7�g�M?�
���i 	�Y�l;�T�~Ec��ȝ�5O�ң��+��>x�_^#�-�2C��B�/_�n���ݾ��LxdV/0]S��˝�*�F�g�t(�Q4X�K�l\-}�͌��9,wi`�Y02K��I$��5��,}>v�m��\J�e�5�E�?"�8P�X�
i/۹�i�4Tl�&�9[�&jc�źn������u�w�����g'��8{�+{jV?�QMMyJZ�~V4۞��63���_Ƙ��d6�X�N`�W��� ��h�:�����nu�V6�O1e���0ÅG-W�I�*-ޞ>SW�Q�f邯��k}-�^N潳\�
)/:�qq�U�I�Թ�)�L���^;���gU��'�&,�j���]=�z˖�5oW�aȝ�QT��̅�Qֶ����3x��ۡ|&�k�gYM���鮐��e��y����*T����>���I��w:AJ'�����M:���aԱ�(Eg�^�7���S�J�u�]6Y�u�2M!����m��/'�(:�t�.���J��?�:h��[O^?��N-7��hS^��|�r�9�_=όg�=�|�������c?,m�_�����f�es^|}�7�>�*���ẟO�\�HܶY}t�����]�A���Cto��_u�7�=,�f�PG_�0�������p[��^ᓎ��YȞtsY��rU���p�Q�'	G����U3?|��rq�j�c�_�����i�W�_|�q��K��{v�I:�?�PP�7�#��ul�,}0e��}���~$sƢ�2֩�5(��a�#�=�|����lO]f-k�{�����\&B��b��SGs!�m�z�����?ͻ�J�.�4���?���j�����a]��X2uS��������!]%�hR��˥���R{�7I��4���l�ג'L�-�q|Z!C(��mWj��ٙlA��X��.j{z�5})�Z3���y�D�F�O]3�'�1't� ئw�������f1(,�⾅�y;5r^�	03�Ƿ��[�Y�KMy�Z~w���0	�;��ke���c�D�X߭��߇�?�B�-H�e��/��NN����#���A׈,Z�U|�l������SZ������Z��`4ï�C3vM��YQ��ٙ����e��9֪_��"9�y��]B�e"��j��J� ��9�`�����o}��P��p�I8��C�Qe ��� ���� ��lvj�p��-��s+����콐�=��ԺfC��~Nl�����Pd1��>��24�QC"��х2yG�~Ua�R�)�s��1��o�O����!Lh�E��B�C��5k%8_���n~[��Дŀ�D#��nJ�'��R<�(����Z��q"M|�>�~ig_a��L�����87D�+R�k{ܶ�o���
C������l�؝*�}�f�lA�.l�U�k�Q�hX�.��k�}ݖVc���W����2�X�����������4[��b*sn����$j�+����*�O�v&�����vya�_�`Q��p�`���Sg[YN�����Ş'����^�;�&[�@�I55��Q�woE#���Z^^����f �}�D9��+�Ȉ�Oxf-��޻v7��7d˵�9p�a�D�����zy=z�W�4D���%QoU�}i/Ϟ�k�#���P��|I�$��	������oJ5�[z�'u|^Z���S��H�T+�Q�����-�َ8Ҋ�RQ���!8�t٥����窊�ʜ#�]�<8��etux%j̓���v
�"�(�����W�v8���[;��Y�-)k��U-���nZ��2�a����ד�vh�؋4ӂ?O��c�-f�����)#���:�<3W���Y�2&c���^RF}?4�X]�y�#�ٵ��ɰ��iw���
�%��� '�-��vҡ�`!�@Qc�����2t�a-¹6��So�4�_\�T+��(��ߝ�^�� �Dz��_�.=�P�a,}Ĝ�F��p�b���Qv	h2:�r�n�[�5��Zߗ#���N:�Z�.uXqE�ߺBC޶G��|u����y��z���ܓ������G�����F5̆��RQSd���Ф�
�(�Z�����$�a�T8�s�I~l�ż^���� x"$����^�6]%Q���o�H��3�Y
��T��2NM��ƶx��,#��Qk��o�]_��G��<�(l ȝϸ 7wA~djH"�b���
�Hxۆ�ݪ��� ��K�G���w��EO�����^�\��6*SGwQ��d-ϑ�Z������]ڒ0ma�������v��H�.Ul���2T��"=���Ŀ�('F�dq������3�A��!٦��#w!�@}�[�M���!.�� eq_U�o��@_t�T�1ר|X��x/p�	�"��<wl	��|����-��`�����n"^p�7��n��{��N3���\x�Ez�yz��ʒހ_���E~�s��I��r`A�&C�{�;�l�f��8��]H^�Ϡ��i^;����M��$��e읮O�'[�����%�/���!�7nbX%Ԍ*+n�����u8@��wu�-�$��	�ɋC��ɈP ��2����Ս�Ӂ|�5Y������7�|�������/C�������r��Zj�-�-rė��"l��hQWQf���Ac���h9I����x�
�vc^��|��Q>Ll��.��Cwjoc!d��<��U5�,j�Do���u�*��w�o�	?`�R�8��*od�
�9�Nh������l��
D<�|:;]�=ͳ;�"	K�<͉ѝ���h�U�@D����\�EE3<���FC,��qS�V��"<U�A���TP�����8��� �k:���=���Nvc���7���\�T`����<z$7G�K:!	3���d]����1o���<{�&�+Y-ԝ~�ٶ���u~n�&�ӦAwսzU�Na���wk��+23���d��V�nq�Gu'��U�rh(��g�h|^�����?	gY�v��smdYK��H9�L��X[���B'z�ޡ:�JXc;����N�c
��T.��nl~u�goz��=gU�Η��̹���7�����!�^S����dKM:���*O�����?�lk�<�1��d�������>�� �цn����Q{i��Y�lM�����]��K�q�6On�s�������B�X�̪͢vtB�>u~N	�S���X�e��p�'�-fz�]�,bء���3`��n�vR���@��Y|�6�P��Ͷ]6���r���n�7����nۙ�H��&젲�3P��R���a�RD���3=,bP��7~��]�C_�?n���'���.���Ho�\uO�\JV�����l�f$�Re��W���ʫ(���O��fN���y}�j>�s5_��`ee&��$88�k��zP��U����i���5���3(N��#-��Ƞ(S��L�|~i
3�>{�,�؄���$:��xQHd���'��>��n�V��l�t�K�$ۻ4����H���޵O�KZ\�� HH ��<��Lدx�&�]2#�-�N�S��8.TS�3U�T�qO�DO8t��P3�.��WI�3���1�f��>I��g�,�"���K�LH"b��������F�9fzY�~����K�^�������ds��⻳�C��u��־��*Y)�Z�5�}�s0s��m���S_�J�����7�-1�@驷�!AV9ɟ5?�ߪ �u|W�_.��5��H�u\
I�33v���q�����Xޟ�ϾL�DY�^��~}�ϧ٩�"��4���m3�8Q�3@GΗq�=�g�gsu�����th�ɣ1x�QVÉ�W��f6����Lk�]gIC�G��\x4>*����y���=f6	��?8��/���w!8|�7��l���p�_q�	G�q��i�\E(�G\�^1I�k��{��v��[���\��僋#R)�����]��Tm����T^�x�`	{��t 2�wg���"�ͷS��#��]J� N5sPT�#g`��H��F��3/���9��O���9[Ɲ��F���Q�;6��,�9�Z��6��*��ww]	1��EG��3C�O���$WL�R,1���y1�v&׍f��y\�;}�i%knj�2noy9t��T7�GY�~jn������G���Ҹ�X�ow(��	�Gc:�I���Uz��p������O�Ti�3b�g���e[��H6R�D^��Ǝh�-M�;)k��f�RE�08��fmZ2��f��ߍ����R��s��f�{<��+.�0�3�xa�լ��B
�����BЙ���&"���J��0'��`�(R06�aH��5�_xK�<7����)�>���JV�3�"3�"���6g����u�nh�Ha�=�R��{t/Ew�����޶�P�b�ꂑ\'����Ӏ�a�d?������!7���g!C��t����I���]�͝c]^}Z�SIM��̈�s2{mwC��wU�Z��0�������N�	w��m]t��u�D��PF�ѱ�	O����d%W��&���N�p����۽^rp��~�
D?�8!��i4�������������; P+/��B-G'ݽ�7�,6���%/>��J�M��e�C�⑸+G1r�0|T�iE��2Y����G�� �)�Ia]��1�p
��fѢ�KS]f���s���7�S��>U�3����b�ܲ|�A�TުJd�΄ :�����Z����6���~��54F���}U���9�엉T���Ǝ�w�pYՖ����sx��j#�ϯ$:L�u���`�vr�tx'A���ʣ"]��t%�����=�z��aۭ��ڌ@E��_O�(4r�*Spܩ*&]+���)s^�cXQϐ�id�2����(U0�B�va��=�i�1y��\Z�&c�Li��*d"'@�<�`\�>�_|���� ���R���q���z�q�{R���6��еy\�Q�1�̑%��K+�N�ܼ��L_�?�=��}-zi,=�b��.[���b?'II:OI;��3߄�Kd�H �B���-g�xP�vD-[�羁����.Z���7��:�٥
b8q���3x��V��`��K����r�|�V�9��R�q ��WE�ґF0θs}��+^{a�F���%�o2}��ȣ`�5��5z+@D��0�N�~pK��Ao`T�R�AM ��k*��oF{�����,�T���m6Z�<�*��`gά5n��|&^60�3ʻ-I�2�7%��&�x�/�}�6��!D���K6��$B�g�9!l�U���Ed6e���87j�錈�i�^\�ڝJ&�I����O(�tc$gߵN���ئ�l�pu�.�*bH,�`�D��B�P�N:��Z2p�G̊:���r��on�*D����3݂v��擨�C,�DM3U��Ls���9�2�Q[9���/q_Zap3{Z��j��.����w����ɜ#���Wȫs�gHn�/�����iz����������Fq�E�s�.TQ%Cփ��D����!Ag��v5����Ą�hS��1��V�D��\ev[lU�ǈ.*h�+k�R[�Bw��,��:�ie(}���>"k���W���mq��~��6*C�^���W���v��I�|�R��;k�|��y��������MX��m�:�3�#JetiJ��O��G��z�C��s7�>��!��t��iW/�8��@����G즴a�����Qz����*�x�[�kx~USٟ!���2n�֖*4"��_����A��]Q1h��\�MV-4jJn��jR.+3ݵu}��KN��y[~U�vŸ��v�6Qv���]Ň��_Nb]y��!~)�<��y/7���VAqT��}VU>�����/����Mk��o�`��F�?� ��j���b_�)}�����#��d�-�����*����#W��D^���s[���~�����N\�3����G�����f����o}w�#�y�h����{�e�{�6�1�TS-:�e:|p�{�Xho���r2�4W����`}�OR<���`D��؋�}v�߳�?�L��٫����[pM��17����&������&���d�bN,�����_dK�C��`�0>ů��֨� R;K��ͧ�w����4l�,��t%e�ӽy)\������}s<�bp��~Y��?��y�9�����1FI'>���o��ϴ�  X��B�oVI���+l�ҷ���;z��!?�vL��G��'��F���tSL���9�����߁��^�L8�u�;y���R�?9�dR��t�B�sn>��7k�}{�{�pW���������1���Q����IH���P?��G%g*��r�d����ʽnu�gk���z��Yp�lƨ_��7릭��۝�Ĭ�%g����(��e��5m)"�d�WJ!�+E�s(�·xR�_S�5���wQ���Q�bJa�B���И�u<�[
"�n��9��\��[�7��>#15e�hm�b��v���(n�Q����x��4��e��<D�EUEቩx[5F9�e���ā���Au\`EQ��+.����_����)�����\�1'1S��Xwz6��3���-f'�?=�F�>�%�����n~�8���y��*>%G�V8\�*f�s�����1��qk�k;�n��6�G��k����6��w��:S'�4���lFw�	���۱W��Y9.�� ~��oIœw�	yF|t;;K�;���)t�jM�:hAp���G�=�P`�-(���/��E�{�}�*z��Ҟ�P�:��B�pr��&�����ɣ�'�n"�d���iB���טE�5����N�؁��-Y�����;�a��n�o�*N[��љX��>�y�MX7�$��w v��
�	������Z
ɜa??���<���ʦi�y�bAaHu��Rj�YI��J�EC�ǀ���ܼU��>4&;8����ޖ�w9_�L�!�&8H�����1�$b���h�G�.�?��&��\l�zq�����T���iH������o�#U�2I�b�ѥ�.�b��\I\����������J}y�0��s6x��}r<�=BL�r���]Y!����=�\'<?@xޞ�ǧ�ȗ�Mfε\��9�'��KJ�u'��C%@W�!���:qJ@�Tz�wN.�L޿� Y���V�
\��{Ԗ��Qr�K�=3o���f�ef�=`��>�l9�
a��C�E˂��-p���G"���Q*i�[νc����[~�E���W��5v����&�k����k�b4�)�ʣ��w'��X�������e�9�R�<=[�����	��ݾQ
��>w��ԣJ���e��;rtB����pq�����x�Ym�me�b 9;�n�	�滿 ��Kr�h�����`#�|C*�Q�]���+@����Kt���DUGU{
���[u�^�ܣt.��F�Q&�,��LUy�
5�Q�6��!�z�A�BK�=���IۆL��N�8� g�_�w?/q|��[�kgZd���o����(��_Juר4<��W/�0�-�3� 'rڝN��ˮv��,R�ׇ��C|B�x}⏞_�'G����>�r��?	���L��t$�X�wv��>��Rbq�����"��4�3�T��R�u��ӱM�|�=�l��$�
^p��H���z˿���x�B�e���{�B���o�d�Vh�)k��X*
�fؾ��.�D_�7J�O���**t�E�K�?]���avT����0���l{W���7u�B�����F}x9��c}�:w�����U��&(�TW;t ����N`�Z�gC7��ʣ�9����y{r�z���4�)���ʸ�;�Ya�Ϲ�ޗ
�;+�Í��lG�?��7��嬫(��6�4���	az��o�pXKH��iu�ד��פ��e1�潤�������5�d}"E"�z6D�7�����x������t��D��^2��y�^Nc���X](P���qd����"O��Z=O�_�OU@+rp]�㌷�X@Su�o2�����u�r�A��@0H�� Ɔ5}�[�2�Tn�dnl}2Y��9�뗱����.�WOĹ�e���㑻Ri��]�&��%��o%�Vau�-|�_�?<�kN�]=�'�B��q�2��Z&g{��se���ȂcɈ#l�Y�a�څ>�+��v��ma����3\�m�\�����D9����s0������HMj�u���XD���r��t��,�����|�,�����:�����1ݴ��7_����E�&#��^�bB�~q��n����(t�\S�Q�W�UO[��pw+��!lԗ��ܶ�5`A����Se�k��)O��l�V�`��x�ɭmĨ`�셭MOI�Rg^.��!��4�A�w���]eUJ}���.�x���k)��Q��GA|a~����R����޻��)�F�5a���U:�^EK�^�3���-JJ,��[�t��;U��I~o	7�X �[c���ѻ�WQ�6۬:��S]\�J��e�}�zLG����(�ܥ��*}b�)��h+_hd>
@��H��f	&�̹�c��!�G�(v�I/��|�Qa���n��V7m���dEx�^R୸��h��Z�\���R�9$/}�4��.j��hd�ҭ��bj��*��N���)`_'��3��hԢ=��.�
��c��M�X���Y�M1,��Ջ�>t_f���/�v���K��[�"W/p���V�8�B��wӮw���
+Q�;�\i�1�;k�������K� 4�波���]����(��c�����>N[��Np�=�ˈבt�xF>T<ƅ�O�`��ð��R����\�F��ga���('`qb��a����*�z�Y�*Q����Q��2&������꫒��V��xu0�ݫny�)�r��h������FH���]���]�4�[� �	�gۜ�T�[�Ky8M��v��߂]�>��0��[�HU�m�Մ�e7�B���#��ּ��E���^tBd��e�󭄈��P`G����I������b�BQ�g�|[ܰ�Ǚ)�X.	>�W�6b�����ڮ����q��[9���S|��@��Uř� �U�H�yD"s�ii��R�݇wA�G!�o\h�7�=�G)�}�;y�L��8��YVh,�%Jw�{��EƄ����X���.>�E@���fh8�U�S#/���בI�c����MDN��/�%��Y���[t~��%�h9yw>&Ŷ�Fd_��)T
�M+�V\�&�@7i@�L1O����5O�Ό�����:���[j�ǍÛE�Owdަ�5,ݤC��tL����)c��FģA�<GuRU�J���� 2��Qګ1�d/�����*�sRֲb�Vw���Q��(�/𽍣V�{�9Ȣ����d@w�ہ����1O��1XP8j���Wu�Œ���QNdBC��������u�f��]mF�Yyc���`.�S���4AӖWv6�m�;�n��߰1�ǫ5�ɗ�13m~*] #>:���hmY����R��4�Ϲ�{(���
��X�/����s9[lŌ��?��8�Gܓ�,��{�����kݫ�E[�һ�
�_Y��w\]$�)�VbG��\�b�M���nyl~#/��u%�(Q�#�Bjx�&��vQf�b�/���y�)�p�aP3�C�0�")�����;��eB�Qz�;Ύ��^�k �s��+�s��?԰�\���{m��
���v|7U�r��9���F1I���볳~K$����Ѽ�d:�	y��5�]K��R�	Ai8�������t�L)t>���N`$�#�KS/[1��0Z���i!%ݴ�r���p+.!�.�hG�o�mʷH�0���H?�R0���i����>}��Q+��-H�6�1���9P"������_̾F5�@T�N����ˆ�n��5�~�8�ux{�ܘ�������۶�b��H0j�u�x�|��e�������G��S.1)ި��I�ū8�z�P��\��o���&��T8���fY��M��f��=�U�Ex�A�]_�Q�����Kbp8�g�bM\'A+p,���q���8�F�A�W����7�DR'��줝��r:�E:�C5���ٮ��xJ��= $
_)���>
Z��Ѷe�/XT�a�u^�b;e�wdO{^}f���!�aM5�L����+�:g{����~�C��׬�/�}�M�+oMʚV&�h$��. dM"�BPa��~��'������m3���3�5K�(��'���d��6�����ebr^����xr$��[r8�_���3,�8�xĤ������-��O\����1Br���>�s�L`���A}��yS����"E��ILKI]l�6�E��h'r��~�2ttQ�����
E�Y�x�qmY��?�a���%9x��cO��(��(\�=w��Y���t���8���N
, �f
0+��s��itZ��}��m]{ľ;�z��z�w�@|ǅ�z����_�|8}ZgOo�;ж���.uJ-�9Mh�H�މf�Ӈ�FVR��ǩ��t�~X _ߐ���� ����M��n�÷ط�ang$��5��]�˫���W�tޱͩlRw�T�GG�di`[l��l۱�r��c�:5P[n1�K�G�,�0_�-0��F�z��	�T4�s����[̲���{�S%����+�;¢��&u�]��I"S�PZ�г9��N�]=z�]��؂u�p+s<�vRЅ����2��w���1�?J���*�������{��m�;+Xdk�}"L�&�Z��s��G���#�
Y��B����J�*;��lǆ#a�0}t���+�d�U�3A��g��V����xg�'m��b|�A�k�n���2�� ���/���ԥl�η�DYF�ۣG�(��4�FY0�($v�s�A:�g��;Ŏ����[������
��>'��@��+�/`tT����CR���&D[-,�\)�|u�\����e7lq�K��Y�V{/��=��8|�3��������.����P��^rvOߏh��Ca(�_ɪ�M�p��O�P�/���O�@�{j�z�a�pb���zP���\�"�#|�B�6��N�-�
%�)��|�֪��R���3��Y�����5�rR{�o���'�9<����W}� ��$�)��#��#��SO�k�V/�GcM�t�=�4�v�ށ@�L�G�%�K��x�E��"S�E�zܙ���q_�_�����g
Vw�M�(O�fT��p:����qJ�>�q�;���9deP��W~ %!9��������%���m��?\.)�5�/��hTS+?�ʓ������R5/s���;�T��t�7xf����lT���h�]+�c�r����ѬBk��5=,m�p�c]A
�ө��_Q�FNwn��k�%8�<������҄���Q�����z[R��ǋ�ӎ?CDJ�/��À=;��o���DJ���?�0CCq��0}n��$8���G���s�8�x��c��M�,�mӎ���:tt�;������4���N��.��#��:*ӊ?�=�LS+�wfE�13�0m����^B�����$�z�$�6v�F�-�D��z����7��C�H R��l���R6i�;���鬜����O�w��[��}�	wd��k�֦��ԓ��^��^?Վ�8z�#Y-�v4�*�w)��2}^n�A؉񧯟�¸_�~�ö�d\�>_�sɌ�ɫ�_lr^����޹�Sug�����	����RX�O-�(U9[I�|׼v����J�ì�j���炞���!�D=�ƕ��+�j2 S
�VH^}#gZ>��S%�9܎�W���>��6[��@O*�����춊��`�T����Ě�r���[���5�e�]Eف, v	�����t#�[#�fVM������6�1�	\pS-�	C56�V�#^u��{\v.p��Q`$�1<�sh�A�0�@d��:+E*��eƈ`Z��^��$�&��M�'k�{{$�>������,p�%�h�qڊ���<;ۊc|���8�N��2�FF!�xH��l>�L�Q9$9@�ٸ��S��{;��I��?�a�s��np-''}�;�Y<�~~t������ T`�|T���td4uy[pm*��Zr9g�g�d��O&;����/.���g{
����p����^��+��/v�DɤZ~���G�[]_����z@�i�wRF6L�)�ܫ-u��Ҳ��-?�w��ξe��z�Պ(�8�3q�bs��m���cd4!b�axvdW������6���L�!mm���Z��`���o̶Bxs�;�8��J��w23q��t^$֫��G�y��U,p�1e��"�X��(Zx�j���E�(�CnD���N��ę���-�	YvGUZ�HR�Q��Q<�}�M袀�3vWJ�S��T�ң�1���c��o��h�$"�]�N�sH��!Rx�Ng����=�L�N���"8��I�w�C�Ww ���D��|X �}�(�їP��ܓ�X�8V'Q&B��d���M��Y��4u	�K묽1�)��L��U���R0��V����)Q& :���1�cφsB�`�D�j�F�nQ�^�ۭ�c`p���x�l2���:���
�Bx Fd��z������s�T��๱�O��>�Y	����dq)�lI������H8�L��Bg�n��ؾGף�HaB��x1R��B],��=;*6C�ZL�R���'�8r�)���d��0K���{�Jn��5<27�!Կ���>�}%ꠀ��
T�o���o�k�Y���|�C�fҖs��U���O�fG0H�E��lG�8ݦ+�3�7l-�`Ҟ�Xb������\A�����������iǄ|����¥h��ImUՋ4x��W�\�~Be�#+�Mڛ39��:�~�,�H�����y�w�k�W�����,��YӆicS�ᤣU<L�u�yUA��?"纠���7�ة��iR�h�����.�4����Ch4��ҡW�7s��"��T;�Úx"��J���l�F'<�1}ُ/(@�=���6�T�j�����6C��%�D<��e47_�X�������19Ӄ����Н��V�A�$f�u2*�T�8������XT,���m��|�/�M�0!͉N<�@���2t)�5[�!u�e����bp�X���{ƪ���ƾT���{0K;�;"%=C��J��J�zj;s2Lj��c�A��6$H-�+U��6^�"Z!1إ�-���i$�����+,��[#	�;|�x0蜓��{��.���|��]�ivI�^���������P��`��Jz��ll�]�HJޗ���$]�Ǟ�*�W��Ʋ��} ��Ș���z᜔*=�a��m����ά�����J��0��}_�5RX���/��U��O\��⽊�c���&d~B��B�p���v�-���p��e�q��:�Lt�.�m�����D�]�sv���7��[��!S�Q�a
�N9q�v��!;�ʎ�uI٬V]cXr�3����Rw���f;b�.�׿>E�����N�F�C Λ*��11p ��ș$~l�V�v�-���H�
����Sl���юg_>)�~��`a|~qJI.K�K!=������;"?���xV^kT��؈�ݜY�5�;[�8�a]:�㢶��� _�����JS��gb�eH�o��=�5�g<w| ���cםyMg� bE�;S�}2��\j-Z��"������U��?7u������+J����o**�-w~�f;�l��	���[=��I}�����X���3���~i��E$��X~���7��!�# ��j){�u���sX���%�!\ӧ2�|�F~�3�n�4��v	�("on��&�p�y�&�3�Ű
G����@[�7e��v����/����y8�\.�̥���Z\�ZX�ZD��8�Ck7I�Tc�MU��HN��GP&8���t�=���'�*x.]�4�:
.�2h��G�\V�P�T&�n��F���wb��><�zK$[wn������9N#R4�S�og���R�1�S�����} {�)��BT{iF�F����?��'4�Y1]T���*7O>l�QX��ػ�S
�03^PwB�������k�V��I�� ����X}�.�t�$*^�}�'Gv~�䄤���5�RE�R:���������1�
DO,5�����8���#��B�<�lP[L��5O�o�Q�C� �ƭ���kiCMg������L��vV��=�a�Dt�$m��w���'k�6ϸ����֔�Xa���K5uOB���ϚH)i^L{Z ��qiZ�C{'��}-�L�� =�w��?s���v�K'b��pq�V�z<�K�OX�7�@�.�ݾ����|��g�,nl�nz��O�x�T��z����R��P�P�20M���"(��KZ��A|I����F�Uhg��c�=��S.R>ߑK�W�
-���jB���tV�F��]�����06�rs�,�4�� ���Q*�"�ð�����&۷}ii	IEJAB��!  �"--c��)�)���T�F��F��������������<��8�nV�:^0�ɵ�Ts~& I�K�R�]�أ��x ��А�:� o�~��uQ�{y�Q�tda�H�l�ɺɐ4l`���,"��FQ�%M��O��Z����, Q,�M���;�1�} 9�vlXA>
�1����9w�gD1'P��w|tk�I��F��+-\�˽����������.�Mg"�c	,*wW�3�h6qF�Ye���+�(��G�k#?�)l��
y �	ٙ,�<UOX������k~pB�f]& &sM}�	rZM[�ge���F���	�U�$	,�c*���"�u�~D�e��%}�P���N�k���ɬO4���s6�����TçC��%
������zCk&���Qյ����y��B��l P���_��5�a�7��+|�IE�`�ÇS3,h(�JP��u���B�_��^9.]�?4딊nߒyד�&ڸ4���NGN6���l0�=K��.Vr�u��_ֺr��C,�f�;���'Z�2�RbIP��},�ꑤ^��X���S�Nx=t�����C�/�*(�K���t�dX�5w�m�qQw�Z� �n�̭ͫ�"�qH�|��l-x�q�;Y}�|�}ث�&����<�_� �	r�Z9�����,|JY����^���G��\c:��?+-�����9<j|xז�N���`_��5�4Fpу�ۃe�y��l����ߨ�F�;�tfD��|�Jri������w_��>�A�]�V�љ1��H0'|��4���b/�ok�ؔ�Rֺ�?���K2jx�e��У�՚�4ҫg����g@���l�O�^4�텩\3�7�����N�'�9�����O��`�ZqT�[@�K1?�t�8�&��=���<���G���8�
,��T��c��`Sԥq����:�<�޽���#C��]h���em����a���q���@q�J��%�e��D�6-�UkkW��`ZU��?G"b^��*��ڤ�Ds:���L���w�&{�v�j��@<��T��,N����R>|�\�����$+�#�c���0��ǧ����7���q�In��{�k �?reT�®wƲ��zx�Ԏ5�Z�O�\y��:����g�[V,{�(N_)v�@���ya��VŌ4��DS.�;I�	 ���	i�������S)�YJ9^-��X�T���=�*�����J��q�YYK0;}��+Q7:�2b`]�В?C����0�|��)�|�}���Ns��]��YR��R�w7e�}��Ѻ
��0<X�f6��tͯ(Y�>ʴ+�������x�e�;$C"��Z�#�]L?_��hu�f��!c��Oi�Ӓ����W*�����n��w�R�ߒ�[W�G�6ܐ�|�\:������?�cs��i%y��z�����W�o�j�&����O$k([Z�O��w���������`f���rg��Y ��Q���QT���F�y��f�Sn6�(Il�`����Je��8�
�ݛe_�[��R���CG�F}S�3@��GF!�#��L\=��������z�l�fyr~鲱��o�Ӭ+y�@d<�}�gm�H\OC6Fe[�x�@�ʭ|�$�浝���l�lW�������";ֳ��)���[��p�}���"o���ҭg�bM9Ae>څ���gz=���t:Χ;�� 3�Lm��\��1�>�Fl;k����ېS��?�Ҕ��L�P�l�IF� (���|[=���-�D�I��E�_Y%���sG3���4&Tc	\�Bg�$�ӺÐ(3�'�e5�����g78e��_pQ\�E9�[��Z��>{ujq��O?�;Q+���xPO����[�@�R�0[`s��%�ʳ�gԚ#��L�?�3)�NL,��d�!3iY1�8e� ���X�>��Yw�,��?�~g"����\�ˣU,��7��@�9��+<y�FO��]�b���P�����bj_��7�
�Egׯ!�8.ܾ�bŤ�7^-�,�/~ufkt��Ʌɴd��mX�=���&�nvL�]?�A:%�ƥ��,Q�ϥm,�c惖k�B���|TW$9�����_���NiF~���O���i*^��5�����/����C�D�$�wk[����6n����D�ϴ�r�� 8李�o��u�
��i9"�G�7;���o!}�-�?�G?�\��g�X�Q�u�3�DԂ�W[���}X�k�tv���h������rJ�����]��L�ڧ�M��:�ҰW#��ɀ���x;+�,�X�#�_��_?&��1�  ^Yo��
�_Y[����=�����lX�#Re��@m+�ގ�/�y����E�x$W���7<�RU��%�&���y �j�2����� �,�>���M�r��8���2yB&��,6���|�R?���x}�L��T�3c���I�2�ye1Ҭ��ї�M��s�4�ּ�a�]����/ѣ���訨T��6���c"oa��C��f�,��h��� pp�$��8�;w
�*OX/��\vkko��'ߎ*�]dZ$=�&�����yޞM��GX�䤒`�5��\;Hޕh������*�Y�?��^	�	3�MOz=�=���*�l�4/�E �AaX��-d\�k:QBF�͛�?i���/��s��_�Ar�N� M .jzU�8��ʏnԤ�"�G$�9|��|l��:>r����%-�k���Y ���`t��KMm���~�=84��Y��O������P{�b��"3����O22�ml�;4y�ꊦ�;bے��ߍ<X����^�s��f�Z~�1�����c��A���6��5et�w[~�����~���׳<Fۆj�]�:��N^���;��߄ضS�;:�Ʌ�	]r	���Nt;pRc�Z��oIɇ�X\��~p�z٠l��,�ip��<�Zz�����KP߭*�uȕ�������z��'}�JU����>��.� �U�Iy�k>]@�IS��~]s�(���g?L^�J���<�0S4iͻ��Fێb�
�ޭl?c�38;u/
�(J�1���n��O+�����G�B)5C})u�qj`�L*�P�rF��{��x�Wr��*�9?����}�;vӅ��$$���(,E�w������~ا�$w����?'])Z�U�Y��LkW=2����ޮ;�e+jV���q���/PY����S�l5���6Z#T�q�J^Z���4^�]^~j����B"3������O�4�ͰKm����1�~��P��ó�x{�����z��Y?N���`���P��ݿ[����ߊ�ډ;��]��%��}
��~?X;��a�;�uT��塀����}����ebp��N���G2��I7=�^�!W��gB��+VňV�ɯ�1�|���?�	̕R:	���X?�[�t�nl�eiN��	dd�ۃY���*����q`��E�3��Uf�� B�.ߺB��_=��;��Ԇ/_
�j32ķ3̛�f8�v/:�Q�t�}vBUe�2���v����V�&����9�����. ]O�k���mw*�Η���IU�&0����C�����OM�y�g͛���WY[��(~����']E�>qa��'��2m��F�SS�/Ь����Ш2�*}n��z��[��Ip�Z��"�c��@�,}O� b�0ِ��C��ã�F�� F/z�X�rL(�4��١G�����̒���/"��q0����zب�6�&�hB�_f`��ӧ	��e��#ѥF�9���� M{K����h���ζ���<�4v���J�5�|��*���6��}����+�5����|�mf���z�r���������[ڟTcLR���ƚ ?�af�m�қȤ}7/�o��	�����/���]\p4��o$��������$���}��Y���Ύ��1�F�4���Vl&&�ap�*����S�Y^�@�U/(v�%�)��A����ی��U���<Wx?��1C"a|��<�n�r�� �X�F�[�b�u�V��_��-���Fų�9`֚�,�îj,��j��x6<�|s���{�M ��⤿匞����}�6c*��`1L�nv�"�Um�.�L<� ��hM]�m}4�����eh�4�/݅�gm��˛0=)/š�͈vG{6�a��ie]A�L��iT&��wf�zdM�[v��|7)A�A�W�GV
��m�
�kvm��y��[�\W�5=�%�"��xrDy� D=�9�ב�i��ݸ>�dJ6�:H�7V*Mաhq�����v��n�z1�7�^	q1 �k�_�ҕ��I27�*9כ��:��qְi�`,�箄6�Cz�K�#>��C��(r�*��W������Q�E*ܑ{w����5�m#��l��"�C {�L$¢�Jf�+Q�?�ܑ\$����W<h������[�����a��!�������(/�&���_k�k���i�v��`�J�T��H^�t�<�+��a�H L�	�A��J-��ӄwar����(�q���]��&E��U����D|���89)�I�2�~�v�y��\<��_��5��n�[��9bB���彿`�Mn��ׯl����� ����lp�߶ɷz���|���7R=�B'y����fq��^�1t�
�)j�V��I(d�9���$5��ː�+��
��i��6"�����T����u����\�>��l��Ȃb��#�%���$�WW޺���\M]򰻷�͉J#�J�d�����\�����E�Q��v��.�W����y�7����2o8���p�x������:D�_� ��!�����w�n"����M�껓n*�k�|��kð,ЬQJ7���|�����O;�B��z�7�r���,Sr=���Ն�4�ՕOϝу{35 �#��6�뤔�Xw��/Z=�Cu-��7���������"��?��������B�Td��v������۴�׫V�S`!�` _�v~�U�\��pyYpF���(l�����`�>:���߳��k�����^s;`�:�>e�Gɛ����/my����_��|f�3,����k,�y>�n9>����U�]݈�X�f�X�1��T%�HX,��>�+g��$����>�6^�#n���"�c�����m�j��cmB�b��E;�t�}���©�_�E�y���Ml;�^���o�3p��+�xµ����ћ���'Y/Y����+\�+���F�8��Z�ޡ�H��B����Qw� ��	55u7��jѮ���4���������D_z�c�-ġ9JW�K��|Hdg����{2F0&�)�\��'&�&C��M���;c��Hg(FE�3��#p�<�嗯���b��6�)R9�/�`4\Ս��a��ğ���Y�ǎ�?R\��&2h~ﶔ$㵛D������p�*m�P��_���"_�Q@]O/��ծ�$�Y�%����yN�0\~~RR~�i8q��{��i�:�F׏P	\K�Ϻ���M=Nnҝ:��ޑqf?������D�{����&���R� o-�ln��+�ƧT�^rՃ�cZ��f���-甛'�d)����͙����3��K���u��?��3D��Ͼ�����+�#YӉ��A7�v����Z3����9�a�&���]�oI�_���� PA��0(X,eD�����+i���� y���I�f�1��5��2������ ��@�oG���#�W���D�o6��0�ν|�;�������a���1��ٚa����k���w�3���~V�d=� NIn�uS�y��>��\�;����o$�IxJ�."�ODgH2�@1d�-+e��Y1���8�h+�\��=�:y��޷���G��V֖�Gǋ�qQ��i�+�(��N��R���1_�����(+��ֺeK�'�pUmmNm����t���%�W��U����tn��Ug� �gdy_��Ӟ����q��e���!fq�G~7��T����x]���/W5�8��l���"r����L97�l6�L��	ʭj�&�Z�{�u	��.)�!P��݁�l�6�A���+L��ٟ[%V��\ؐ�L�ϵւ֬��n�,��<T�}2� ^�^|�!��]LQfQ��}ݽjzm=�U�@B��F���v\����dO�bB�	�ё�{k#��!�<���64�}^v�ǜ�[��{zJ�2��Q�􇏓�Gh�������7�q_ ��#Yv�w�R7֝?���/��|_>n60o�����:'m������5|��0��:L����q7;s�?{�v��:R��y��#���i]�U�"���!5�����q��V�沦��j���kq2PM5���+��{=u��3���h�)��Ȯ��
B�[��Y�}I���@_�������̟�A9�/߱L���'\���m�ζ1��)�͸^�m���?�H	�l�ƿ��S!��(ptW �e�|����|AA�2�H�w�R��.)�V��S��ɥ���"�_ߋ���_`�H�V�-��w�ԩ�Q,WY����1"-A�,_�qoT+8e>�Qw*N=�a�ʬ�ҋ���"��Ou���"�J�F��Qc��xsz�_����
�E!Ќc���ɢl������y꾈�Jt���ES5�o*~�Ω�mq��C�}~5{��y�ڹc�ݘ��(N�x��mF�ۥc~�Dt����8�����9�A�1�k8�M�y����cd�UǍuP`s����vO4�h{�X�!ׇ�'�=W��]T�T�b�_�l��hɀIE�O��0	d���)�	�'rO�����>p#F���ӫ��\��ʌ���z� Zt��Κ| �dR�����=q�� TU�Y��jk7��F��w���%�U�T�\T�ՠ��pץ�"�H
�Qb�73�W0Aa��ɑ�g;�E�?�94w�r���.![7���81ݜ��y�;D^��@1D�qSD��;y�P���A b�e��z^ѹ�9�AJ��4��jm��Ӽ��s�}�X�/��6w�1u6��3�-��������:�hj[��8#ӥ2r��E�G�;_�:n�v5�Y�ב"xI�"Qڊ
���� �=Wܬ��|�פ���G��:�C�W�|�/B�d�
��l���n��E�S_dL�E-�L~�h���,�����A�p`kzM	�=�q��89�m͡��݊��1��j��2�����,�����7��E r�տ�������s&Q�;�O�0]�n�c����q�LL�,�NUV���{إ����V�_��ZE�a>�8�5��8ͯ9�D�G��2l!(-�Ё�T{j�V@h��Zdd�	"��+�z����h���ac��;��Q�O�Mza:b�u�@�:N/�c�ne��,#ƖB���C��H c��S��H!�8R��o�	h�Ao�5��J�z3��~G��~�*U�3����nv(k^ow�̄��/���_��ˏ���q���ǵb�ٻ<��A���F�6Zc}+ߔ�f�z��`D�E�39�hԓ`��ܹ�N�t�u�7��d~&��R�}*տ9J����-_���6���5�l�;7��XI�t���.�^��ѡ�JXj�/����m��@}�1�<d�X{"%8���rz���)"�ʙMt͞F���H듉��t"�1�{0��w����s{
�T�E�"f±S��DNt�V�M�X}L���Ͻ��.���<0T�����l��~ILH���� �TdEq߾����Ddo��ޫoceGb.�`�`0Hp�0��*D��"r�fZ2+�h�u�ୟ�}B�"��CN���ˀ#!J9����^���W��O�61�"{DX�	t����+yɀ�h��V���h�{Z����AM{ϫ/��=@�ay��0=(M-i�<���k�zR��_�%��U�F��w���]�{K3xE��*z��˰rØ���UT#��!�7�/���ڜ�s=i��%�K( Ȩ�=eQ�؏���/E�ҳ���7����J�8�C��<��w@�C���ߴ{=����g�	���g�2<�����j���~Nr�Q��2�zů��`.���]�Q�l�ц���X��	�G�>���دz��O��b�n���ר+Wna�]���rv��'m+K*2­�JxU�'ș�,A�)�Ҙ���8L���FI�ʚ&2q���k��e�X�due��	ud��G�P�\llx�{�Ō����$�z㣫a�֊��s��ɽ�z>��!�����;-��v~ƌ�5n>�A��#+�ס��c��<���y�Ql�%4O0R)L#���1m����p��[ېڸ��SGZ�̼�;��QJiq0�{�{t��m��ki���z	�_>_�k@�X*R>?p�;��}�� F����aVXP �H��z$a �B�ňyi)j�z|��ϩg��ؖ����p륝3�dߥO�8�܆���>L*�z*VUX�SR�%���d��쬣x�u�VY�	ɣ����A��^$��c5'���U�ܒ�6N����z��G�m�u,�碵:��V����2�4%�#Պ?�d�"�L0h5ߜf�%kd@��^<������奸�Ờ-����T�����ۈ��XZOw
{:#1x��^	_�$��FK�6��=CZP:�7L��>�g�
o��'�׿���1����ɫ��2ƙ`:�=��H�<�XG���>P��h�<��hU�8^��P���3r����2��{��T��;SElm�l(��#� �@g���לn~�c������櫡��V�r!G��Ce����]����%u�0��x��&��s���w�e�lOUj�yø���FQW�ǷDS��_���r�;�5��QU&_�6�p�IU����Y���T���2���:��mgw�a�JL�=a���c�����ѷ&��T��������>����ؙ��'�#􂫼z��C6���j�:�u�$��:��t{�j(Y��c�wJl�ךB:β;0:tX�Z;Î�f�9�Cy,-��3�����*�y�Y���Ɉ|���|UQ��f��\z�z��&�����jģ
ʛ��ȩ��7ϴ
�QZi��k���),��(�
#�mJ_mx�7�ƫ���S�����)i'ڤ6��#X��,mx�w7~�1���l�5x���漗��=��Z/@����}T?d�;����J�-����^�'�?�?<�R�f8�ǾC�-=���D�e�8�����X�)ș�2SЈ��I\}F,lU���~P���	6v���G9Yk@��?/�+�]����8qR��?Kx����8�{Q��߂.��^�PQQ�s��Cbޕj���G�t�	:��zK�,G�P%����� �Y��]����!�?�ȁ'����a�MpHe��H��k�Nd���@�+���G���7������!-M�_����s��1����b�4��(�!�Z�_n��X'� ���~���һ�f:ǖ������i��Os����!���#�>T���k�0�P��Ra()y	1��'i��a��t�n=�[����������gͥ�oݟ��B�0����A�[�0NL��U4zx�@%�l�E�WT�W����v��S�L1;@��$x���i]��}c�N@�="�b����{E��蕃����=m=
���K}��X�g�Җ�6�;ƞ~��^��+(d�O�����닳}���6OP-�2b�2�ҵ+z�Ȁ�:�l��`+K�"��߉��l��b�	�c���-�uF��'M����X����L��s�o��й�
�.�_��C�=��מ]��g�#�#���\���ي%����K4�*>�e*m3_���9�ޅL6�E	�ba�K[[���:����􃢨��������߽ɸ(���\����ޗ�&��:q�z�D=@����%�QD�T�yk`<�f8:0�
~�(���������>0r�tG��rX8�h$y��I�Ou�S�� �8�������*�U�@�5�_�X�$N���[��Fļ;�z"x���G�#�p
MK�̰���Yb0��;|�F��dMĂ�F��K�ڟ�O�fE��i=&ٴ�������s����ʩ�e^չ�]q
o���u�f����]�bu���f_��S'.X�t����9����**P+�F9&p|?�RQj<���S���(� ٸ��ϟ9�9y��C��4w��XY��F�ߕ��� ��X)��4���Ы>^>�"���TF��#<����.ٛ.�:L�fRo��c��8��'ġtB:��<�Y�oWL�{�t.��p�=#��L�@~ �t�c����3X+ړ����Q�l���8��L��}�@��_&秒o�TP��X ���m���L��NGmJqm4R�5K� �S��N�3DJ���n�P�h�6�5�m�p�Z���cꔥ�c�����y~��q�v����>J��9�@���kM�����k�݅�X:�?e6��a���o囱x~��#��RE�F&�<r��k���H�ls��.����!k%�h�='`�B����;�h+���s�l�Z�Ş�Ĺ�+��jȟ�9���`��Ł^Ƙ�۫pQ�#�%u)�>q�%��9��D�9�f8'���M�MD�<�:ۭ����$�.-�u�Ap�ݤ+[�`J⛧��*��}F��eD�ëf�uo ^��9`���öa��gt�a�]w�n�;>����N�׳�6|���}Z>�pC[�&��]l��eX���4e��&N"��3G��_l��l�1�ew�ŕ�*6)P|�}<v��$�|���o�{�Qj^�������gd��+�[��jf�)3��l3}3Ç�f�P���A����u��%�KX�2a�ϊ��q�<�'@�F�l '�����v�Cm(��n>z��;@�fa������O��*�Q�_Ԇ���b�9�:�t��!�1li�Nhl���iy����n��8�L��.m���e@�Q��w�:�eṏ�{�\=F�hO����ؐ���y>lFy �?����L}���/w��wJ-�"_k��7(����U��ʇ=jw����H�ei��J��K�G�+�r�k��X�4%o,Ĳ,�C������χ?��d����
@���9��Y�POSfƖ������;����fTc�ǚ������*��p��,��=i\�s�<u�T�Db(��|0�me�|f}�̒���y��ˣYŸ����i��Z���:SU��S��Z�j�ۜM���X���F�S��B� <xEA�D��\	:��nO��{Z��3"��B��6I�-�>��n�yrS�m���{j$ɬ�F����}���aN�e���I��ƍK��iK��͉�ȭ�P�U֟n�cnG�I�cՏ��X�:�rC�zR��OJ�;G~�N�u��ʞ�2k� )�l4����uT����sQ@W�rI
�T�(�j|F��%*�%�u�a�ٞ�_��"��N�����.1P�EY��:�⊈/O������I��
�9H��0�gW쥫Y��)zH�Љ��}ڴ�+_��82!�T�[8�6�cd���wG���6����D;�#:@�����k� ���T+o�a���o��a��O�~4IՇ�?r�s[p{eFW��1�ִ�1��\��O�4���f��vW&�g��<ұ��/�iJ�IJf4O��B���$�tP׹_~?r�@;k@��zd���R��m�G������c����m;�����f��z��~4�~ǧIuc�A��<��C�/��}�!�O-����޺�|XǤ��AZ'2��VO-n�F�n�b�4��\}Q���Q|j`�"x'�q����6�����i���4?Uq TٽpF���X��2¬�H�j-�v�`���q���n7s%���$��8�/�d��%{go
���='\�Ey�*�?��3��ϛS�_��D��ڶ�� �p��j#v�6�����,�W#}�,%]��s=-2�x��?���E��Ba�9�GH�w�6������A�Wp?P���ߙ��tG��?
����'���WJ��1MwaQa��@�����v�(�����d1.�.k����o%����@�C�g4�X��� �ѫ�����م���ug�̝���=��[m���$�����m���d���t��w{��<�\NJb��o���?��'���J~�dt� �0Ǹ�tg��Y��2��Y�.��9���]�41A{�v{�B )F���K�>9@�v>9mS[�W���#�9�����98/=j�t�����ح%���Tn��m����`Y�hCn@��'�-r���W���B)1?Dd'�F48�,�ë��.&�Až�-=-��o��� 	�YV+i|ˉ��)гL�U~)2�^F�5P���{����~�i\��Z���-*ֱ�W`a��Ie�=�+�n��?����q---����Crr�g�4g�����s�\`Ŀ-E|}��o��s�K�E�0����]@x�4���?a�V��&�3Wϋ����슈l�8���LU���2x���I�M����ډS�[����7иk�iGk��F~C�7 �����(�T0��Ѻט�ǯ��Nu%�=a0��*��O��Nw&+h�s��*X�M��.]���+�T�b ��V����z�u��~MG���'0�Έ9���	��g Nf���l��8�78��
1���y[^����S��˴z�(8��OĻ����a�iz�~�b`���3�@n(s��n8���E҃��p���Xp{)� w!x0!c�Ot���X�.���HZ��z�O&?�t9��O�z��
�Qb���;�����R�.�{R*o�K��AO��-UZ��o��B��Z�%"�~$��E*����K$|�)[�����=_�g9�E�}M�iBN�Q�{�k3��{�����i��Jt�aR��kU��|t5��ܫ%N�}�(>KלS��ٙ| �O^�Kt��w{�a��vq�V!$mz�e�Z��IT��c��:r�}���p�g�0"5�ޒ�R��k�����Q7��׍`��_�Y��sί5�$♜��D��5I���<l��j�k-��sM��5����Z&\��< ��X�
�j5b���,S9�mw�m�3�'���p��j����a��a�H�ޱ��Nu6���]���� ��}z���-��q�T�tL�*}g`���E��zSƯ<���gFѽi��	�v�p�گ�m�i�~��å�e�ɤ��5����/�ފu]�^E�-M%�&��J5X��q0���uKPF����	��-e��l\�HkMN���#�YD��S!�`�Q&UبY~��0���U�����d���W#Cz5(���s���U�e�Z���ׇ�<dUͭ->��U;*b��K�ݍă�s2X�T��x����FG���@-W�nP�b~��a��b�F�E�P�竀�L���ˤ�������&[�2���믬���|�lw��֙/+�j�K�N��]Z+M���Z`"WqEV�Q1e���j�:]��oByѧ�{����hS��ϩ�^pd�6�Ǘ>��$���.1��4����X��j;��ӪK@�9��P�g�g�z)��+�B9����1���Q��M��wS�ٖ��PRԕ������o�'G�0����}���$�Z���W.@�ˬ!+�����|��g%��
�>��1��3��K���,�=b���e˳��M��@�f��	�X�k�`Vnk���[���	�d�ɣz�xXb��ASqS'өB�H�l�Y���3���I�a�{�h�в������]�>f������ �>FdPu�� n�К�W��`	�w�7c�@簎�"��9V��?A��_v.@r�}��vG�4Sn�0郦���5����f��ٰ�GW����~�`j	>�h?&௾b:�����t��O��Wu�/i�S��[E0rsU���F�<���1�"�9�MCKw��|h.�*���c�����6-~�n����3�l�	�wK��;�ꜵ�+�l���1��� ���-+J����6��}>��W��ݪ)J������l��>@u��L'J�_�(s=�E	���]>Ŧ%�>�S0خU>�-eg����@��W����2B~��Ϟ��a5)�d���{®G��˒4o�.z1�d�6��)�G~��jd��&SJs- ���	��R|�D�������o�L'f�����<��Ң�no��[�<������ _nPQøV���%�=�2��Ck^�G�/-͈ͬ��c�R��PUX���OX��e]XX�8Om�Oq�-�8�ٷ�4�-���њ���r!��xQŏ;p����9<�a�ӳc} _�ϡhX���1փ/z+d�����G$M�������p'���'ߗ��9`��|+� |^��D�|���Z1���+1t��g�	���x��s����#��X�!�ݓ-�h��?�"�x�Ne�Y�~����# �>[9�8�/�H��=;r]��i���ŁX�^z�7M�	��x,��G�-�-�.����J2��:%o�ҥge��>�Us��I�v�9��NZ1x��?8�!�%����̽njiaS�-�W�]U�N�z��nA!�mqv��eb��| -��ŚGE�6%I�N����0���O--v�j�!�4����<[�>��aN�;�+��s����@�I�v��O������"����:��1lhci|���.�Mm+�r_Ŵ"�[�-�%_���o"�!x��*�y�+�b�f�x��D��6LE�io-��Z��}v2�2��~o�5Y��"�ӝj��Yft�2ضZ���^��bn=�tp�P�I`�^B�~�4���v!�8�IQ������=@T2�=iς�n��q���^?��+�W����̨�!ӣ�M��e��o$��&��=S�{-'��f�y���m�g�/�����m��f��~Yl��T���&��F9B	f#���`Ii[�Fo���xc�{E�O��K��}�[��k�q���� �}��L8
��'�q]�CI�J�F�K�t'���U+i���:���9%Ă:���%�m��z�nY+��̃Jc�|��[5��F�kV�GNH������=�����hV'�u>P\!��lA�y(d<��2���q��4'�Fb��6����1�p�ݏ{a؏]*Ckr^�8�����Oȸ_���j��I(�6�ݢ���E}wIm�O�	ϴ/��H�����`c@ߕ�C t�m}����A�M�wkF&6�λ9�{���n
�����2�n��e��X0N*�"s����� ��dߥ�����W�j��F���e�.��U�)�;�0zl���A�z_-�&�K!�appcA"1���c���M����yg�� ֻ�'M�����~�}�to���Ā~�Q��N�-I�2 +���]��z���%�.�p#�2փ��Ӿ��3HJh 4���X����x�w޶=��٥��dd��G�.8��P�<l恇����K����j� oM��	���GW7;@�S�*�{��Q���:\6�cUa�̈�Oa���m#R��{#��$=m˞/Rtg�B)�6�9Q����K$$]k�m�3c���0�<��K�T�#�HLlm1&�'�0�g�
��g�_�Y�C�I���v��B���������l&�:�����G~�0/qD�lI��O7��u�L��n/�M����?Z��D��E}���O���J$=�5���rBs��-�
޷�
VS:��˳��a�&M}8��^mE���_Y�n����8p'�!�G�Y�3���i&�G+�y�~�E°����N36�U7����H>K����U;Y���gRU��v��f,+
W�7��ST-P��3��p2O���2���:�OOW���C1�\�V�6�7n'99�����W9`ת���j��:!j?,(�F�H��G�E��F��,@_�we(Ҟf����Bs�.��>��x*��HAZ�m�2�?�>��\(�������?��,OI0���N,w�����0�O�<���^L���J�y�zf�#$��/�;��#�m��[��&����7�Aw�r�t�?|��=�y�w�3dt&��2��K S4W���xD]�m6�yY�44��N���;�$|"
�h�#W ����3��j.��*�f�ړFP��	`����!j�F,}"+I�*ڲ^��5���9vGkfߝ�S�G+����VV�P;ٟ6��_8��`D�oHr<�Q�(žx~���WB�2�:�0e2V ^�D�|M�U�u�]Q�tD���6���zjT��^��~2�>Z��.�z��I����h��J����}~>�Yj������ٽ���l����P2�I��m���6��ٍ�!��U�C���H�Rח9y����O����n���Q�O���Qy3�g�-�vX>S�(��S����ej��h�T+n/�$R��������l����� 4�W�8��.ߠ�bVuDᤩ��ӆ׈|����T�/�;�)��M<F��F���~����qƄ^eĴ����21�3�g��l���[�7ŚR;�1{�HL�����3��mK�llןTW�A[(6n��~���O� �/4ڏάڶL��"�ooUU������H# !ҥ�t�p@��� )�!����<tHw7����<��^}���w��c8�g�5ל�Xk�B]�8�$F]ag�'�������1�i��B	���F��q�����b�2:���>���P��ߥ�w��>��\HW�$�[P���n���u\�HmL��^�=��oD?�Ju�l��&?s��DEX�P�E�[��!.N������c�bL&�����|�n3��S(F(m4�..��X�q�E�K�6����,j�G�(|;���|"���P��SX���_�$�Z�;Fc� ��n�}1|���?�<�rw�v�>����p^	T��V�Cֆ6���io�zct�r�}��DmK�b%c�$6+�yX����%j�=�œ��B�8����HW��a���v����W䥣��9��1�ݦ0R� ڟke�dY�vZ��|�>�u�X���W�@���Mw����L������-�>�	�|�
��Ĕb����2��1*�1�ޘ^+h���%:{�w�aD�J	}��)I��슋{<�}��2\�Q{j���h���)�����>��s��]t�h�Ŧt�I�P�v47p����s_S/�ʊo�d�
�<�D���^�^`f��&��8/r����{X;u�:����(?�4� ax`i��1� 	������[Pj�Y=��-T�~��^�������KP�B�&ǋ�|�E�ͽ�{��a[N�{�b�� 8�n�M˂d��;�t��i׃��N'Ϩ�_�b���6����{�md�t��칄D��^�جt���DC~��.@ ؚ�L��"v�kaq��P=RQ�R�xxD,�����:��z;�V�K�yo�t��"��)��+����QTa������XK�6��J�0�:��N�\��5B{��l3��J��|	C�v0ʙ����\��/R嚈Tu�;w(���Z2��q�8Ċ����<�H�f��B���64�OQNe�y���� Y�N�-�1WNW��$�x֋k��m���#��Qi���|�
&={�'��澨5�smc�&'��:쫇�Z�ߊ��}�X ��5����Ű�\"z�ҧ��x&���v/�zk���)��'�5��񘻸_K��;�ؿ1n���t�u�4��B���G�����zuu<J��_̓��0��`M��.t?pP*��c����h4��S�S��_�o�qL��Ú�1(cj"@i5�_�[�<�v/��3��y�]���=�>�}��x���MX_� <���֨d�Tv��M�k�#&���u;��� �Қp4�a��P�9���	��0���?q9�9�<V�����-�c����-�V-�{
���q�B)������Oo���+�*��������D����gmV�����S�Z�u�r2��|�H�^�&��C�V���E�<!�R޸�����}@~p���[dӵ9q�<r9��.���_�lܾ/��tq(5"aCڻ�p�U�{��Gxa����,)ЦcR�>�NƕGO�L�"-�-r��kw����[֏jD��Ӿz����Ntx�J�I}�D�0�:(�m��}�e��������7�p�`���r����;Z�ˠ�}�]C�>Wz�k|�k��Ưi���^:��Kp0!A�X�}���y[�����Lt��d(�������z���+�K�QJ�+P��K�"��Zw��������FZ�Ɉ�Q97�Ե:g=}�o���J�׳v����
�o`�R��.�+h�����3uH��~�ɏ���O��D��uHQ�7��s�d�;/Э���C/��Mks�u����[1,0��)�7|"����sw��y�:���r�1\��=���Fu�^�,grZ�`溌x���y����I��=��I$U���H���zlgb���.���߲�*�ݠ>�iC���[^�]����*���$Sw�Ͽ�ԭӽP��^�����4ţa���-*>���-���tp���Ð�[�@��.�w}G�i[.Dn��������P_��z��H��MWT�����c+��R������|�癇�1e �KGLkTtH@�i���\xz��2O�<ل�>v뙵�W(�cחBm�$�Ѓ!G��������q]7��%�i@��*~�߳����r:m�c��".Y@չL:�
��͓�5Q���Iw;�/!8��S ��CE���Y�Uv�u���jo\���yD��
�)L��lɌQ1Ab�T>����ȕ�f��9�#�V���\��O!?��l��=O���g23x��1��A'9n�m��`c{|��؇mE�`�<�[��I�Ѵ=taa ��։/o��_��1��S�M9�q|�2\P];�r���ӆ�.�C������m)-��+ق-fn���^o��޼��]��H��k�vK�A�?͂�@�2Sr��ծ�u�4�N��I�:E-r���H�-Ȱͣ]*�B�:_�k��7�.�w1m&�cH�X��|�kB�(�_ 6��F��pa�����o�V��$m��Ao��˂kPd��6"�)�hׅ�ͮ�`�:�$����b%�נ���_�!��bZMNO7'��t1�+j-�:gy�oM�#�69m�cf�tQbZa�,���z𙥓�g>�2C^��\�^�|lШ��~��� �µ�Kr�uӃ��& c���)w����+��f����+~���4qe$SQ�z�d�]U'��e{�hj��Z�~W&޹�;��7a8/v)�*���eɟ1�܀|ۜW�b��Z����mI����bۺ�}��@�-YE�?��I����=t����J`=����c�ʎ���m}��h����(�tV�Z[��unY����A5��OPz�J�\o��a�2�-M��
3-T��"w�0ĳZ�K��"�#(j�)4B*�Q����P�N]֬�����R5������z��R��ͫ>�d�ju�іuK�C��K�(�N�#��p@�I�R]�j0�q�v�}���(A�t[$�Og��s(�|��t
��U���/�{��tz��g1�����c��v&��8߼d.xʘ
mzku_F+�6kڞ�R�z�h��]8֭V�[V�텞�1Qc��!˟P���hi�x�<Q��B\P~Ѵ�5���$v�s�i��D��B�AjױY|_F_O�ժ/z	EۤJ��K�X�84p@h𓙋�g�!>�q8�=�M��ӆ[��OFm`ޝ�
m��P!~��8d�җ*�������	Ͻ���E���̽r���Ӣ�P�^�ܙ��Ud� ���]��<�-��:<��}Ԏ}�Y�#8~/|�s��=Q�_��,�8yner_��	���t#���y��j�W��M�V�l�}�����o-<mWL�3hX�����%��gˮ�lz��J�@T�"�B�.��1ʚm�ԝ?�T�Tu�8,��C�*����/
�z&�V�
�l��hQ��/��l O;u��l8軚�ϩ���,�rW�>U����d⭵:"�NKq;�v�E�/�Í�铁O����r�~�=Z� >�v���E�,հ��ض���zS5��
�sz�{Gi��;.w�b������Z��T�>��5bڱC�����r,���\����ՐY`A�yZ�I�ocݹ�Bc��4Qז>�3xk9|��w�/3|$��w\��G��i���؀r�qﱟ����,f�ȱ�����Ѷ�f�I��b�_$ݮ��ۉ{zI3	�dy䰿rs�<��\Xg%�%��Y����U?�R��������`)�'��UR*��gU�dw����t&u�G�[쏏 �3J��A��,ۃ�q�LN�yq����=z��89�����syz{���C�����aG	���K֊2�bV
^�utQ��>?F�"���w|�=�5��K�母}���$�Z�� Kӻ���Ѥ����a�D��kޟ���]�A��y(DB�	�?�����w_&i����iag#�`�;�8��k$L1�c(Ya������x��Vt^�됥�0��T+n�+Ȕ�u��#_�%j��r��Pc�f�m����K(�cSʹ�R�� +!���(�8�wS�r����k��ڣ�m��$�F��*b�<0� ��=\Q�4����F�:��D��-�O{� ���mx��=�Mt�7,��ah��B���>"�j�8�y�4�Y��� �C�af��^�Se�XR�h�@�3 l}�oV�;�'�3.Ь�.c�O����?��w�S�4pY��%/��|.�	����"n[���3�1O���<v]hb�qw�X����E�6�:a۶][�]���1-���u���?t�ߣϠ
�2,�m!�.�IU�]r�����c���"�p�r�d����,9VH�#���ny��䈠q˕A�l���®+ÃN�����]�~^|�����������[m|�� ���b��=XQ��ϣ��eN�~^�?��F�@���SS�|7��5؀�?<���>���� �ݛv��C~mC���Zt��R_(���_� ���h�A��v��UFScYPqp{���*Ao��9���k��B��/a,�5�$���J0ȏ�Apc_��6�i�%���T�Q���
P��ex��-�x.�]p�ԈS��?|v��0�|��8�7�*,	ց}�z����h�<1� ��/[X�82K^�ղ���e�۴��TsL&e����O~�ہ��~�R�"NT��m������3����3/B�a����Kn����{��f@Y��'[�ϡp�fK!U"Q��~��,q��փG`�Ov�{�"�p �x���K�"+;4,$�����i����tr���_13��/�|��و��at� �`P`FZJ=$e����;ܤ�_��i#DS`wK۷��@���R�ċ���9�0/�j��n��Vr�i����@�y��$�T����ӕ\��u���/7z�=?~A䚐��YiۀH�j�UC,%�U)�tA[�P�%#������s�7a3ywU���ox���U��GL�R���K�A����C�Nx��ԋ�ӏ��,B�L����/�� �=�3���{������v^��Sb�.��<���Nqu9���1]^�| ��k�kk=\�E�ԋ����&�*�b�tL�T:,G��1���?MY���ai��������$�߽k /�[zGŢ��d�O�qN��)|�;d���K� ��2T8ߞ�Y[C�r�,)������0'��,@�2.��Ӛ���ef�g��	��h�K����Z�uYbiS���Q��-�)~������L������g���� �7uN��ЅA�4���Ї��ZUO��{�%;�������`]��|�p%�œh7��L����l? �,��ǫ��|���Sٹ�k���x��<F-itf��xܑ7�]^���}�j��?������B� %o�=��{��se��OJ�~��L-�2�a3�"'�|w�yн�X"���ц�ڟ���?;�1z��}뇋�t|Q}��M��T���6Ÿ~[f��S3�H}�;s�8���7�����3.ΟF.��1M)#-H�4���K��HX	=�y��-a�R�O�e<��y%�������A?��J�=���ɧ\x�,򶓚^Y���vv%��7��j�0r�����D��QE�ui+�8M3I�v�Z�J��-�Wjj�^p5O����W'q�`/X�Y�%[_HU���d'���ru�.F�N�L��p3�2���(���Ĭ'�|;�3*i�BL=��9���O1�x����"�)?m#��;���i�C��$�mx U��k�\?d��Ցٸ�_�4��{��
�����x�B�K�zå����ơ�q矵`������u{��v\!��:[�����z��l���;!�F�mI}�lH�~��wR�h)w����8r,���{������_��n���+79�~lQ��0��x����=Q`;cR�Kj=�ٚ�2�x_�pc��x
�]Ř�	�E�ě�	Ɉ�&����?F��3��7�ỷx
mN ܜ������u�dDBZ<������XnF�я�$�D��&"�����)��h�1wjUs�7p�#<�XW��9��O�h���=v3��M�rU��'hѶ?��B^M�<1'�!+A����LM��ʿ������D��:���{��כ'A�ϯCE���e�
�˿C?����=�#6�?��_G'��gC���[puS7yD:*�^�Pnx�*Nj�K���@�������d�{(���isXF�H_�
ڂ��ɭm��1^�O_�t�{{�{,6�B"����*Q0���=v�����;����l�Kf����[}��=��H��<Q-�ҿ������_��O�i�"˿�8.��A��� w��y�B�ɢ�XTԧ���>�;����䓨
Rg�P/�������ȵxô���e��y�FA'���Y}�2eh���$R~ko[���}�ܦ��՝��s?��F��K�������~94Ew:��������e?w�t�^-K����s�JC'�����q�\�64������&��%ז����âb~^F����>��"$t�wwJ"PB��Vʜ���Z DS}H�Q+�\ �����>2���=8 ��5��E&�C��&�3'y=��w��P��?�s�|,3tQK���<1U��?K
+��kVk��/��AG��,^&�]_�~�c��=*��N�76j����ݞ^ߢ�e���,����<�竣��o9���χ��I"���.�����L���C%ÎZ�;��%c��z��[��B\�"��U��b�=к��7~K�O��S�ǴH�� �t~|�豼����\(0κ9/~j'��x|���64�i����m������U��sټ�W]t�T&�R=�-��Cֿ���Y�@���#�![U5|��̈�T4Ӎ�ܺM�z{lH��1ry!؇�����-6��v]~�J%^�F)u7��۟��XY~�F�gaX�;˩.�Z�>�E��n��z�ݶAb���Z�w�?c����� �5g�>�x�+�K4�;\��4����WQeu6A[3K_䌷��iu��w�>U��R� ����ʓ_Q&�t,�w|R�.D�V�/~/b�b��D�:Q�? ߋ���=�K�9��;�gܲz�wH��U�ɸ�0��=�;8��U�����@�=�0Q�_٦'s%֏��&��3���Ҷvcy�q��5b��.C�V�^N_�RH2��6�v�����g�*'����?a'\���ۆv^����ЧjV���{ 耳��gq,��]�/�)��$-Gee��*���NK4d�T,b�
y\]�w�N�|��^J�l���4	F��ĸ���,^+���x;���Uɟ��r}�}�V�
�qR��"��3w��}��qЕ�ye�t`2�K2F�H;�ΰ;h5���Os�e�m쳦�t��	���D�ذ�\�s�>c�������Bz?cR�jPH�X�����A��C������s[�Y�K|(F��l����o�9}�2y�H.�p���;����cS^}�{�Aq.�d
��fÇ�(`�,���^ر`:��ŏ��J����1�� .5oz��q�����ryt_f�ږ�ڗ��ʍ�Ku	gȨ!�.�r���n�3�J�I����q5�����7W�c5lE؃���i�����.6���ዔ��icC@a��r��S�촵�9��5BJN\�}>%��w$�����y�H�b��*�J���Lp�wH��;<<���6�N���BV�c����V���-�D�͸�y6v���p�-P9�o����6��&�C@�Յ�P]�`����t��.�M��z����2y^��7�80`���&���*�ih-���c�2�0��>!���Sq<q�ْ�
;��₫Fj���>�9��W6���=b�Ǵ����SI9�J�q�����b��F@��R,+=� 1L��x	*��L�� �2�>���rZ8���� 3J&K��'�5��г:~���	r[�E0�Y7���j�R�ݻ���-�0�2��#2;�����:�s6v}��y�W)�ަ��5t�j���o���!�҉S�N�����Ӆ_tm��l������P���K���f��}��Hg�Z���zk�"����A������Ͻ�X��?��ͯ�?�_����T^|0���kh��a��N����°wڐ(��sc���G�,��y�2�p紫)����`*E���X����¥��`�w�A��F�rr�:�J/��S���݆����i����yhK�Z��0�r�kh �b�S�S�HI��-���,O�|��[6T98S�}n�n��k���b���*]�3�I�ui;|�6��������)_�-��6M�AH�o 0�Y~��'���{S�dv�S��kp�(������FAW�v�I~`�W3�L����;j��A��i:/I1����l�6	�w��f�/ȢQT aX�V���	3�x\d�y�-k� 3&W'2ߨ�|bI�;di�P�[,�����]"d�$	��h�UJ{/��y~���ꩆ�����س��;����o����vM�+�B�a�0�'��#�x�iG(�����q�ߞ��UH>��6y�]|���l7����YL<�`��=�-G#ќ���`l�f�h��D))���T��(���u36�����d�vK1,�	E�h�]����b��N��u��U�Um��:�f.e&�T���^�w,﬿ ���SW+��W:@��� hp_`�"�KF��� �0\�$����#������(#�k�V2q�J4e��mG��Z�v �vl�:���Uq�0Ͼ��.~G���@�X�ў�W �>y�&\�L\-��R=��A���4LE�3�u������g�?��`H~A�ԵM{�?UeX(v��i��b㉒�����֑�����J2/V���.��b�Lc?G��:l}��3�f �eV� $��PւF{n�/5���X�6��0����wQ��jt>4�kg���������9��.q��z�v��~,�l��l�_m�,/��^�,��a�����O�e�IfMʲY��NH�E�B��M)�{�	OZ�
��}�OBJi3�));įm�zOo���ELV�t�s`��U&��+�AJ���k������ā�^��l�c���t\��v��b�be���)�gPL!͎�>�(h�*�Lp��S��a���_ SI�dP����G���1T_UU���_յ�G��J��MA) ����(Z�nĀ�@'آ�|��'�4~#��3�����d�Kb��V� ��z�0�+�sa
�z�4�9�{pl}����[/Li1�<���.��t[)�X�@��+ǩ��JG��������g��~�ў�Jo��A�d�I8�s�[°�K\�>�ߠ���dʍ¾����m��覐��v�9��Ӷ�������{D�������(s3v������(�r�7�1O���-�zȜ�B�JjO�l�Uy
p ��RMS5S�%d2 K��I{_��F�	Z�-�HZ	����m�n ��tT��O�LqF{WS���0P�`k���G�K!�:@u� {���#в1�Ҽ�/��H,\`7ܓ�J@i�E�={�����7���LZ�rW��I���''Nmq��&�D�4;#k��"�#%Z��U�	�j�. �H�������y���
��f� ��Je�x6I8�Ɣ
���.j�}&Ќ}�t��Y�A��%���5b��ņy�l����vZe�NW`r��0�旳����8b�ú#j_7lr��`��gi˓�)%�U��OR�!���h��c�Q�Ã�s�Mޗ���;�(�[��^w��y�y�=]w
_��}X���kY��:`���vJ5�n0�i`�s���[����e��Z��{��Q�y}�K�e����hJwI0v��uA��5�Nv��N4[�=�0dYR�σL�ǖ���$���I��T�j��K����E���cYؚ��"�*�L�x����R
�i-���|�7#�QX	�:�\%
���r������L>}�� �v�R��L�]k0����M�[7�D2�I���h=�0�ST\\n��|u�(��a|���ڢF[�h�tŎ5x>�)-��I2�����}��Չ�H���7;���P���.�D]�z�u5'����K��;�SoNkt�{��}��]��N�@I��_�@'q�<��ohy��fTe����x̑�������6�O��6�W!Wu��؆������BJ���z�.=t}#J�V����9DM#���"�$�FNN���R�;$-b~�:�QT�d��������A�a4^LkC�ݣ�Y3{�M�>-I޵�&�͵d7ϛn�_�^�	���rV�����מ�ӻ�rٞu�;i���X���z-����]��i�ДH�`�?��*kH�N�n7K��n(��nh�����7���
Ur�n� E��=��-�ۚ�E�G��x�� �/^�4�����/,���3�ww�VJ��H��w�3\��#=�ewhK�X�@�lfHiP0I��cd����["�0�lͩ�>:���ȶ�T
.�C��C!їi�t\�$zR"�Fd��IZ�b~/�PTܦ���<���`��;�l�`������/��>��^����ٽn�]�n�k��gS�/|U�>�Fk�Be^�A�*�g����W\���##1���J
� ���"�zXW>��[�g�|xm�!�{.����2P�-��x��N��]��9���S��=a�L�{��+FK�"�f�J��{�������S�Wu�i-`��_wl�ϰM�5�<=!�(�QwA��:�V;h�>-5�hΐ,8�2Q��؉�[51��%�hĪ�v��o6���-7KQ�����J�
Jv��F?V�Tw�x��H�P�s��J��-.^���B��.�[K��cJ��,t�%kl�
�[�;q�뉆&�-M�8���ܥ��=�D(�d|��g�j�����y(?�����x�>��"�P_��U�gk��2(?m�D	��D
93K���+N]V�~�����j(i&�`ݢ�5�+2�����������U3�{Q޴[L����<o��� ͱ����Ϡ��!g�^ڇ�n�z��/�|��O�}�L�K�Ɋ��w��e"��܏1�z"��f���[K�6���gj������כH�����W@��H�{{��H��E�+Și��������JK@���UN��*��D��e��7FE��)�&�Z,.��{6���{�4�1�X��C�о��.v)N�:��+Z!q�Mf ��4Z��ߪ�MTX��"��R�B0g�&�u$ ���ƚܠ���p����. ]�u(�ԛZ��I L�m�K�sd$�G1cb��t�#S:ovmE��+˧�/�y@z*d���z彦��IvuWj^w�/7�.���	�U{Yz��{�*0�m��b.OQ�t��Xc����faaf�M&d��oA��t��@N.p�Rj�!�x���o����vgYc���7�5�^�}�S˭#Kγu������➀���f
�eY; ]^�S&~<^��]�ê���|�8�X/��%�TAS6�C�������Qh��W��mF� ���+�>4�R	Ƹ vh`+P0�^{*�|1�����t]��p�,��l�gM~?��<��ʳ5^����������5Eɝ)�-5���;��2L��V�"\��g�����A�G��Fʕ��=�_��]����ʟ]6��Ъd��^�V}����� Ӟ0y�T���gW��,��j�r�����cn�裞�Ν��+�t���ܛ�! �jX�ė-�����d�
���&��9��=�b���%��kx�*$��hfݴF�O{j=�����6�ڪ��F�#�^�f�ȃ�����{����?�w���7�{B'��KWD0�h_�Z���^Bq(���Dđ&�bn˽�c��I��ݓ9Y���R��۰��V۳����������zߣw|�0�fTЮ��pmeo�s�#��/�1�׼-�E�@�6�  #��y;79}��|�:���������j��A�6 z�K�x��k;�ߴ��(�M@L�b�t��B�tݥP�*p^t��[sE�K�s�i�O��1�浼����B7 �qI;����7&�q��E ��3K�������ԓ�Lbg�����C����M������4�?ѹNj�����{_�x�a)7NS?RLgUE�X=�_�w}!���j ��_�'��j�$X�ꊨ�x�^��������Z �Vfd� ˂ZWi�8�4�=�ډQ�M%��7���"\ ӿ8,�L��M�)��V���/� M�:)���@����?�� ����<�w��ZΞ�[<U��n+��G� ��$�T�[�@Q�͐��igOO�։� �0����>NǼ�b��6@;�/7F0]@�~���$*��sy[�.H@})X�ԑ�G9���.��aއc��z1�p��z}�wO�N�J���T�v����F��ܓ���;(�{N<�6yu�~s!3�P`�ڲ �I����a��7�aVk�&d�%e��(�Z��%؂%ik=B �M���ǉPD���ѯ��-��u��B0�e�S���6V��"A1�2<�h�ܭhME�}u�#*�����]�?q0��%;A�Ŝ�.o���K#|�Y��ncw��e�G�"#&WÇb	���m��z���db�İ+l�b��ShB8@�c��n��(�<&3O,�C�1�jQ���������y���h��x��ݴ�B7=ӟ�X�w���$΄��&�/1��m��ZEZY�\͍�2���
!%�1W�)P�(&���N��<�WHM)���䡥揘���j�P<$zm��G����)�>�n@�(B��3�):��q=G=G'=�^Hi�S+T�#�Q4�	)��@���2+y���M��x��$,��2�����m�?�Q�l�v!/ҵ�&�
	����k������/ ���m��SU���%UI)FNV���c�T��TP�>����=���˯_�bV�V=��Qn~��Z�7ƾ��C�%�s:#�Y�4��j��z��R��ǽ�+�'��>&0C�.�g2YP��a���|��Ty�*���k:Cq�UC{8��`]_r`E1�%�V7��\P5��h��٦u!�+����{��ٴ�{�ū!z�bLv'��ׯp.�����_�e��O���Z���J�a�˨Px�ݘ�Q���@E]�ԛ�#����N	� A~�yέYzY��HU3P54���8�T�<{��݊�]����K�&��[�:gF���J��l]x	�����wq�Zy�e^�a�8*7�̝w���阓b�J= MGp?Մq�{�J�.4���~�R�K�m�,X��pX]m� (�_4	�qM�#U����`��L�:��Yl>�~�+yY�Ǉ�������oʒ�kƶ��81��cx$Vy�/�*�������q��6��E:����Y(�k��a{E�Ї
�wZZ�aP�TB���]�ѓ���J��AGĖoj�������@�ž���I�����L/��ʉ��ԉRi�$m�:�V�؂�\���E������pPt����snHW�6#��<�к�ХN�/4�����>�������Y��s)Lum���/&�QV����/�Rl�?Z�]�F���m�fW3�l�~`�9�'��n0�v���ufV�N|�bo��~8�ˈ�#�� E���h��������2�D��q��்}z"��z�U���:0L|���Z���zc��!C��Y����]𢈥��^��w��Vv��%���c�#���%�Ξ��V��Q���|��mp��K�3�q��pH~�dP;�a��!�s�ռ�m�����y��Y���W0�R��0���f!�9Yz$�,�\�u9 ��mL伸8�m�Ծ��|z2�m�y#1ϐ�����4��Z���ʪǘ�s)ot�k�����|���+ D�����ZxV+I�6��ٺ���C�4$��)�ۘ��e}�"]!5x*�����(��������8C+����3#�
Z<��l�宫���/�����pғp���s-@��U���H�U�X��1Ht�;y<�{�늗!Y$�Я{ʞ�u=��(���I���Jtq8�j����H�ۺYG)3&W��&�h�=����N���8�� �Hw12�{t;�L㯚����[�:���m�t��'L���t�.�?���Ս@ŖJfS�6r!��y}L���=0�Z�H� �M`�7��	�K ������ŌPɰ/���p d��~��W=���2P]ě��I�wV)��^V�� nl��U��D�h�������j�k�����;-a�ۣuB�ć�	�l��XAK�)�1����G��F�֔���3;�Ga]\.���I����|���K�M|���#YK�x��P�g��3KsT�a�<-wl��G�����C�E�ʥ���;�Ye	�S�Yam*���ϫ �Io�A�>48�V_}��E��<�2%����s�=l^��-LC�\}�ؒ���L"g��G�Qw�)�}�́m3��4P7���ȁ�P_F�M���;��͟��gH�|:���b�/����`�P�B�����<���XI�ʼ��#���BN�y�"[�W!c���_�3�/)o�����-2���d����3�Nh��J"�lVb�4Qw�YZ�)P��wQN��j�5K)*���B�"n�^�XX�o\4l���n{�g�$�
�ؤC�kb�xh^9����t��l���8��c���Lx�Y���=	w �=�ٮ��LS]L�g�De.��*����GWRm�[�zst���JM�%[�r@��T��y�UB�~����{yS����p������$j{������i�kg]�x�U[�K�_��:������aV"$�m=8����L�?��$N���>��)~V��<o�G'���#,������"
�;�LIJ|dB��=�� 2�.�K���=�G���Z,Ij�)dC�ae����h�
�v�"���<��9�;G�mVa�]%��}�\��n��$��>?�l�cۏ,<����������O��<�K|�`W���>�m�3�G�_Ie'����G�W��^��V�Ψ����I]l^��tM�Ugs.>�}ZC!� ś����/IeU�y��1��>���>U����%�����ْ���|���Ė˨m!��c�[���J^�����	��b�V�u~����w߷��F�A���5�H�Ac�֕1����:��_{w��B	Fp)G�q��-��d��o��!�ٍӃ�(o훜����/(�1��Q$ػ"�t0����oXlͭ���*�_�.���_5�Y��h���P��y�]���O?�d����#~���) ����O��[�Y�wq@���A4<����ώ27�@��d��|p"��#)c�q5�������9|�-��8�C�z�mC��%k��j�|��#FJ/��i�����.�e�d�%}�I�'p�������8 c�NI��=mܪ P S��P���h�Ër��8�o�a��gTk#&�p�9�%�����0�4����\�$<��'x��]8.�f�j�&�I���7������P�
q��ވ�f��  �L��5��u�M�ݢ.��6a���hJ�X(�x��(&�F��Q�>Y�)��C�zSf�]�����z��C�� Yh��t0�N�2�S>Q�o�2Ɩ3�o�V�`R��ŝ���k�>M��=���WpM���F�0u�n|�$4��-v��G0O�XX�+���67cZ�#bp�:hE%��jOT���<"�[]�G+!��p��x���b��=�AB������^N��LdK��L����Ѻ��ܙ��3�����d5�䅛5T���5�u}nFc�<0�j)�����g��F�ʻj�9�nt
(�/k�?P	��f!���/p{Z��@�l��4�'N�qM,IƧڃ���VV����ȶ�~�\0�����v����<|�̄�Aut�L`&�Y�è�JS�}q����Z!�=�.��k��o��a�v���3�w�o%�(-"�vM�B�����O�y� �B˭s�io��i�e��'�q�W�M\�+�.�V�%�.��LYv;nߜ)#{ʿ"%r_�+Idj�M=X����=M��������`j��}5]�=/�����8h�I�h&���E��oX<<��%�Oα�ʽչ� n�w�̈́0P�nS@�c(�`K�J(���_�N>��!N��Y�d]��\Rɀ���Tw�R%�Xq��7�e�P��@D��y�A�����L5O[/p卵� 7U�P.P�Nݒ��t�<U�:)A��h-Ο��m^L|���҆�
%�͓-��$F���no|@.hg��@�:G��4���>�٧ǽ��i������x�T��Y;���q���v��l���t�F��v��Xa���B�b���Cś�F<��Dq8�$`�,AC���"������2\�}��v[_N��z��0{^��!L���ؒ76	�!��m���
�R��a<ũ��}�O�US�fB&�T�>=:n��4ĺl�#@���v�������=<�>_3	:C��t�&������(�%t�S%S1��W������v��RQ8�Z���l�_*�Z#��s��B��-��f ��/�6���㮜w�_.�����E���4[5��*Ԝ�	�{�܏2�3Q�}���M>W�{^I�����+z�q������J	��P����f�?�����^ď��>?�we{I�Q����Q���I���� 	jG�;�,�6z?cx^F�e��J�qK9��4�֫�^s���:���:��Om.4����ɠ���-QI=�nk�-�����/*�2*�m��Ƃw�� �%����!����=xpwww��yo�y�w��#�F��U�j^sUu/Z׎F�
��h��Y�v�'Z/����[����Q��7.��(�o�F��?n��������c�a�*�������mce�Y��6{D��/7�gEI#�Eďi2������^.�Q�bС��G}�D��;~��P�zCyoɹ^�PW" ��+��{d�,k��>��m��!s�˦6Y����Vƥ㥌ǩlXo�%��3���5��}��G�U��st�G�%���8ޜ]����������(���6���j�x��A�j�t��0������A�S�V����&��N8J���RԳ��+\?�W��Y Ồ�%^ K���V��r�m��+_bde���_�\�2��i��by!����Բ�4�����:�����P���@�6���sBEfa���Đ��c���@�ʳ��Q��欪#c�)/��f:��UJ��&%u]������-3�O�J[�Gzz��(�`��h���F	��%� p�G�,�ws��>� ~)���w��hQ�
�΍buX2�7����e�5��E�7�N���N_�?�͚p2�3wwPtn��C�6�r����]Ę���,N��Z\].���շ�	��R�]�
�\�N�kȧz�c����S��nr���|ə�i/VT(&��X�r�o�F��|<nz�afV�s��#�j`X_~�I{N��tXJ~�'�i�כU�G?"(St|??�:n�'��+�w�u��1��}�4�G�vp�~X��O�Sc`a��w�Z��*�}���a+�u��	�J�s/*֢����}��m�_	�ܫ���b%�(�׾��{��)t���1�\�g�>�m�W�n�������8-�����L�ۂ-���ǹ�.���W�;�wv1�kj߬��Z�:/`-�>C�Dmp��͒�����t<��8J�OK����=]]�:t�.��D~�a�r1��������x�'~݂ea-�k� v��)�����{%5�hM��)�P�EdP�ُ1#|�ŉ�߂E�(�z�7�����׭����r�-�3Q�i����L<ޮM���ա�p�����ҡ��E�yL�t2p!}u`�)�Zb�V'�{���Sв�����i�aFd��ѩ�A�ɭ\ճ��7��}�t�Z�Bv���P&�#���2��3Q�,�|̢m6��b�����j��K���s׍b{f����-�	����}+\M�11�q0�{j��;ײ�Q�~��=�O�vS�IQ�I�~Y��y�X�p���S�8���^�A�C�+�D�k���Ā���%bx����n���k;�6�=!��[?�o�;�ƅ{O� We��g��I����>nf����RR�C˘�֛\��tFpLb~8�����5���P��d�)B
��Mҿ��{_,�h�>���,E��\���IŴo����ٓ)J�$�"�~?���yaHV�L�����������*V'W\�و��72�,�se�39��0gpjq�Ƶ�ɨ��.&�\�L#��7�Y�r��{|n�Iptţ�O���XP�
���5��[+������qm�o/9[jGG�hM5��\�-�VO�%��ن4�'Τ�ȁ��ô	1_#N����,D_r����N����$���.ގ��n�}|戀��,ao�C}-��e0�����SozCr�Y-yi�� `��ٽ����#�S�m�u�Z�t}ƨ��)z�c�	&YS*I���'������f��B�~��6�+�m�p�����hjo�_ϊ b����љh�Q��v��n 4wF%�pO��5L&��J���>�x�r -eq�#ɟѲsj�ʮr����ȸ��5�� ;�6O	�6!0a~���k?��Ю�����l�ʼ_��+�����l���g�-"C���;o�QZ}�fcx'?���"�k{��h�t�6fB�}D�k0�#��6�K��4�{�kǪם��E�v�˒3'�}i�P�p�u�X�|�o��Ţ;�(�3x�3_�I�#.z�$���)��o>Y���}X����1�ƘG�r���<��v������JגӬ�5�C˵��Q�3��[��v�x�?7ihV�̟�*�#g��g	w��B�p3?hC�`ևA��U0�1s��ZhO艊_ �y	8��VU���ն�VM��ƑǊ�VuГ�OG�7g\8����u⢜��i^ʖ�%����7c�3�g�A�ye豪�%�o�.��c�} ��7*xeq
U6�(O	�s:��|	8�g&�zS�J=�N��o�L�����66����҂���~�<�n�;:O��<���!�8�����.�������P�L�	��S��`oZ	v.}[�ׯW)yI6��~����Ӧ#�~du�˝���hUl�� �^�������gط���4��=ǵ����3��?�����N8~�5��ũ��n�[�=��T o�	&���Ri/OH��.��v���N_�~%i��X�
p{$ܙ��]��ezn b"ӂ6�J�+w�H����f�`��^��4��i��j��`�/�*�q��H�ԙ>�`T�9/5��m��l`����yY��Si��Q緝�4b��X�#�7���4^�z.��<k��q쿠�M���i��d�|��<�8�'@ԵJ�,��Ym�K���.��c�˸\����)��fE�K�ܺ�He�9��]�䦫(�i֟�,� /�/�ۉ�.��Zl�M�>�Z�w���7G�i�irt	�o�?͸a����o�oOT��o�ܟ��`�KKK�L�-e��*;����^_����M�QU�8�^<��g�}��oW�oײ.ڬ�x�o��n���\����Ѷ=�(��T���[GQ	/�$��heR�#�ɪ./L�SN����8���z�yM����� $�rB�����Y�PI��	F��*��@�Z5�c��Wk3��'��D����0�g�8ӊ���,n<^���=D~.����6�mE}���'�g��zے�sg���m���x�A�ڑٝ��e5mα�sa�����.�T��5��j��X.��
~Qq���2��=�k��,���S"3��auq??~\Wϑ�4'���[\�ź}����3I����@e����6#�x������b@�]Tu	��V���R��mC����vp>��ｾ�H�n�~v���}l~a����>�kHf���k�pPϹ.Ki���J�.�hP�^r�M�2��	Idzr��x���|gw�=6�G8.b,��$?��5�g�vAxF�H�����^|��l�����*O҅����G��-�,�����x���uz/pW��\m��@/W^�E§��ٵ8��Ǻ�`��%$26��z�'���8O%RF!��;���eZ�*���J�8<��q�2_鷌�����?*+R�%�Y��Y�RL��$�ƅi�LW�g�q�JBp�4�n���s*?4��ܑכ�Tێ�9cE��4�Y5>���N��Q2!�3A/��!�)À���d�o����&~�~�"��7Y�`�M�Ȼ�n1;od�V�+�v9�דTf�~9_	?:*�=fK�Ny@J�В�z��m�qs_���	�X�L�˱^)w���iw9=%P�2ee�_�ݯv�|�s�"9=�)�9�ë-�*n�[s�b�ymdG-�!H�/?�1`72�0��a���B�bY�ӻ2��^���F͵�|�@E�s��ڳ~�1D�jvh���oկ̮.��`��ڒ�ҡ�_�'r�v ��w�Ca�1+��{n��B�u��?_����\>m�w��$0n��7�.�� <ū7��8��j�ǭ�u�z�����f��@7괬�>��}�Xn`����_v�]�����F�jn�-\Iύq���̌JZ�T�:��I_�B�c�8֗K��H˿��}v�V��� ��񊽏��Ngx�mB�O{P�y�a���,P2�)���Yj~���i��iN٣�i�������/V�Q��~�uL�ǣ1�|o�O�����vשN��.r���0��zE�۷�B\ԁ~F�F����uA;jp�_��;61�cc[���2���-�K�.m���%� ���#�W�KN�����I[Đ�3�ݫT�Nя����d�d˥<*:���h��s�+�7D��G�]̸�.?�����O�D��D9��	-��2�Q�b9���}d��dk�&Ն�%B��5,P�������'�*'7fi2�GU,��}��'n�MBrXG��m��慄4�Ѣ�`�Lٌ����H�oщ�SA�����T -��U4!����'`޶o���y��U,#�.���a:P�o뿕B��k��H��7�.�r�ы㷽��f#>o����읁.'�~���Ŗi��v��/�o~k��PP�%u�WH��}�xQT�F,�3c��mՠP��:N��v@���N@���9��g/�Y�F!��m�����r����3#	x �4}�:b���jw%���0�掅�׉�p�{��;g~V��m^���@]˶��;�Z��Y?��h-�["�������jȞ����"Or��N��kW嗞������ۆ-�KzF%V*�6}�#�;�1��Y�α0K�+���겔J����-�<WR�8��f�^��L�7�����
)e${�"�5>�	mF�j��5@��Êb�H��~W����f�����B:�bu�^��-��/�e��oa&| �jJ>��U���Jd���y৙o`hZVCy1�����]��̈O�PžIZ�T ����v��~���C��EEح0��"djuX�%�j&�ըBÑ�&S��d��iY��,'@w,�������W�����>nm�"���2�����Z�r�����3�B��~��d웏a�)��o�Y��h�z� Q2����nc��~$X�"��!Ҥ��.l��ۻ:�����Cmn��ٍ�޹�R|$�/�͚��?s���{P{ �}�P\IV������Έ�f�p�3u�p�p �+т~�Q�5 �F_�i�f2Ir0���{�w� ��|�ҧ�(	 �p~%���b�����7�;j��L禷2����7�v�,���X��˚xe��r�QA����?~�;.~�m�����w��ә����j�7�?;y.����j+�`\��fh���i�Z�?-�m/��mǽ[U��jk�W�ƿif�x\{<���3n]/`D��V{n���=Ľm+�����;��={��s�'�gc7xI�t���-���kG���Q�����`	Cj��>����m��;�BG;m��8@b�F{rQ��l�oWr����D�@���>`�5��;�<��vJ?��}�W���dZUz�Z�YK��^_n����v�ly����>����h*o��Sa�!4%���-ˁ��2/��R�yQ���D~ys2����������ׅ�(՟���UK>���-�����ٿ�Q��Y�mr�UV36�zι�)S�]k�g�O�KZ�0�{��������M�?��}Wy���W�/�dp���&M���aVҤ���N��UG�	��[���u��,��<�+�S�Y��7s�jJpq=I�U�j�<�^��VD��W}ĭ�`G�Ƶ�#i}��YoE�L��%~[��?���|<�c̷�C��&�v5�����~h7�Yv�B�+��Ův$�+ӫ5`�&�{�m�������>�w��A0����iQ-J��ϧW/C�{O�����z��=����˦6dn9s,/s4�4��!1:�-s�~�)��)�5{�5N�giw%���������Xn�>(��<�����#�r����8�H�<`�F��,�w�S�:ÍŷZҶ�8/���5�bP*��<��ݭ�	i�P���N�R��jL	�Z�,(�� *�+y����0FGI��B�i|��Y�*�������^,���P��@����ތ�<T����Um��t",���\꫐�xn��)^�O0| y��\{}��D�K��"�A��kk��q��y9iXX�5������T/L�������:�5��|�vg��V�{�\AN$'6��jB�ኬ]m �6s����R
�{v����-݁��*���պ�ӄ,���XMU�l��(.Wr�G��|��9=�ܡr�Q�qְ9��v��M��q��r�P��G����e+W�>~*N�ȹ�("Ɇ9�c�ɼ����w��L��Ⱦ�;�b?�X=�>LÉ��j�<��> �~b�U�뇼.HW{lQD�y+����pA@��T�g��6��F�T�O�/<���R��<��p�"�8�$c����J(t�/����S�,�?_�h���R�M$GM|��C/eϼc�!�DEF.����B�+E����K�v��,��h��W/V�$�}ar��WC\�,u4W>��+y1����,Fыa<��d5D>9	�	�!Rh��"ܣٓ?���դT�]�Z�����;mu��ĩ��aa���O���/�n9c�i��"�_��54�
r���b�<�)�Ӹ��3V�g��-��E���"mX=zQ��a�~���ʏ�M�vp��k�b��nf'�j+�Ȧ��R�.[!H����Gom�_c�;k|���8��#��X�1W\�p�t-��cPq��Q�Z��ԏ���I>����Kn<+:���P���-�@]�2��I)�ǋ��`y�!H����*��[�A,�$5�j�sW�H5�V$SS��x{k��%w��aD�WҴB����/9ٓ��Ѕ��� vg�6�J��h���`��oC� ����^֥�TM��KS��n$YS@���26b�0'8uL}}z��7_�k��?��A�K��O�EhT{�0�/D/4��B�""�G��y'�9�?:y_��jֱ�ᝍ[�����."�e�x���4^p0�͕]}�v���	,�!�`O��Ň���JL�����Yi�F����=۵@��&��j%kǥU�4\�ӽ��n��bK�溑h���U���$���<Y��c��J�e�yl�B�&}���������!/�O�3$P�,K3�9�Ғ���Wh	gmW���I�,Ku����	����-�I�R�ΩԷ��u�.��}�*�ϻ�G��XE�,����V6�6��
J&�uM��Ө��>d�|VY	��&��Q�� �����ɼ��lt��#D-ӳ{6���7��W�v���հ9��L�@J�T�A��#�j'qL=R��AE[︅��b�a��^��M�5�U,J�,t��X�R�.A���s���w���B�(.Y��T��u�=����冘0�~�Mߣf2$h����Nx�2!�Z�wm՛_G��U�1�V�s�ȶ*9��g��(��-�D��&A�t�����Y+8|4����fݓ�Q���b���T��ōh��ȏ�*�?�X��%YQD�$�5��'�s��6|09�
X����ۏ�4�O⥙o]u=�ߦd�ka`�7X���r�/�БYߧuܸ�i�D���O	�'V�S-�_���5vU�HU��.�Y<�k�['�����:'��gY�9�$�ޛ���h�Ξn&�n���e��(�������㎜F:b4�N��_��bV���8-+8�PÙ��Qf��2�'�E�W,x�$��>J�~X�aے�nQR4Õ��,�:�;�����9����R?�K5S5��s�����á��쏶4� S��!��}��>vx�5iC�&۶D�����HPȣ���/&UݵL=�
��ǿ�M:�/������XN6F�FTF�n1��|���*q����(�
1Βy^�
�� �U��z�kk��m�=��~�T5Vf����xKH m�[�������-��#@�/��)�t��{��x�4Y����z��Q#�̈́��\Z��s���|��r`�㵧e�C����A�a*����i���t�q]�F�eʇ�b�����0�@�����ϊ�������Y��O�A.g� ���5d�vGv������Q��k�^`D�K�������1�8��%���@�X�]�#��Dpg�"Þ��uC��<}�ґ%��x'�&P��m�Q�u�������,���8+���O�
Y������8�����2��mP9l�lm�Հm����Y.\�Z$7�Y��� Y�R�f��$�W���+���_	 �E����ƻ�=�kr����>�6M����j�i�����ZZ�*-?ga=gȧ��~�����[Pt��i|AF�}F���C�b|+ݑUIm<᱊] ���@�!�xZ'��~w��I~V�8�7����n4oLޔ<�B�%�LŒ�Z��A�{�4��k�l��IГY
���>ω��m�fX�vA�e_��v#}���i��\h�^�K��N�WX�	C@@B��W�c�H��؃/i�-��9�3/��lY8�e�@aî �'+ȶj��8"�{���O�������!��W`�xE�\�aO(����������0�c�H���@t��d
������4�P�onY�:��MSJ=( ��)�]ٯ|��5)�7�E�
��r��C��js���Hj"�NI_՞z��Pӏ||��k��o���̔ϯXDh]NL��#53�)�X_��៟[}�
��*�7�z�by�¯�2�
}6A���|�=�3���8[k\*�:�G[%��(����s�n8�'�c�|*�RR`��E�{F$�1���j%u+(A�	IT�,�����B��)󈗕��O�v�H`�h8���&�W������?#����l��%� B�"���>�8���aHM�&�C�R�6��-j#
<�'V�/_	�B';����y�W� #�r��� �Qf��TNd ����5'�&���S�6Pf��Q��M��`�L�ǣ���1Q���b��]�Z\���-����wf(�*i�����p2�s��y.4s�#c�aKA��� Hї��!�;I�x��e���u�ە���6D���O�O��9�VwrXܪs�R��A2Ԣ�2U�tȸ̚�%"�%�
��VM�*#B\�W�iˮ��*W��	TS����q�a�y-�Ez�(�~��00�],��D}F8RiXs1�&�]?d`2�T���ȏ�~�&��&�[݁y_ ��+Yh�a��VtX�:k.��<�y�_+���� �ԙG��~N%��� I4�ݜ���J�W��-,}"e�<�����m��,����E�iE�J� ��YVÚ�Vhou�ƓD|K�N�������z|��j*�������Eʘ�Z˱��o�;@���+ *?�X��H����􃖦14���d�׊\����SG2F��MI�lu�θc}��&�����\u��HE�s��;�m{�`#'�����)�1��;уנ��J���_�r���mV3��WJ��
�N�����ٸ��ݚz�?Y����	���Y�W&V��Þu����#��q0Y��t�6٥�m��H�X��1�����i�X�H��y�!>�FSnM�{dߊ��.��F�cv�;\8��<�"4>Z�4��l8=e�@�x��̛�-��_�'��;���F'\>�zg���7�E��{Xx塙 Yjw~����?��|�I��C0�/˕r����R�����Y�4J�OKB��dǵO�(E& ��h帔��Я�͞��Ff��9��2��
%���.��#�b��e�ԉe�^�c�QK�<��g��!��� wl��z�o�:/�����!F�N��]���/�RX���<���������k�,��/���#~;��)��&Ǵn��K�?�gE�l�X������
O$�1�ɔ3���U�[̳������M�r�*���I�a�:���Nv?��rul�7��������'�0�U��G���|�,�-z��[�x�B�����8p������d�ù\����0:�U�/f�Yc���i��qB &�eq��`���B�KC�ND8��i݆�E�ˈL����W�	QK�g�B�}ڻ�$�Y4U*$���w�Z!��מ��[�IX�0G2���U^+�JZ��[��Z��"O/�w0\���5FY-����y����� FVlS�h�����I�2a+v�J�T>[�Y T'�f�������j�1�1�k�D�'<r��Hx�8T�'"�i�H1�;����9���Q�D�.#�!/�O"��D.f�ǟu���a>��8ˆ��`�]�.����|nCB<�����&��_�lվ��gl}m�Ӡ�R��M����-�x _]���G�2vb��nRVJl8e� Y���Z��F�Q��PH��#po�?��^
���Q|S�ϻ��{Zu��њ�{�/(E�%l@"��ρ���uq�>(�or\b{4��lpw�Iۜq�Du��fA�_W���S��U (,��|)�=H�!-��l���O)���|�p1�"�\�~�ՠ��5#�pԇ&�[+��_+���R�z���y���^�y������,q���;OO���t�3A�>s#�ɒ��(�����o	��%�-O��?�2`aX�!%�|�65:H�� +���u�TYL�����џ}�t`��7	q�|(�uD��Eƛg�F��u*���;�����IRy%�����#3���� �&���N��/'Wh��6h>wv�q����dzJ�-g;1f��#+�#�5����¹��@!Jʼ�x@��A�ó���
�}i��`F�������N;<L���y�������wW�$}&��}�<�,���_�x���7⚞�E�Sm7�g��I�� ���r�������=b�e�@C`�r��zP�x��������{}EDӓ���Ә�6L���*�k}�&U3�N+���2�p�n���\&�	���t-՛W��h��Ts2�����K���b�����S�$x0kR�&�QU�LG����qh����J�Cu5S�7̘?CS�k� |(#%%$�ʋ��]5��{��$|B�&�,���o�1�iφ4z���P��}K�J��R26�&T�o��[y���pm7_��������ۘ�I�f
H_C��cE�ٳ�NK��F� C�B�q	B�TC�Ǡ�;h�&��4Xa`N����3_�9b�s	�V ��z���r(w�8���%�A����㘄�<h���Y';#P���=�@��\����r��ݡe�L,]������:�F��]G�n�O��nr�˻�/m�>�v�d@��+�5�ԉ��MC�'�S��5�92�D-b�=������V��p�R*�#�rr�q���?a���t"ȏ9K�):�k������&>F�{�?�+^2H��SR,����a�=(���6{�,7��چH��F,���g	�O"1���u��]cs����}�n�#��F��(��y,�����'�����6���꽎s�_N��釻=�Ο�{{� h�)		i`Sn9�"5�'�ı,��&�K�Y"oU"vbM��s)�:0n�	�%~9Xio�K�L�����H��>7gg�����T[�AM�:�J5T��eP�<����<M"[�K��i:Y�R����UVo�W���g���XU�5�P�����N�ny"���+>i�0��)�G�NS��c����Zh��8�<e bhp:������#S�Y�*����-�+���F�ۊ������$U�$9"CI9�����C�3����:����2�Y��c��e2`�����s�xz�Y��Cy��Q'#�_t��h|�5�G������]��x����f�x/j�n�ˋ��.jXem����=���.I,R�7��&��4�1>t�,O\�l��!�)a����@�&H"�t+�_v��|%Sʕr��A٤ޚԕJ1�`���I:�����P�by���PK@�i�]nF,�[_P`��ǐ9�磵`M�R3>k�K���0V�:�o]��GT �5x�Ș��~�HNJM��v5��w{�����[�,d*s	1�ч��V$cϵ	����y���xu6kz۾CM�F
��J���̺͆�e!`�MnL^P��ƇJ�������40Clh/\�������SD�f�#ƹ3�b�����Jf>||ev:R2e������ ��~�NXR�A ��l]������:�������-���r�%i����}#l4GT����6(�l��BQ#'΢��|��KTMi
wI;xm�^�@~��.d{���^#��5o��n�c���_Y�����r���>�����w��z@NE������{?�e��II��!��.`cs|
a�RJn��1�w�Y�>�Ͳ=��\\���@�X0�j����+d,0%H]��R1�=c���E��yfy���I�^46��$	+4(�P�ۘ�m&���ɗ`k ��#d�)ҭkE�DKy&���;϶t����\��[9m�C��*L���e������'�=5��N�o^>���1�σZ���n��d�\b��G�]�w�,h��l5u��&Nu�ἳ��Bo7����JPN�������M�f��>�'c�˧S� �{ �3T#Ja�ַ��\���bJ%�t�)uQ��M�o5����n���7�j*�kp�l��%,�u�\9��8.�tBf\��O��N0g���Vr� 9�?�ý~w�(Z8C�����T2�~�7�IP����eN�GXDr�Ͼa}��-4<akr��%�T�z��ҍi�}3����{����+##��ʓ�g�3R�&&���#��g;��e���l� �Q?RF�+��w�9a��
N�?y��&i2p�{8�ah?��	vwx�/���p��/b��#O��X�y�-!"�y���&9��H�>�f����k�v[�,(�"�����������7EF��cE���������!��Y�V2���U͈p�.�u�+����"����9�$,׵��)�%�~�q��c5`i�#���/')*L*���29tR�*�������7}LJz����Z�G�&,�ݒ�K�x��7H��H<=�5���1��S x<�""���P��Xo:<����,���~�B�U=�rm�=�'��C��x��au"�Յ�DuE'] &�����AhQ?ݟvz'Ɏ�5�.��x�at<<��N2�e��5$���H�=V(j��rE������7������O^&� H�IK5lu��O*���v>��j�!r�n��uH/%G����E�dOҲ��]��:G'}��o������"[���[�%(,�����?���V�#�s)�� zT7:�u1�5��� >�K	�Q��l����-�i���#ɥ��jc������	����P%��!�F�Y���TRh݅�+�/3��Oغ�jiDS8[�i���_��s�7Wfn���0�N�W6D�M· �g�މm�Tl~� R77�� ����k�hM�\H �,�T��0�n;H`�^=\���}�#}¹� _�ѱ������uh��GZI�؉�o��X| ���#�󧤼����g{+Z��q�����`���C\�H��<����D�}�%�'�~�V�����n/�dvO�Q�Y	����M���a��zڋO�����-�b�������M����,Eǔ���Ž�/���`�)�� �4��|�cc�]��?-�F���WG&�36)��ng�*;��4���\&S����+���gp�rCMK�ÝE���+�v�;a����N����R�,�_�N��q����,�ӆ@�(f�uu�F=b��Yko������L�B�B�co��oʪ:c�
��N�UJ��u̗pk��hr��>S4Դ�΋��!U��=WG�����Y��1$�'Kp�y2�g`�>�U���/5��S�~��fڑ�͉Mp�
>�T�<;}�ҏ�X�����(���w��g�L��]����H�vr-�MI�8�ǹ�A�N�g���� ^+�N>�."��Dr�}ъ:��|�Y�*�?���Q�V
��Gz�@�;�\<�!�$�`�V�a��(���.V�x)��&tK�DA�� ���5�cͳ:k������''�v����3����X��4�u����=!>>܀Ѷπ�hZ/e?.�Oa�4��M&c�4�XʟD�>u��<*�i�}����:= t06�7ҫͨ&�b�0�8��D�f]kD��Xl�(``���
���'�4x�aS9��</^(j����� A/' �?�@���@��VK�ʓ��v��{���ؼ{�'����Ij{�����Ø�+.���x���#夹�D,������>z�O�k���@@�I�Q��-�_b�JA�/�Ϡ�`��PdEJ�e�(��3I&��]Ŏ����T{<����G~��5_{�@'ĢÃ���z�	p��M��SpP�Txˋ�Wk��^�3�����г���Pu��N�mU�z����d嘲m�ۂШ�|.GE�QVh�{���О#	B��������7x�Ǯ���@��~�䉂�|�F���}Q�W������MPd|���E��0����Ĝ���E'߸L�~B�S�@z�f�ס�3���?d�� h���q��[d�@�E����v�Tm��=Y�ǋ�ùz()�����������Z�K5�#y�c������UP�`��=����-r;�&$I�f�@s����Lt*�c�!����/�R�bZ���"�R�Y�����i���E�m�����2" 9W\ ��y?�+�9M!�s�]ΗG�J�.#y�NmNK�~�m{��e����kp�n���QP)�{SuO�_�����[3}�Kp";�B���#.�t�N�a��|��ِ�6��2��NO�d{2upە=�͕��a% �&�;�en`��ԗ�xn�=5�ˊˬ���?�J��u�,ƪ>B䷰�=L'��Q>�=D��$�ƄHP�>[
���Hw'*h�#�G~`�G�"��/�yJ�/u�/$gx�Xrl��/g‬q;�T疂��m���A���kzv�DJ!$.:�������7\B��;�7��ծ_E�����a�Ӂ7�'�0U��)?-�e_���ń�[�{G��2knWcf��=X:�%��W�K��jE��!j�^[Z�O�^��cz���1-�����M�1�������QD�S���':O�4 ]�.Y��c 4�w}E�>�f��=zO.�q{�h9�l�s�$]�ۭ^����ϧ�c�>��.v�⧿J���xO����)Z�u5p�+�ohW�nw*��.��n-X��Y�]D��n���Y�̰���7����H��=��,�o2$^"�aN�!S���R���M;:�1E�Ym�R�$*����6Ɍ�b�1���6VFG5���s���Q����R�o�]S��F�ͩ)��ʿ��w+6C�a��I7��4�`	[�RQ�x⸿3�盹z~1�ڣÏ�X�0|�H֢}o��O�i�ժ(��u��F;P�j"#�2�=@.�?��ć�ū�ˮMrJ����&�����r�����#5�/��j��G*������s�ץ!��#A�u`�t	޶�bAfp���Z"������r�N����XNI[�_B��#��λ'	�E��
Uu�y��Ȯ�su"!�n>�vQ����a����K�r�qwx^3�)�#�XBJj����7�;�~�M楠�K�S\9<%�΍����k,����O߯<���˕0�P8^ � �{�2IĹ =4�<�LSlk����o��.=�9��mr����i�18y�>���c�A2Ի���)j����|z�A���%U���:�N/-�3��B��k-�c���� �7�1�a�A��%2]@{��\�$����W@���`��N_F�R��\�]�ks����)fCqݶ���(J��iD��;dAjAu�3)� �'��a͞�c�D&΀f�7;�-4�{��;�E7����=z武�*M�
�F���K\���]�Qk� �?�����0�|�U\�$�&�8��Fr\��mwNW��++^�OW��W��#��/� ��T7ցB�õk4�3~���<U{g����	;�9��s���T�~]���aj`�H��:ďZR�^��ߵ<#��x���\s�l�1���������"�xT,
B��Zv����ɦ���H�^��ʻ�\Lv&Q<+���|�:���&�Ֆ� \�l<R�[w2N���JK��U˵
e��y���:w�;�7I�h���2>��Uh�bty(}�N�[� ��M��
,Q�$��v��X�KWh1��0�^o�"RV��/c���Kۥ��/f�H���-��.i�+~E�D��×�̯2�xž3%K�٩��*U�k^�|�ɁĊ`�]nE{<�K��r�JHPL��Ί��h�X.Ә�im��g]��U�����j��� me��4yO=��%[X'm2�ًO[R�E��~&;Q�O��_?��_mq���R��'ǲ��Y;>F9���^x"=��yPu`^�R��[D�����H(��x��-�.�-��+𿲱O�?\��=��T�G �m�)�4���?w*�t��̓ޫ���!�D�j|}�20���&�c�qͪ1UȠ�`ǾVkz�l��%m�R��S��BfPY���=�#���v��^�.���-�lT��AK�S#f�$��s�%�;�N�01�:c�ێ��r��+Q�=��%���m�&�nw�奄����Ĩ�� 9����囟{�j�]%��Op���[�Kǉ��H��it7������%�4!�V��vB×�+�oߏ�\4=1�t׋���B����ү{�t�����A^�_�}+�x�R$eś��"�p6��g�hИm,�k&��uҷ\�ty��5�׊\�[�oÜhbW��b��|r�m}eT\��.�	�@p<�K�w���2!A�wH������0��m������ޜo��?Xt����z꩞*�R�VQ�E���/�&3���G�Ƃs�_�X�}g̔�=�Q�4�V��aB���9A�c%ٟ��a����-� _(a�.�J(|�Y�H�i��c7���Q��%��C6M�3�ww<�z�n���� f�]��Z1�+|�n�`:�8I�Uwe�'�/��NL3sѮ6�fu;�~���M�h��7%�1�E�B�6�b����Q��"ͫ��u,@-~�Q�'
(
^�/ȅ ��9���J�B����W�t�`qIg�r�S�&�(oy\�cP7��G-D�W�Er��FM��wqQ:�t��9�Jz�>$�?�����$�ǬEX��ܝ���3=�ҁVg� ������h�!����Vڿ3h��y5�#]鸵��VW�<����E7[���j�8��{�����8+z�����t^�P��Ng�� ��@~e'*n3�w��zlFir��+���d��PòL>0(��m�����qp�k��E��Yb2BQ�ז&�M�X.�"F6E}L�I5u�%������t�*Z�<����-�+&f�lk�F���Or��k9õ���b�}=�)�W0� ,�P�*3(�4��W��U���~k��_�%��D�J��J�c��RR��`��Ϋ�5g.�}l~�}{+��y)}�����gj���l���Ǆ?+bO��	�"�S��8�b��پ[ �ex^�hQZ�S�e�c�,XkBU���'�p�]����~>wD��,��T����E��6^���JD��"�pY�d|2�J�Le-����yO�M���r�f�^g�nS3
LLĢ��W�z��1<dv� t�)k�`0�	jq��wsm��]T��T �?�9P{?�uZ}5��\�z�ʇ���|\_6�D����`����xǯ�ҝ��U��:,�h+��G�E!� ��T�?J~�{�0�,�(Oڌ�U �c���O��T��<|�;@�!��ɦ1�;���z�ܰHe<:8��c����������!�֚r�ߕ�Ո�� �d�O�l|赼ڗH(N�n}��}�o�����7ed��ud��Ќ�^�%a���j�(,WU�����=����**��CYw�$)���~/�&*iy�o�x�r�̛��-1a�7ۏ��=�qAМ�w�C�IG��QH���`t�q컎�L�#]P�^����v�����R%`����w���/.�d�IlB]c�^�!�Lc�R���YW�,DA�(�d�����N�6Ye�<_�;��f?uPN~F������٭yE��2�6_���bZ������m%���H~ ��b��|nC�ZW�܃�|�o������7w���1��@f��=�m�Ê�IbH|�~�9�$<c���;kQv���͖��i�2�S������	�m ���|ma����yN��o\�~�<��q"ա���uf���O�T�5Q��A�¯�GQ�����z��s�g���;��ۋn��Jq:/��qe�ȽYV�N�"���0h�n��m!��<�^؇�X
5pl���[,ϳ^W�Lێp2�nY8a�A�`��'���~�~<O�&xd��t �����_�.::��~�&Ùi�U����s�������|+��|�����NYE(�q���-3�X-^	��=�U��
O�UWA��'A��S&��%�������s��0�1�ҫp��Hg���O����KmukYܮ�$[27_�ƒ��!D��;᳍�/@�_�H�c�o�xfj�Ź�H��v�(�����;l�\��<�)��ƍj��� �����Rogc��:��&2������V��rd���8���7XhE��������ʖ�W�#�{�@�d�n����ÐFoOs��>��6V���X��G;
��ߑ��&ϟ�!�:`>(�wݩM���X�����~ʅ���Xg1=C�7386o`��G��A3��Dp�HM�o�-����c@�8�,C���:����)z�g�$�Jd1"bb��Т�ֹ'�vI�gu�R��g��z�\�� (|AZf��I�!�f�Tx���>�	���/����������e���|�S�"��l��,>O�5��@��4��L؆�O���Q,F��P�W+)8�`?@^�?�*>��H�S7�j��)�����A`z1����`o^���Cޏ5����Pa8�Jy��~-�&7��4�qd��}��+sU�������I+N$�/�_���t��C�-OV�{n
����=c��ETZ�����H;��Ӷi;6�/�u��mO�U�D<V�D���ߝ��n�P�s+7�FB��]��2�7��7&⣯�����n/�wf=�P7��Zg�VGdz8-�0��#q�~����ܐG��9U�Zz�YXI$���*�h𓲓���qCf�ͦ��{�!ǷS�s�5F��7�(l��7ʝ5yݥ�����޶�t:&q9�6)P����2�c;A~?�<��״���6`�/�q�$����i�>�z�!���<�W/$�[a&4����/�%�u��N�����I7K���j6�Ĉ�;ϖ���c��>��W5m�υG��5��ľrJ� ��V�4gQ�ygC{��ǔ�)�j&��Œ��E�ͤ�-��hဪ��k�r�6���!�r����r=Ἂ�m�8��=��ZGA1eW짷�>+���[�,�V.:�=/9J�@T�g摨�Y����=-X��j��~���٪#�O2flg���>��F��_���=�&%�W)_��D�1>�)ɂ�}dB�,&��p�Φ⪨#����"��"�*�ȖPF�(/��ꌝ����C� *'Ϡ����ە[��M(�n���~�'-_~��w5�����nɏ]̈N~Z;���s�I;��i�)�ə54=���iZ�>�94[� Y�gM��������QMj�������+��bQ��\УN#��2WR���V��\v���~��G>,�p�M�F������u�"��N� ���#ȵ�`=s�#���D'Ȱw4�'ثx4���eeo-q�4�X[rxxO8((�T`:�c�);n1>>Rܷ�%��Bm�ݣ��*�K�[����[~�=��X�{����<b��x<�O`��j�/�
~��X�3n8H�r� 㭩x+��[Jꔋrp��^F'_p!�Kkh{ֲ���ܼ��Y�Ї��'�ț[�z��a7v(<t�F��k��+ƴQ��#w����Z������L��2�M�����%7f�#Z�Y9�ۍX���@¶����n�֯eu�!��LY�G�9Q�G�p�Yx����)5�D:J]��I��O�ς��t��ej.0G% )��Z����9.<������6����)�^r|��C���=�I�>&�3��a�����[�<�ځ�|�:��n����|���o0��O�X[��1a5��^�{z�Z���)l s�tJ��
�B�dw� �hH���ݿ�<;#Xn~�����Ł0�����d]9϶!0M��]�U|��`A�c-�eFvCv�S�����+���y�ѧes�/��%e�� �3�#����2��Gzz�ྋ�9�����S�*�;S�AX�V���y����Zsd���=߲��c�K�<�_���,�c������k��Yt���C<�����=w��q�[p�
;X9�����?�ړ���ω�$k�4`�ƻ�{Z�3"yxM"�/�wv���$��ڝڧ�'�U�Ʃ'������b=�V��)�z�)��7q�������v�T����1 ���}w�&��w�[?q���6i�Y���^�0f!�Ԛ����+u�-p�I#_q]�S�R2zү[M��
���ttt�	dS��Ir�+U{���J��2WKU0oƽ��M-����Fk<ū,��6,Rg�0�,xw�������>�2�i�T���~� G\=. cmoCY>��Mx�g��-��F^�����'����nW�w-@[�M��LS	 ���/EuА�ٜ�VT���̸��x��&v���$J艸L�8��k[G��ddW�������?����nie�=��̒�9}����ƌ���o�η��/86�"�-:���,2-�ߋS�����v��xW�����eH% G����ėQ�1[W�l���cN�,�%��֚�As}j�
	�!`D���m�w*��axh�,����ͻ�������T1�U�{�3'��{��^���Ə�؈� i}c&���j?^ח��O&��[�I]�q^�t��u��4�S��'�b|#��9��� ��������D��v��	����ggH�	n٧F���?�l��$2A8������2���Ҽ�������5Y+�^|ƪU&x��}�@B�����9�����+E{��Da��5t��xIu��I����7���ټ�=곗��f߰]�����[���+���?S4T���Ϩ���V�H�f�;�j#��0B8�9$���Zi��U`!�yN�!�@"TÀճ�}lJ��2�kWt��S�N#�;�XM��ž�t��=[��� ��~-e���=t��뻟���9�{����%Tl߆�S��w>*Yl�S"�8�q��=��lQ��Ԃ(��0�u�?aZ'��h���FE�<�D�� L����|Q��ͽ|C�^8BV�v�
�������2w�;��3��Z{-}E;y���V�����v�{�u�q����Z(� 4������9.!#\k@���cI[4����ۗ�gQ�Ry�_��%�/�z~���A�@/88�+�z��i�� ��/�շp%�5����16Ⱦ�5��acZ_���(������z�U6������X ��R^̵�%/���?��oi/K��������7Z�З�䭫Q-o�����	���u��T�<�K�#Z�7�udcN�[	�;�e��� ����ں#�����bM��Q?�m�ܟ�w�3Y<��ZP�I�I�(� ԗ�b�� ���b�3�7�Y�|��$�#d|&ty��/P���c�� A�뻏�m�OY�S��oĳ�v�6"�6��[Bu"���C�*�ّɬ��;��H_|Á�.�m�W����ϼ�N�Ww����Vi��D5}������O�YƖ/%���_m)��ӳ�.�7ZΪ��=# 
�!m��Q�/�AK]k�NRG8�̫vC��V8�:�
䃒���T��XD?H ���0��1����巓��y�T�^$����gy�"t��g�F#�459>r����l}<]��oy&�tW���C>Mzs��<�s��삹��+���T����i������T�����
�{�h�]@����`0w��y��^2��Z�jv1<�<C(�.��E[�e�-��T6^ؙ@���s�L�7�}����}�,�N�<�@Q*(�1|t=����&jtU��;���C�-����]mK?�V��ܞ�D���ez$�z�J꟤�=u�T��'�
����Vk�>�G����6j�q�ׯ���i�PH��M3)=F~���B(���$s n�G �̟d�_�&Z3C�"q	o!��
%�V�_0TPB=���l�pZ�Z-O?�� ���M'-���,h�҈�W:�̵m����eU/XD�Ծ�f.#�	���@�ZU3��»��|����E��uٌ�ܑ/+b��ͳ8l��u@@���:�f:?�э��r�zS�8����{���/G����s�v�'�����Ĭ�ȈF�
�aƇ9�.�c )X�)lW[�����S�Zήaq��\d{4�Ε�ϓ�c%at���7��S��t�zW�~�S*f[����C���|������V���a<����167��fh��v���Z�d�c,&U���uK�k&�L`��,������:�8V�T�g:s6F(,��!BZZ���2R@Z�<�B-Ɖ\n@�#^!�?@��<�s}�k{��G�N�P�[a�Y���L��bx.117��$~��J�Q�L-����zD�c.P���{oyMn�'q�?���Z�� 0���Ů��G���ϳN�g?DJM���$�`d����h��G����,©B�rlǱ�Ă���E�!f�שbH�<{��h� ?�Bw?��}�si�i���鬯p@���T��"h��KB�<�sh�[�o�,�%0�
3r[�U��";�
7��_����;+�-�z7�Q���3��n�kP{#J_w����b#76<Ù���"���� ~��Z�����*5[����|̙J��{�+��*���)Z(P1�;'4�NS�o%bW���~)ob�­���=���0tk.�A��c�/�Ҟ�ONr��?�<��������|��Ởh8t~��y����ƍ0�0��`�o]��i����ueP2;U�������)m�w���ּ�&��MMsVg�y�MK���G$7����� �)O.R-�7[w�CH��x<:�C��jI�U��JY������z�����-]���!$5��o%
�idc���Ncn�;��V0rS�GʻŦ��S}��AH�~U����Y���Y�r����c�X$o|<�(���\*��v�;'�@���c���ί�y����F1]�f=5Qʖ5�?M��s����D6�G_���Q��ݚ��Փ�76�� L�6��K���Z(���9�һSA�5�}�ɏ��I�#nF�x�9����gn᣶���W�(�p���b���F���p��K��R��Jc��'��a�Hq�"S��g�{�f��c��%���6����N�^Sϸ~c|�R��m�<�2��D~ÎCG)ɫ�CmH��;x�7�>�]��Y��[c,�4�/�35d�_�#P�8<�Ό��^C4.�|��� V~n�(>S�W'>95V=6�ɟٸ���%"l��e/�N�#E|�q[6�y�,xz�6D�&J�N��9�-��ȃ�r��_���:�d�%������p���g�jQft�Z�@�V����ߑ�#�6$�`OX��}��Z�,��#�铭]j���5�;$L����!2��1�EI�
��|�{T�w��%FQl�)�ۢ�|6��冊C�|�T3y�5�êTM��������C���r�V�7 �?��t<�m�6�l���,�S��T �jվ�݁&}A�<������N���	��W��O/�غ$�o�,�W(ϞJ�m�
�#��Tc�?kW˲21}P{��:������[�Z�ْ�dy�"�P�Gq�����W���<�|��,2�ng�j����Ԕ��h#È�L􈣞�#$��
[��^m�>Qi_�d�J��:Y�� �5��#����5�g@1���Im��n�'0/G�6�6��T�I�'oT�Es�iBl���s�������4�iL@-��"e'��"�])�.�����fmU0ޡ'T�ٷ������j�x�������xd��MSj$Û�;D��`�l�IiTY�DѬ��7�WzI�ZZڈv�m5���3�Ao�H��%&m.��+�>�>e�h�!.�"eG0e��3E��cD_���u�䃓���iG�-���e�ע��A?�{{�ISBo����m�fU��6��[Mi�>�`�o�&[A, �ʇ��x:��z^z̹�.S�S�S)ڍ�ݓ���j���ۘ4��&L��K*��\7����nI��vM���x5��v��c�Z; �M�SA�ޮ��_��S�jr��k�;]�F�o
k�]��_�^�j����*t[d�.��DU{�\�z�1�ӂ�ZB ���
���^ǹw0p�څf�*6BEa����g�����OW\t!����Ǘ�/R{��=��(8����=S���7PN��E!n�a{4����Jl�a��?2/צ����u�H�x�?"�rlzҷ7�p�ld�(�җ� �ﺁ��
� dFp[N#	�W�
6(�F9Ö�+��ht ���[S.$���I���)�(��x�*(_]�����f4�h�Ǽ��K�#�)��5�ll)-֐01E�я~�x�2^��=ON����`�m�1��� ��Hp�-'\0��C��]J������Ca�Y�:�ɷ��@�Ab�ꯏ @�m�q�1Ϣt����JE��FW8n�/�>*�ީ��k��dy��1�;�m0YX�$��>�h\��侏����W��%����-lxϼZ������Ĕ��XYE���6�i���w�O9J>��}�f_]�FP�`Vu�5�b	�5]CDkg��1U����>��D�@��Փ����Uj�d� (QU�Þ���V�⠟��1�s33�r
 �5�^��J�]��B�񏹵��TN�o�H3�w�'�>��~X��F&L�T�0&Azʬ�+T��Bo�$!/��F5�k~24M��;P���B�X�ēb�� ��9$�6(;�}���/$l����K*�o{���E9KΙ����|/KFSBbrr��]��*E�i"8Mg��tSC�;+	���t����1��F�U�^������̇I,=��Z���j#m����T��g�2ebʡ�#�~ˍA��C��K�O�S���[��m��<6H.s�Wb�>���	�~�>��E�7Vl��/*�e<|Z훦�������-�8Q�W��5�r�_*e��8Sa�|8Yˠ2�c�rޟ�.����f�)�c����^Z(�IU���Sꗻ�C�	����apa+�ll\`\���9�Ĝʦ�q�'VJt��9���=���տv�W[z�a�m]��6}�^�˿�aN��P��e ;�5:�o�Zw�w�.]n�T�\Z�q<E>�x���k�@��3���P+������Mp�[K��Eg�x`�=�X��Eȏ�Ko�U����ؔ����n?ۋo-���r��-m��ߟ:
x���n�J��1�qqkRc\���;9�[{=�kw�\h�l��j1j�~-�_9.�E"�3.��[��n��n��`g�TX]h?�%~j�?�zVб�L��_� ���̬��J����{�~���=!���:ۺ0v�U閺���I��ڍ���1���nsa�->E��?��㫩�ٛK��E�_rJV���f[��ޏ��&O�^�Ɩz���)����i�p���&�$th?�/5\�xK%D����>���S����|+���c�M݃��$+/���j��|�N-ՎY*���h��t���tn{f�ux}��	�Vn<�+}�rf�0�2,�ꊮ������{ё�s�e�|2(s'p�rҬ��w!{#/k��	�eդɳs�ݍw���S�q�b��|���3�V�R��U�t�p����G� ��XdG����/lI�]/�׈eك6�J�x�r��	�����/��j��Z��d�J����v��f�R,G��WSN��<E��C�Ƚ�{���i/HɷOk�!��U0^E��6%�oӊh&����0~P-���cǐ�uW�ש���o�t��"�N�3w�G�%
G �{���K^P)���U���j�k�0j�1��|^�ڈ�-�_���V�e�Ε�M��<��.g�!݇�D�b��x����Q��m�ZQc��[_{֦z�U�ʿ5ldR��0,<?��쎵{�q8F6���]2�am7
ޢ�xW�q������<���Fu���I��ڗ�����CN���[\��� ��{��؆v
��W�U��l��y�j�g�r�HwXCj\����"����uS��!Hc/����B:k8!�֧B��x��p&���QF�����}���E���L.�x��ir)� +��ᾯoX�\k��k��=�A�FZ�Z����ٯ'��k��i�z���Y�k���@	�'{�F޷�����'�V�RN�d/<O��3EҧŽkK��	�a^��9�EQ�}����ʢ'w^�=�/��q�$��[�����B���\ؾo���Nu�(.�^.�н�����\vy��6�����֧�rv��e(�,E��T�4b���W��%o!�<ﲎ�_c+L�d�j��'ҵo�!+�ff��ETp?����mυQ�b�R��-��{yb���B�7������I���K/�h~5�Wiv^^����sf��"�[����K�ם����p1�76�N�����9*S�����Af+�X�`8E�"��V*�-y�R���^J��������������!��z�ڶ�8�aF�5;<rX��$�.j��m�e���jw�Mi�+bO��E�#��k�vM��^d郾E�[���ݔ�~������Q�F\�:��vϛ�qǼD(�੩���������y�5!��p�x���Vc��*E����L�y�C����=V����E�������a���x�k���[��F�$E�I��d���|��+���{�b-��{?t���!:J��g@����l�i7�j�v+�����I(�������ZN-��@�k3b�u2<��չ�}�@
�K+���}��7țE���Gܐ���q^����5]��t�^����'N_xAN6��<':��DI�ْ�D��!0�����Pe��B�[�W]+��)P��^�u���,A����ޙZ����G)f�=�w	2�ȗw߈�W���LF�N<��QƓ�lZ��?Si�p:�C� ;`U?+�H�O!�>�.�R���}�P�ݱ��~�'S��B��&��HT�v^R�(�F��9��!���z�e5�*�_���DtuJ����z<���s�UK�W��F=�zB��8�1�_`;_��my�h�'��+5ι�ޖT�2�g�ms�q�F&$_h���O����_ך��?�.U~���u@׿k`^�?���.\��`O��w�}�az��x�U��� �[��lU9�z���뎸��\7���{�9GyQ��x֟,�%X�q��[���H��o�|AQ[���;h�ߥ���s�3p�^��Q%��&��?�S�)��&a��r-��!&���IK��8�LeY����6ԉw.�jZ��jͥ4>kx���mȻ;����]��?��u:� i�ᖜ�v0S8S���t�F��fƺ�p�l�4�w�	�G� z�:�gm��<��j��z��b�r5�r��^v����x8
Ц�j��������הy%���л�e����4�j��w����A��[�lC�'ds��S��x$���qKxώ��R��.�0��ҹv���)�Ia]+�ݩt��Y�uO�L�����x8H�_V�xk�zfxR�%FI{v�_��&�i9+Q���į񔳲F��~� @B2�)/?֮X�b���,M�NQ��,Lu��e�%M)t�.э���w�n�*D�M�����قc�I�E��"psH+�i_PVVVE�8e�G�� w^�lry*/(Ǌ����Иh����Jn�I�J[>��l���+5��?���Ttu��T��ȥ/�	y�d"���9 ��X�h�h��2ڗ�Ʀo�e
Ξ�k�y+�5w%1���_���"� �-4�n��,���bd�o�q���v���9��WH�g���JIwz�޵Cl���r�����O��(�5W^��u�s��Ǚ9P�j����.M���8��6���������0�G��OEo�-�iA��I��n_��n�v��8w#HD��J5���h�.`=�ߦ��0�Ey���y�����2���Ԃ���fm�����L�>��lw�5Ħ��U���DZ�|�>E)���ջ�/�� �����q��S�K'x����E��Y�F�ۀ-lϧ����J35��O?}�~���Z>�p�Dl���[����UД6��Ǭ,i�QQ���;;�Aϐ���A�X�bm㢎��(m�D	`ޮn��Y�2��vx�W�"��6 {��L{GJ��_�{M���5���n�|�z�ͧ�Փ{��7ç^��!m��)|T7���ƌO7�����t.�g�鷊�fcPw��ysӸ�2?%>��һ>9�^�=��r���f�0�9���~֏���1��Dc�'HHxw�Z�ļ��ǥ&C�sSE5�&V{6�t�Stz,e�aa�)Pgki�jX�W<(�3� [�	��{�TLƱ���"t#����,�Ȯ�zV�{n�Y�lTU�WW���3���⩜����:�/��O��B$x�#�\�{&�2��6�e)����8���@�~=�H�ކ��zo�5�����c�Ґ����)�8� ?^�AF��wB�C�G�HH�;.`�+��Y�����L �m�%���U�&�53EL`�1��	=��p_<n?�A���J��7/���rE����ii�q��\h�'G�Ͳ�1��Z��u��[

`lk5��k}�����Euy�$�8-EZ.��~�K">�bt�JGf9��=�`�ǋ�*��c���n%Ā���F�}�^8���K�*����P����,������l�D[���EM�?��B�ڼb#ldڂ�.g��2��a��~	��w,(�XH"OH;��"�VN�"bL��K����0B������oE�I�f�B�Q���c?�.��_��c�/?)�}]� ߼�+^��z��	�H�x�M�@(H�y 7�pZ�Ԭ�0�FO-�<����5������_sK�^ϭn~�����>�Z�ȩշ�M�.,:����,�t��Z�ٴהP���MBf�:��]�����[��+�Z�!(z������W��Ojl�C�� ��3�٦Z����ðA�dJ�wm�қ�t��ץ�������p�s�Vd�IzȒ;�����PR,$�:��s^�L.E_�G������p�`_.n�B�J�7��V�ř�'wj)�`_�^QR�����Gg��Q(Sίj�b
W�D����9z$��kui�Cb}Oo��I�g�W2~�u1�6C:�E3Bj� �$|�1 ���l����9oٖ�m�p��a��:`��1ۅsYM��X�w �"@ދ�\�}��.�扏 }��0ac?n����9�{(D�͠�Ak�5�U5`#��D�kV�Y�s��צ�v��������h�4�F�F�ɩ��	�jTs� ����D��,���$Z��H
�ϵ�>m���W�(��ok~�Q�[�VՓ���}���'rC�5�w�ۚ��93@3Y<��B:��L˯최#�� �:BU�W{	Ҟb�I_�JXx��]��QL�u�]s��!��ł�xDtohС��	�:_�j�R1���c낇e�.H�-�jGn'<�P�)����#��_7}��h�%�lY9���_��+v�]���#$����	V�2���r�3��=F
��l_��,$�p����ža��Q?�J~r��O9S�Ap@����)ߝ}��KE�?��.��q�-.�Rr�Fc�x�oiI�d9F4�6	2�ݘ��vw+�տ��ũ@H�}S0@_+\�7g�ȕ�MOێ�`_O�$Z��R�++�i�0,��ظ� 5K6��v��3�ޜI���qb � r�.�����?�l�iU�;���u��������F�ț 5�Sjw]\`%�����8�|�����>9=�^�^��O���+=_+zuqc�ɑ3���/i@�N�7'0�vf�y}�d���NOZ�¼~���St�4S��?����Ts����4��l�PH�$�u��t�	pP� ��~ј��s���nh7�����*x+���j�AO�5�jŔ��1�w��o�cڟi�84��E�ع*9��;��c$H���)��Aj|~� (j�X�Z�yr���.m���ZJ,��a{8���Aff/^	2-�s�]�ԶS����/��6������ &��pY�� 46Y��w��D�*̉�	�K+a��A��v�E��VG6���I�(�NO���$���R�<� ů(��x.'�>�Ep���}���B�dW�!b�7�d)�4���T��.Z�����Mo�dTO���K>�;�a��g_d�|�ۺr�U�]���M.�R.B�C1v������TG�A�/hC}�bm���Oߖ��F��"1�+�
�u��"�M0K���6��T�:�9ٗ(b�
kfI�I���U3�^�.!�6Y]���E�)�"g�6���WЯ�E�lf7�n�^��Y����?�$�@��Bz%b�W��	�\(�e�k&��HL�|t��J���Dr5�}Q2��{rS:95Q ��2`��T��(ø蛀���J��c{w���XDJ&�Z��� MM�˾��&��Md��D/�պ�����|j!{��r��	"�0���,�g~�a��[���zx߾�|?��ئ��N���ϒ�iu����gb�V$�����,O��c�ɍ��)����+��_c�*!$;bc�5H,���J��L�w7��~��y��1�@=���܁<����^��[����c�>˘.��sB�^4��\�먌��CZt]݁�����	�zE�\D����n����s��̢� Ӯ�թ��_��8����� ֯��X�_��4���i�1{�s�g��Y��i����}�1D�B0����.·��g�E�B�lJ��a�2y�i���r�Pl�0].mӚ���;e���dT�Ǐ�Z���Il�`���Wߙ&�J���5`�	+��@M�Ҩ7��P��t̿_��A��
�;9M\�zO����lO��[#�٦L�����i�� ��ل�h(Vy������ ʾ�3�s�1ً�}Ϗ���S�_J�x�oo�2_J�Jdrr�[�VU��(i
��Y1�n�!=:-�X2F�G�:E<Ѫz��sV.aJ#	OcVǖ)�#�,��U~�v�����&k
cW��F�x@��t�eg���1��Z9�ze����מ�%
��K���i�z��T~����w�ȇ1��5H�㽄��3{l�$�.i�y��Q�ZA�댤�"�0K˃�>G���__�0�eoG"ٔ*|���bIX���Iؠ0��s��oA�ڻ֢�k��y��X��Y����",��;m��Y�"[����"���N#��1����<�v��}NH�9�-�_��Ύ"ɦp;�b��r�)�۵�T�N������m��dl'�eb�����U�|�]4C���M��.�l# �ժ�q��dv�$-.j����%�cQ� jr�ݵZ����z�a	���i7��l�'�ͯ�9w�9�M^e�3=�Ԃ0;[N�)��{�������򌲜��Aҕj�m����u���W�I��R��J�=�j'�t�����<�R��^�w�2u�A��Z�P�A��g�Њ^}y)�r'9s��.l��B4'��Ѱ�1�g&U��J����H]U��]o��1��M�2��.���?al���B��%mӡ��b��Q�����+AC��Ȋ��9L�8�:9e��r�!�C|G�p9���m�^�޿7�]�v �v�t�z�VN����E�� Z�KEJ1������4�|���T�G�2�,	6�ʶ�뎩z�M�`%����wt�JwBN��������C�Yśs�q9+$	ߨ�2�ӮSU�i��{� gg�̩F�]b�C�^^L����3�J����%�Mp�מ17E�#Љ|�j�j&�����[��W�a�Xے<�s.�. _�zB^+p��{g�Mˋ�L���X*�����v�WU�����;l��J��<Bu� �AvgW\������T�|L��8��n�=�n�.�H�IPzp�l#��U�TEB���9��z\��I�V���ow���k���WUU���r\[}5����T�!2V4��ˌ��n `δ:Eo���=�vVB&a���.c5��]���ۖ8�*RVψ�
��nLiJ�/#NUu��Sy�;E���dWY����z+5�uig)�x�R��;*��EZ�� �=�yՕV��d$�u͋��n��RˁY5���:��ye�#b|G��ޕ��Z��Snk���;��
"Zl�%��n/O��1�@�{�? ^��lF��-(G��0lFB��k���d������t2$���/2�E;�E]�ꖩ�6+3ص�fG�uq���;M���%k⒌�I��l��[LG(�2ߗ�5�� PK   ��!Y~��a� ٮ /   images/dc707dc6-8489-41bb-a5bc-77a0670f90d6.png\\\S�� Áh���P%�lٲ�LX��,��
BX�Q���%�A@�� �0Leʎ�gb!��b�����p�=��y�sB��#=�=�{ /��E���-��|��@�W�]~�a�<����7x��粅"������	��Q�K��&�����N
%�����p��I���%e^S����iP��`ȓ��P�ej�l�{�y�o�!O!rݢY��بߚ愳����}���r�Wk괡XY?�q�?�üh���!͵�/V��xt�e~fc��	�O��D�:���s��;%!�E.�o���˘��P\hV��rɘ �;����TS��{k����EA�n�Z��2���|��k$8V�p�N���$&��������Q�9�HO�	��T�{���M�*��o��f���̑��M�<�!�f(nQ����P/ h�fvh̜�,`�*�Kp��e�Wc=W*&���s#�pSx���]jr������Y�]`7�핮��jʿ#˰?!!�\Y0jn��D� ���Ȳ���h��87Mr�q|h㡴@~�K���g
�	��Xy6\���J��ځ�ӏ�u#H�u!�}��K�����%%%v�ou�V'���'���$�
����vv:o��Dz����p��r��gD�*������Tc����u&�17Jw-16������p%�8Ec��Nl�B�{Eُ��^�LG4� �s3�Y&Gބ0�F�٨����?l�HIƾ�䦚 Y��q
؜$ȁ�,S���fDz|�e,�q��傆��Vn����@>$2�r$t-�Q����a��o!KʐĦ���H9�mb�����m�Ž�u_���is��=ۚ����1�r�|ϐ�B-a9~X
j�MD��+	��#ҍ�֘	��1//�����")�	p[�e�5���(ۯ�N3�� d�)T�����ɂ:�x�f�h/G���%�����	L�e���fx{���}~~~��J�1Ε6/c�&�
?LDD�˓��3�{����g?�eB���Qsn>��>�2�+Ȯ�\\�1%^�+���q��>�n���R6��]�]z�}B�u\����uv�Y��H/$�W3�
&d��Z��v���#����ї����k̉�����ڱGw4ʂ��W/��� Ɖ��OP��m�*�E"7f�TU�����a�@���+���=�o�a5sTL̖=),�Ek�k�:V�[o�_�#� �zbўׯ�o��Z�Wud��x��CU/��Z��,L�s�ŉ�kY�����"NN�9�s?���ma�����i�-g�1����H$_g���d#0[��n�����S�Y� ���>snBj���ݗqt2�0�׏�΁J�����7Z�|�2��_���R�t��� p��Sй9;��q`;6����@��VhS���[�0��o��V�e�_|B���l\�Qq���So��D�����[�m�~��B��D,|x*.F�Ƭ_�8��J$�Asp�y�f
<�]U6��Ka����n�����#	,�~��=w'H�g`��w�z�<s��@���Y�Y��F���#����e^w ^*����&���'�
o��$5�8����j�����	^�,-�%z�h���K`�kʋ��Z��**����J`�W	����5��#��i���h!����6Q�#l\Q�¾��%I�>}����t�=y�y��~pyĒ;�H�Xc�u���޽{ͨv! C'����|SE��u@��;�u6.^��~pG��
� �ژ�m�@[�:�������EEE����G������b?�*���������6��7)%�iv֣j�kP~�Ӑ.�Ă���:�tD�B|{B�B��Ǭ�A���*�m^Y	R���_
�~�VP@���1���(g���l����ˤ�E��m6����@��:9߹���п�YL	�i:��fdZ�c�Z-Eջuee�KY]���mUCEUUF�VT����206.���J޲DvM�d�|�v�3l/��i���9����ϴ��Yy���3�;ǲ���9����vnHa��zC���d�?�{w~��|2����r��,D@���ͫ�P�[�kᅠ�,1z3��@Sd��o�<��Z�x��Ey��(韤�����H@n��̮��0���k���TM����PSc���q�h��m(�Y�
-!��a�؄c�o{�����;Ϫ lv�R�
�eXR9N��6��c�ݽ�j�y묬,�/����bF�a���؉����7��Bl=h����>�n��P�J$�\@���P�y�m����_g.$%'7JTc�e�NLִ����������=�g�'?6�L��U��N��=��g�j4B�- %�O��@%���7U+D���oM�"\�"$�p�� {��+#1���G��P������G�8�f^U� �!߆P��ɲ=�Lb�ض�>6ʎ5��-�m��X�7�E��EvQ�K����(�����- E��ռ�*���к�01>�s��� ')���.Nb��̔�98�p@��b���w�X ~*lD���w��-����B�@�=v,Wc��=�M//Y�o�+����R�U���^_�&�}0sD6�h�I#ql]E"k�뾤�bS�4�]��IU�l[�I��^�7���z�5M�뱂��@��l�wTh���8�4i=8�j|�ߛ�8I��
��$�
�}�{<ڄ�o7�C�+S�$�qU#�3�FFF�����r��ၞ�Wz1��c�N�M�cQ����}�".��O����*m��A_��o
GϚ х�ie	+��dH����Q�kE=$��m�2�0E��趖�`;���8�31J���̧(3�ۅ���w���J/�:��K�\��"��PGe�m��=,����Cj!��W�cVXU��L||*�'d@��������Z�2_9�^uj�B�.+��!1���RݡY����)�&)>�B�פ��HkU��k`"�c�/�oS"���ʦ��6C,��x`����vb^�p�`�Q�Ǔ\lsDY�x�,P/}��r�-i���Y���5dx�w8���t���6�#�q�n:��������f�de��=�����Ĥ6)3=A��\&�x(�EE�f�z�����FWG�l�2�����0�㥒���E�i�^��QV^*S� B��Uqк����P�zK�'T��I|���	Tb�&��S����<��51��W�H$5��(�>nV��*
x�Nh��@�/DDD�$n�'5!����<y`3����l/`���O-P�>��-4�һ�e�U|�\�
�-<idd���v�Çw�����<��[��Fj�f��������L��Ӭ�\�:a���E��)hȵ��Չa���J-���`�[0,�)����
\[��&�,5U�����JT��;6�6	)���/�^�� ��gz�s������]��`w
Q���J�����>abA��V���rkʳg�)��:�����wL�^����6�� TT��B�b���9p٫u��ۭl���2��C�uX���_#	���ڴ������c0�N�����{�����J�H�(�aԏ�Ƥ[����ϧ� T���n.I������;�F)rh���bi�
�Cܝ�޽ks��qF�G��W��9�o/�W�Rm�F������'�m�(&�M�h��z�4�0��z�n�<A���(o���]��4����a�<�$@�V ��om���Ź����+X��H��ޜ��P���~P#ʸe 7�v/��k�4Tj��gߝ���8D>a.�`aiY58ƌoP��UO3���f�ח��/K�j�n*�{�� �@Bv��πn����w-9�E�mL����S��0��/.���WN��_��H�&X����Hnz:�:;CσT�����ׯ_����ۧ��V����K�G�۹��K��>-���f懧o�v5�h>@��'3�a������f�ֽk�mv�G<�S>s�С�xĪ���J�Z��M��k𙅅�)����6 s���1K�^��@�z��ʵ�*�P������"7�rͽ����S���q͹!5`*�/Nu�n8�+��4`�0>֤?<������[+�/�?^\{�9�F㾲�N�R�������d��Ҳq}-kS���sֶ&t�ߟ���N rMJM��Q(:]|��}J[��r+�G�	]�E��]\�JlJ����5��2���o+���T���|�j�R��F�Q����v�\x���%cn&�'l�nP܉��X��М`��C�����Mq�ي�@hz�`�KЪ�,��Y�{�III�2̭mlFD����g�*,�3�=3�X�ؠ��i�y��0I�����P�0�v��qUI��.zn�p�f ��a㬉h59�f�~�P�`(�	��D������,J�`Y��G���T �a���c�7NY�{��S�;�e����3lgL� �s{N�>����$�5NN�Y�%@X��E��A�L�`��``` }����?}��xWt,		��8�
`;��	,���NM��W�^��	�`��v_[��xK���Z�
Y����W���eƒ�@�;���+X�\��XfyTX���C�꼩�o�gwk��oS��I�/����ơo��Y��Ü"1�<�"Q���_�|^�����TSZf{K���kEӌ�'�2j-o����������n�9��ھ��(M=�%#T�c��
V��%�!0ܲ�ܜn�*�ӛ�|�`Y��� ֓�Y�?��-S	�t�&r�K11R�Q֊ ���V )P�L`�����tn�O�֏�#K��bmY���Wy��`�:��#֌mpE銰ʗ��1�!'+�i���>��Y��tT���@�`"k[��%�2����0�nG��L \X�x5���u��4�3 V��`h[�V�L�ri�{K�Q~�E�1\�7�LykMU��+ �Z0��tʷg\Ē�ءj}	DrL�45SY��]�i������B�,B5x�s|�����5�!	����jz���?���m������	�X���2�JF�Vh��>���`靵�_X]��f%��}vu��o $�}���6��r5q /,�Fy��N���<a�
���xS�K��4  \�C5��r��/7|f�}�U���ɞz���Z���Y[�]_�ե ��߿GIlMȌ�p@〩L_�0��r��џ<M��}ZV��5RO8�t��.�@�w&E�_X�Z�T�,,\[����@�W���M@稠`Uy���7����h�b�S?��G��B9����~�e7��@�)���������]s��a��Z�u�z�$�{��$3$�����COh����ۦ���i#p���&J�!�;�\���f?i������E��M�gj��7�OH��d�rйN �`?�Z��x�%)[;�n`����O7=����޵��Ngg��_6���~�rq��'&ZӚ@S�N~|�8&�v�'��c]��K�W��1��4r�	�\<7��Z���߯�>��X���IFݯ�mۿ�l�.k;���!	� }	��3�zr�{��]�"p���2X]3����5�N���K��-��ɩ�[k`�Nͬ2�PXo*���r�y��P��M�A�Sk@��=d���*�D.��'{�Hl,��A�� *��.=�zs0̑�e�oQaO2@���U��o�,� N�wG��Q�'V_{s̰�Ƀ���6�⥒ң��������6�@ث����#|pI�e�(��	8k_�g���C-tտ6<�'�W_�p�ڡ���YAM��&�jSب��}�_J烜��X���l���S�n�%� bSk�P�1ߟ �he��X����<��7? ա�8��J���X����k��<^㲭i"��۱���S�A�M�T#rrr�D ?ы�\g~�(QQ�fV��O%���,6腟g��K`��<���s90���4X?�B=����/,���~�2y�a�[�� /Wל���!UY6y~ڴ���4$�J������u�g���W�}�8Q;^rݹ���%ǟoO�z���U�}�:[$�p���y쓣<��bmi ��������?�m�-O+�T�X�������u�2�xs`p?@�C �c��B�R�m`��0<ˏs,O�V�x�$�C����c�'V��[S-��K3�k?>�Q#ǧh��8~qnC6�������\K2�L�h��X��ꇶ�˓�C��Z�ִ-��@�Z�E�Y�v�5��1�ָ+��-��ָ����%��E�s��&��s/��� �mqwb�X�����|a�~ds�g{�B�DA{Q�Sqc������D�]���Z��,�)��y�X�O�-��<�շ$׏�i5��ʡ`,\�87�Z���n��`j�\�N��.��o���E�����{�ID�$6��!�?/"6{���a0Y�*�v��_:��ء���~�.��۠f��a�c���B5�:��ڶd� m��V�d������/��R�й	�����/P[uC걣���\Ǣ�H6�e�ϫ�J�PuףF�(#Fk�l��� ca��/x�����&�=��r���3�!uQ���{����J�>Q�ġz�h���I_+�1�L���C
�A�h��C��\m�&�O�j��P'�uE��)��a���������˾�ޡ��r��SbƢQ2�1S��ݐs�;n��D�m�Nw2G�Y�!ayO�O����dY,C~U��!z[��K�����p�<ۋ�|ܯ+��0�gϨ��m�az�	���5�{�RMY� �$�lz`tr0�f�� �G�v�V����:�_���Ƚ]�wC
������r��T^n�Q'���n-�xM�$�����q>!^�h9Q��c�@nא
�Ճl�n�_D�/�����g�k�a�2b��b\�4� �?�e�N맃E�D+����0�j3F��
vz�A*_���p�\�y�;o2nt��.x�9�qAa���}�1��J��
u����$��&ɾ?q�h���}Mؔ���2�����۬$j�_�[��A(�;,��+��I�7��A�Y��m���++�O��,�$�d�����ȡUFH��(�S��:U���w������!0��FͻL�5�=�g��vx^_�Jv���>e�b��Lg�V<=_�8��h��>y�0���61���j�O_��������@�X�p�:I�2�qm�/�}��RT`z7���[�a��V�bSL6��ˆҷ8��7�WUH�]t�PI��)c�1ùw}`��[��9j�:@����1h����[3d�����{"4c2/n�j��;�aw�L,a�p�`����y��C��c�kT$y��3�����8�:jR��e�	��g����`t9
׵=T��
H�w⨟(3֧��������Ĵ�1�Q&�m������߁sHw�7��1�	mK�m^����Z��rA�y��+H�b��j,NO�n�"Į�HJ����s�d��!}/��6�Š_@u��4 ��w��(μ�4��Ѻ�#*���t,0vRd�8ǗC7!�v��>�S7�ǤʑA\I�3?Y���H��U�y�&�v� ʴ�i[bp����;�E:��:Z#&��a�ua�W1ߒ��HUY����ˁb��D8�_��W��e�����eGL8_%���ȉ1�$oWu;B
�?�a��tT���Xm���ޮ��:K�pg�����$̺�w���!��vz<�:KΎE+��j����qj�}J;J8Y�r����B��t��:BS߼��?_�Jt�vMtGF,�*,C�p�G$]�	)���ȵH�͟�O����!KOz�ۤ�Wwzn_)W?(�OG��>-I{�N�)U:�a���;i�l�jw^�/�VCA�]��%�W�g ��/ӟB3��7`DsL�$9�U���er���4`փ1&��Q旗�<$�1�3��`.\e(��:��*���C���3��ѧ���"����N���=؍��%κ��
+R��8��čA�.���2�p8�Zo��tO�v�h. =X��	;�^X������`��G��v�����e�3&F@1���`�������A��;D��0m$�0������/�z�}��&���60յ�� o�v�O�*%�A��ݳ�bz��K�v^a#e2h�8j�O��`+��9�v����O�&� ���T� oA��&G 7;����ϒ�H���ə�Ab_@̏�h����J���/�R 4lg>����Xкщ���̋0KV���.�b�����OF/z��B�]��#v^��1�3�8N�N���i^������xЭ2��dE�+�v����@ƨ�(����H����L>����g9W�1�=��i�Ϯ��o�-M2��L�+uw�6bGj�� ���g!�۽���N�����#��h���!Q�!��w:'�ea��Gb�YP<���W���<���j'���@��c\��uŚ_ND(_�y�[&�O�b֯��p�9���-���´�1�7`�]'x"Rv"P�N(,�d�%��,9 ����(G �XM3�\�����H�;X���Z�ť����>l�W���y���?+͇^��)χ��?y�9}e�yZ�X��$��c�i� �S��Mi�}6~�A�)�����qh����!I)���	�1���9,L�<lL�@"��8�~Q� )vdd�*��2k�Aɀ�p��H��SG�����!���p�M�1��Q,SHCl�P��x��^�tG��_�6��5Ka�b��`� d���/���y�L
,P���0X��N�K�bg�u�B��Ǝ��D�������G�Mc+݅����8#�o�&�25D������jV~b�u�3?y��������$kY��y(��G�01����u���hA�0~l�����ql�ߤMݑ9��2$"�s�h�]N?���D���Z�#��������D��k�:�8j�yۏm��([y�d������]��z�����ioxԐ��D�6/aj�Dk�� �_f�/SFM���l��s	�ߐ�C	�C��v����V���2��5��S�|�����XX5tNGŮ��SE �O[mC5=����	1�n�G&�ô�{���WN� ����'$���o)?�QXH82y���g_k��+��vG�������߂{�=-/���fk<>�d�Obnn!_}����o��r���-�rl�����d��p[O
���kz�����P�W�/\�-�=~��4r�=��_������?�|y�TJb.��H�p�)k�z���i� �=Pأ�l�f�����(ͷ��)p�?j���{��۰<�j����ϡ��צ�g0������\��
� �|��a�b0��\�;,ƕ��8�s��'7��szr�ߞ�M6��>*�6� B��<��9i�N�}��u�	�%�ﮦ���%Cs���$�Qҧ��jm(&Ց�L٩fl=l���8��;ҾlMi����W�M���E+�zp���� �?2��摕2�����[-�Ӯ�_����B�{���W]}����E�H��e{���k��>5]�i�W*>��H�P��ݭ�G)TD>c��R*�����#�ɐ�~A�Wr�͸�x�_t���T4�/�׈v�����Ԁ)7�Lo唏8-"?Xͩ����o���k�w�'�y$2�����,�����Z�b�ٌ%ņ:��s�N�g�)Ƒ����(1�M��ɘ���Z�q�q�EA��{�a�}Y��S>�+}ͷTB�(��T��"�&�Ά��}6��>�}�;�JH}�[{�(�ϣ���%���[��!v�j��(��Y��__t?��;Xȱ"wp�+���3����kֶ0Bm�0����1���q2���@�����I��g3�"�^�NTŝ��������0ب���U�0D���7���aK�F�罹����g�+5j^��q=|;G�= -{�BY"͜B�ή%�,����^��o�l��I��HF2��-1˭�]����=�o����}D}7�����a�߹D0�WЍ�0ą��%F�9�2�$�ך�:h|%�y2������rYHJ����ڌ�)�鄲�|)c�쳻6�8'p!q[V׃=E�;L��K�Hi����Y�G���:��[^G#Z!)���Z�@8lE �^��r��ݼ�C��4}U@#H��*���Щ���W �"H���v+`�T"���/�3���8H D���p���ri�-h����A�� ��4<�X���k�0���u��A�]�<>J�����3ag'2��� �����V>����߯��m�&)�Q�H��r�L��� �g��;=�РS,S^��8Sg�u�G&B
 ��o�d[^�=�+�[z =��{���e�ο�Wj��fa%�>���ɴ��ڜ��i�*zC���Þ�x���Y�o�75&����];�:�
�ŵ.MS<�ͻ��5Lh��M�vi>N��ﲽ J��O�+[�¢θ�*�7�z���yv�%��a����Ӝ�P��Ϻؔ5����~��MDɽ!� ��0����~li���u	Z�AmȀ�sV_���q^���O����N��J3���#��m�؊2�!���FA�n>��N���df�)|z�<�>>��$��"rO���M%���&s���32�1�=Ј�����Os׿���v�ushD4�x<����H����:������-m�S-/M�/I�
�szq���f�@�M��X���bczg^C�:��/�����ʮ�]�f��0����U�	vmCѼU���D�U�� �v�2~��O�ē��ǡ��.���(銎�����hкL�_�U�်�G����^Q�O��(�pT�����]rf�	��Y�)CG���\�MON�&��U�Q=��ݯ_�C���>�.�p5)=�98X}N�󮺺z��R�vF�nC���U�lՀk��I��p�u7�u� ���FS_V�!Ô��so>==ݰ�Z��9��E����b�F��<�%���Q�W�W���f֝NlRް�E��.��ux����o�ᝨ�E-���o8-� ���t"~?���jDJ�D�qU����'������+���#0�3ٜ��zz޼'ѯ�|_�H��uN�������T���kB�(�PiӕCU��3)_ߺ��^��93���X����ٳ˞�����4�k�}����!ct�����1]�/6�a)��R��~�ʸw`��x���'/���.�����xe�n�miӓ�'999Y�$����7�/!6������N��8� !��̤�%�u�����y^�6��YNWE� v������jЎS8���dwGxCPl�Ӿ�˖����̳�u��8�3�[y��Ŵ�͛|��G�$��W�X��,�����ҥc�G�ʌѱ$F��F��,���ʙx�!36�D��gm>�t>���~��bFb)Ԇ}�kY����H +K�ԇ?���@%�@������D����-h��E�>��psE���"1ؒ��v+�����	�,�_`��/М!��h[5W�=x~��	�Oќ$��l�9�:"�Exl\���^���kV���o��l��:���y��8�G搯���3�9� U>W�٘�'#�>/>I��2��{>T��I��!�aBV�c�}��|�PݯIG�Q�Hk��Ʃx���=����h��������Q޷N�m�i�}���~��Ec5��ƍ��"R�?�˶����uO5�@li�4��oyL�Dʦ�vJK����9nF�[��{e)ڕ��������Y��3q]ۺN���͹�WD��
����X��̺W����լ�
�{�����+����3�cqM�b�q�[�o�}B��Ç�}N�&b�����7�Ż��8�+J@+��g�� l�s<�}y�=�Ϸf*�;:�<1�~?�*�)��$��,��(l��P=6�<n�kk��<	.
G}+�=�Μa}L�]���ށd1�!��n�>̪�s���>o��2h$MD���Dj�׾)	�k��o��?)�$Bd-�?ݢWg@b.�t�|�!:�t�	t*��L��s���Q��$f�79��&B��$&�4�6*�uZp*^`�M��)��aa�	�Esqǟ���β�J�vp�T!o��#�'h!����ğ�$��]���М��"?��-��k9`���q�����BeG�K+_(��8�����cxY>��1�O���Op ٘�W�b�PS���Vz����U�oj��uU�.�c4���sw{.ތN	��m$]����r�~�z�L����|�uM�e��u*��<O������L��11�H�3A�mUcz���HʎH����co��m�8�3��.�>{i��/�p���7��Կ�DL]�EtP]]$i���Pl`ĂA�u�����ԗOE\OJ\r�nN�byZB����\����Z��CS��sKh��9l���3�^jn�?�\���,#�Dz�#��Z`�'nPBI�S�K�'dRo�l��j`I-X�j�7�3>�[_ooR�n"ayI~.�%�����RNhe�3$@`�O�k�Z4/r gyt%Dr�Wf���׻(�,�VMryqE�&�}�{(����	����' B��^\��{8YH�[�$_Hf�{?��c�R�kL������0�F'��s������NIF���\{�����<�˖}�s��U��)W�<-��#��&@�$G(��܍��DP�B[��<��@J]{��T�B����ڢ�#83�镴U�tٷ��"ü�h�ZyCv=fӈ�5M���hő�ˋ���mӋ���/:uޓ+"2��PP6[ͅc[8�e�����>�~�������δ>>ӢEP2��|�7�w�k�
�}ө�y�p,���S�<����R��ܛj������w��_�T�B6�tH鷿[�XEx_\yų%UN��]� guv�_���4C��φ��o��Lm��U�)�@�D��d+x%������b��"@�lv�����IR�;d��!���^�����In�B��4i��S�6w3���x#����U�OTG0�Wწ��;88H�U.(U��k��搸�Ǟ�����l���k��sY؄@�1�*�J�R��^�"�/���2��:����5��p؇�M;(kH�������d^���/b0ݙs?Z<�Ry- ���������Ч�����Qw��Q���ޙV����I5$������+�%g�S�b���n��~�qe�(淞�*�ȗ,��!;R�ҿێȕHl206�XX 8Q���1��c�T5nӡ���ȦR�*��SӔj����:0����hI��2$K��$�N���>t��)��Sq����۷��={��u�q�)��~��%������=1��)�I��xS� G�-�?��pN��Ԗ�����4���,
��-�r�1=u�g���lC�}��E�u�ԃ�G7��i27��cҎ�{��Y���Q��&̚kW��ێ)�4]��E�{`Z=ǖ�{�7�NI��X2�·��D��t<H����%v�~�^�����S������ �X�v!4�T����c�#���4�-c�j��3�ʗ�bO֯<.��dT�DW�h�ة2��Ə
g�����=|��|�����l��|Y111A���n{�B�ȱc����Wz1b��j&��"H������,մ��`���Q���6B
�t���Kk;K#'9x}�Ћ�/�M�t��/��I�N	��xC&�Aȼ䪲��zZ��Vr��7����u�h��n����(������G���z=ο8geulnn��W]�>���422b`d���+27�,��I�5�-��8��[��K�8z�͹�-Ȱ��+�w�mS��l>ϣ*G]���-LNM��l�����L��Ż�����}�J�Q�n���:�d8j(�C�c��P����-��-=�% ���<YAJ�t7�݇V|��V{���߄)=�5 ���[8���|����]��G��Y���@���'�kJ��텅���r�t�(��[�| �
��:}j=��e��$�;��g&ք�[��?*
Cph�UK�UK�j.㯜��b֎r�7���}!Dp��
�R6O7�M�k �b�Z��9���1�{1��	���@*gخ
Π���3�}�iڔ����h/ |`S�,�o��L(][v��;8�J.�e�ށ��1_;�1��f�F��6Θ#����&�氯^�����t\#�qQ�|�8���Z�.������R.?�vY,V�7M�d|��S�5�C�M2^cb0���Gu_����d�Ӈ��F"�bccn�K|���_��f�U�V%E4�M�� �"��$������6VI1���|w�Zk��`Ւ ��Ix�F�#�}���m竾wa\����ڃ޵�y�!���dn �-�ڴ����@��=�p��al�n�������O��R(NO����[���=
m,SM�>���ܯ���.Z׍��:<q)o$�8�PTW_m?2��j'�y:;;�}�c���7_(o�z}2gI��s��Z�ZK�|�"�|(�^:�to�+�LK�?��tlJ�)0*<�l�eڻ�y�Xd�35Y�J~Rc� ��~Z�U��(o4lA5���\��G��)��$cX
!�����W���z���͑�G�U�%e����[+�ؔ%�.�}��X������VO�-�N6Q$�=�0�Qݩ��乸��;������� ���@TҨPu]к%vU�e s�I�p?�7Y&�*%��fL8 �e�^�6�����o�2��=I�Mxw<�7&��{��8Bҕ���^4�����<���/F3�8[;i��t�8k��P���P�K�����-����ص�<׿V�;{��; ��y^�՛�Gss	�U��MdM0�{����u�|��<�;v>�=�Wy��,����oyY[�n1uݼ�v�Y��	`��uCa�:R e�t��X�M���\Ȗw1�&6���[�����|fT)�JV��z�6΅��̱���%_��\���s�Yw�$����sz�������;R�UKi{� ���4Dt'����� ;(���*# ������FMf��o�z�0=���wz���}x��`���w[�|��xOrƥ������0��5s��D�1���rϦ����8��zR�⍺=���~f���[��� 5Wx���Ytmk)A���wK>���V3W�O|f$L�XD[9�������{��l^uҋT�Ƚ�CH���k�B؈Ɂ��.A��L�>bhH�Xl��]��ݟyް��D��O�(�^�Y��~�]���c���֯��%��e ����{翼Ɉ�/FQm5����'�$�``���1�ɽ��|�,�t�@������9�\g���h[� ��d���3k�yJ��D�"N���u��$+ל�T���LF��I3	�Ћ2\\�{i-ۣ��9��7�	��-ة�����t�q�ri
]�"A�ȹ&�c���`���`胭#=��O���T�=���0����M��#:)dǰ[���#�V�T>a~�Ź�#��m�)�	�{-O�ݬl�!�0��R,�N���ʙ+��`��w;t��.[���ϯ�h*(���((�}rr2tI�*�@̯�����JG};�����>�M#\�s�p��m��7 �-}?��vgؽFtm���D�쒋�3��ߢ*�Gt�����g�}��_��lՃ�=��Z�.��}�ֆ+����ߏ��mgv����7F�\H�@���n�{-05�N���I<��D�q8�7چj��r���1�9tD�s@��@�����q��SXӧ�i�H?+�~�����T��������<�J�"sM�;Q�|��YY�#d��.`������9�����`m�*g��ܑ9�UZw}�>���][0ӽ�yW�J��ִZ�u�<jӘ�o�.I�n�y*#l�<�&�V����9�L������1���.������7j N[�S��@��myfw��J�G�@���EF#�3����w�ҋ\{��5�J)|��;��'����K5�W��4��: j������F��	�I�?�jP��I�3yb��i����=`����/�>� ����=N��`��=ϓ-�4�����g먬��43�8ywA�뵳o��C��g@��� ��5ꔼK����8��qV�����o߾������>D5t�����R�e�Z����3���kI�sW��Ԛ�m\S`�Oف�(���1qq�CFY;t?ۖh�-����	B6q�ޑ��˨�vZ����S�G�� 3�TVF,�r:�1Q�������]����O��X�,�,�o��aٮ�ȇ����V�5]^�1q���!2=��S�<�z��m��jz����>��~� �G�qh>�u���}�j8�q	��2Qb��x�����^�c	�f\�&���lPI~!)O��m�~lW�KL��� d����g���\�����Mw��Qr,z�j���5�X�QAAvʿi.u�H���+)��� (J��CL��h�摊��59���S�@��000������]�wo��^�=���<�0�4hF�U�IѶ��n�6-�?��8��W�_7���D"l>��z_���XZZ�q�gb�y������=�v�c�Ho�J)%��9��$�?~�/�XDƮ�X9}�	�]@����.�����xY����r-[�eB�d�ۍ_��+F��]N:q"���o������ֲz�a��?�����Mֲ���U%�M���t�*!H<���ag�  A���ޒSS�ǚ�Xᣇ�lu!�.��N�*$5OQ�J�V8>�es����v�j��< �E8/9LA��-��>V!��M�~��߻v�ĵ�$��rv�r��$ Odyy9hy#̗�/NF�������Ϯ|��t�3 J<"�f竾�	�a��+1 {��oY?�$��$�Ν/u|�����U����}��0�����׾���u);U�%�)*::L�~�ڞ�Jw�zj?��Xc��p����S��9oo9�ȰT�|��Zeo�����%�d�qL�B�w�b��sm=�:�a��JX�;ݞXz�3{#�Zs::: *|F?�>����8��7h�ug��Yڥ�#�p�ͫz��hh�=����-rh�:����wU.~qcmMp��8�E�D]�А���m�?Y��Xp��M@C�p/�cmPd��-;-�bd�Y��rH���+��[��R8d�g��YB��$[8[�&�~�2�xN��x��N�<�ԇ�C��{}y�, t��ݞ��"�HK���嘪�h�{��?R��>>O��U���LLL@n  ZsL����I�N���J`�VI��u|����ś�}��|��~��3y����4}w<������HV��Q�){o�P�̮d�ۑU$:V�)#d��1�DI����>N�ؿ�����q�sw�u����9����K��۷o+�c����jxԝ���^��j���mO7�*��&Db}	A� ��'���l����Ȯ��Ȇ�_�i��9��	��.�7��H��h���R��ǌY��b@��zM4��Rʬ�S�&:�:���)��qb��O��Ƀ��>�d�r���3_4~��
���J�j
�
�7b=$��ĥ^�: ��,R-�S�9�+]6�s�0}o�h���r���g��X�+�5D@"&���)���ʎ$�����4��G��z�w��"d_�~M�r�xH"Le*���Y��[���-�Ժ�x��Kz��ri���������{.�Ba�7R�⩣u<u6���7���ɸ��No��6��0�0�<�X��MZ>�a�(
��Ȋ��2������N����P̼;�c��a�o��/��HXy)y|s���=�d��	�VU�K��X��-xWX3i C	m��i$	PW��dI�CF�F@����Y	�}�F%���:Н�*���&�m����|-�~�a�g�B �=�2}}`���M�^����0Raa�=Ț�pl��WͭF�8�ח��lh���h�Z��R�؉dg��S��]}}u�)r���e�s������6�!�M�f��ք�T��X���0.@z�`����1���0v�ҵ�2���T����j˶����SW���"N��P���S��A�k��z������;��謽��e�)��
v��$��-^",nG��TK�Dw��8ϝ��M?L<���A@*i��=1f%��%r�]W��@Zk�G
�:���F>�=K�!�J,t�.SN���:��U-��#��/:�F�n_�񵛮'N�ɱ���V1�P�Y�iW�۩��_Қ86A�\.'�=xU! ��N����g\��I���T��:�:�ם��_�#� P�e%�`���A�?Ra�3�P�- h�4d��Fg�KS�y��^j�#19��=�R���8�d� ���{^�m_��3�$�c�|�zu��7���C�*wBBT�aůݰ�21XY=NV�\�L��%Aqpi�gV���'�n�"vK�����嵵��ű�z޿��4�W~�jjf�d�l��m��7�E|��0� m<<*l�h#�,�kkS������E��ݱ�P�nn������7�sQ�(��Z�ݥ�\�TV����Ѕ���((*���<j�a߲l�p3|
4�ň������=&��yyy_fY�9>����<<��9kSO�|i�%�����w�G�K_;��f�L)b���Z-������c"bq��e�Qܐ]�-�!����ֹ�L�α:�%k
�O�kg��K��XX@�O�\�=8hȚ7|�R�htՌ�H�)����w=}(�G�>�V�;A�����w����bꕦ�����K[A���s��!?ޤ��)Y-H�l/w)=F��B��k�����;=�cn����N@���
�̋_jkISk%�Y�ѹ���7Qi���:1���Η��T<?{E���U����٢��v����Dh� ��oݙ�+�T<�������BXbB<@#�LG�$
�|�yt��8��j?1�e|Z@��~����CK�Zh���t_jl���т���[5u=0 �����h�usVK˭1s�5g��x���c�����\�2�ՒH�������w������^��~���X�������TknPbecc�l#v�a��$��7���1�� A%����C<^���	X����\dGG��u=��M{��^�&_�yQ��y�e�`ޥ���qmZ_Ta��zp��2��{s���A=��Y����%���Ö�/NB󌽩�i�K�&�P�Y�3ƹ���4�C1�W�!2�ٚ�T�K-;��x�qq��x���Qw�4������hσT/��@�G�8rz#K���qo���o��A��8���{�v�LF�"�'����]Avtv�J���y����.��H���x���(٢�M%�[�F��E���$+5�΅��kK-h&��V|�����+�R_m�i�)Nω���(̉����>>�<0 ��ׁ��P�(_���rTn�9�J2�IDs1��'6A�N���iLqޫׯ����B��z֝���.��7@��݋���x-y<<�D�kg�Z�}UUb��	�k�����	8�V\H��OLgI5hb�L�Qw`�j���P0�6��c$��7[���Ν?��l�����-%6�8�I�a��	,'[��h���\����/r�ξY����^�SZ_���+�+�D�ٲ�$�K������3��:D���k���?���g{.M���z0&���rO_��$�A+�������)���h�1��0ڲ�G8�n�@����!CP�P( #��R�=��b���y\S9^�~�b�Y��߁&T'�|�G�,z�I�f��Y(��v-��������u��g�4�C���Z��r"��g� �W�V�N���Ъ:��gF�-�~�8��;����z���Jի�ݻv�͠�;���k��H�1��~�{
�p����h���[�-��tQ�w���R��?���vv��|�6Q,�ÿ�����D�7�:w�}��͸흢p�K 
��G�ݎc���4W�t�=���w�Q�P����
���X����ͯ��s8X��B��>�F�����jdC�eb�\]4�ąN��/��Y��`*�s���m�EqR�R��2��f�(4�U\���	P�����x��GQ�
E�m�]D�=��ڀؽ���'i�+��tޙ���ӌ�;��TKK}�����\��gJ��\ZhGy��mv��S�jyd Sd��C�~��!%������.V)��HJ��F�����<.H��z������7��s�^�*�G 9/D���lv<�.�龹�~w���=z���6���%=B����0ۅ��Ҏ��{@��j��慆Z�Ǯ����j�v
Vy׹�>'��5x�EZ�	k�����ޘ�{�T��9���K �G�L�՟RY�
�D4z*4X��xj�5(����7Co��Ih�JN�o��*�����_� ~�R=�e<,�,݃'v`�LB��9����,���-��M���qj ^�~�/������S����?y;J������=&�me�
+������s��k�4�j�f���=������T��t����??���.Pϼ��ԏsZ�b��=��T�՛pZ����*�>��j��܂H�FMo�/��I,j�B�D���"̓BִY���yd�ʛ!ĩ�9���C������cT����⧶8#&�r�P������ڰS�-Y\s�O5q����Ai��$���jn�0�bTl�����ϩ��v��+�nn��3z��/���r-�6ȸ���}�x����꡻�����nMMM�-k���U�<@D��|�r�2w�!lܜS-f;E'����y@���:�R���q��ϯzt�B	L�i&&��8Y��^�]�T'p��^�z��$t��J�=X[�s; ���H�����F'5��B��Ȳ���S�Uq��P�\N�Q٥�TǗ�[������>y�����~��,�������2�wr��/Ma�9_�[���|P�X8-B:lF��_[�ia)'�IVZ��v�nms���� �7��/���2�y@�VTTdV�����s��bU�M��]��c!nݔ �E��5I�^z�R�K�.b��TC"��R+ɺL_]�h�z�+m�w���3���������9 ��9�o�d��+��� �쐏�����D-����G�N�k�V�P��~� K�p��`��l^0ٞ���%i��l�Q���Q�Yyi���mMf��{yAA���w�R�4i��bg�����n��)��q�����-е}'�I�aJ���昹k]��\4B��-�x��ew��?o�w"B쮉	'H�'@m�y�&m�l����~\!�V�������=Y(;w7&��D`Y�T4֎�Dc����!}[Wr���,�>O����ɣs�S���(���ۦȦ>#��:Ew�~�y��g��jڼl"27r\�󗏿*�6.��p?�"��(�,�[�6�d=���P������h4pN��!�y�����-��,�L��`�6�_�֋f��r
��Y�*q��/���(wW4�����&�B�Ȳ0k��шL�ٿfK7�*oߦ���u���B������@�L�_�޽~:�z^l����P��59� ]F,<�C0Rzi��`,&���x"r(���L�A	�	T�5 A��f�#�M�+ܬX�v��x��y)�����X��y�yX6MJ�ib��6L�<���d��ރ�0	Z���b!;���6���ϻ5F^͟�A�GEG��U�n�	r����oR6�ƪ��LD�`>(���b��w���II�m�����鯘Ab@���s]x`�rb�^ʂ�|V~u�� L��z���V����x�Y�����V|\��NP�+sm��]00��J�E�R,AP�(�]�=4@b��&t֒Pj���8^�ؐ"K6n5��_%;��+�LA,������Ä�8A�6iF���R�K����5P�1@��3�o��݌ƙ�B)�ϐ��>Qo@�d�����{CY�+G=�[�GLAAa��حE��Rc��T}
]�VQ6 ���ߚ;�s-���y5;��{�/��E���Q��h�� $�p�f3�jk�����E����k� 9`p��:��$l@4d�is�2���X&>9w����徔1A���ǯ�#�8?�a`^K�2.�i���@ �6�p5�j�bNOM�|�9�7�P��Y��g��8�ݍꍐN/ᘻ�W�_RR��<AE�N8�l�1fn�oj�o)�c#��'���?g<}���dߠ%B�n�[���W��	�Ф�6i�,/�*w����U��/��6CEF�q�3j]\�Ҍ��ܪՕSf��`�нN�� �F�ޫl666�UC2Z��o�˛�<���ߺRµ��� tg��5��<'�I��Qq�#�`P*m����M[�X �� r�V� )�O������l�KuMM����+3=!@B�Q�S.�q�|��'R"(g�Q��i*��;��;l�K8��������g?EtТ|s-:a���K�*��xU��V�0�0���gǬ"`�и����a���ճ�E������)�,S��Iڭնxg*���?4���� �f���Sw��6�~V#Q����VM��,�vq�|t8����<%`a�X��G(�鬓��2�Ɋx��v}ح4�yt�XvO6S%�ӒJJ���[v�X����S1pC�@�K�9����୏VD#
���߾�������C�7Xl:x����9����1��/��28�u�Ctnۂ��P'[`k6�{S�hw!�h����l��YE�C��HލB�˅�3�TH�g^��cC���7���~�8�n��îJ�8�i�ޝ�$�Ey�R��,�@��y����&�����
:쪒�����qR"�^y�M&YN8����4�q͏C��]n![94�d���q5>����V����^�<B��2 ~���*��zWW�J��ZN�����p�� �����KKK�;��Vl׹a���s�YYYP�@&^�o��Ѻ�]����ޫ��=����4QWW!y�Z9��A��uS �#�R 1��o�����9����CIR�{`��f�4�l�6��R'��l�^v�Q�^E8�k���X�1Ԧ��=<,hx�ʽc���A�����P�jk�1��ڃ�A�<������{�1��*,���gs�������ttt�z�ѥ΢�9�������ſQf�[�n�黻>*@����@�����=9>�.�~��W���i7xh�흝L�*�4 �/6�Һ�0���ϗ/2�%fmEF�:��z�\��ϼ��}/n꧳�������T6�����;N 1����??h�6�.�2O-�Qy�ʃC�*F>O�|����º��K-�g�R��	9Gv|(R�2�!F�#�:��2{ՓrS��aS���I(p dr������Z�󎊊����d�kn�����72y�t!�$���1w�B���w�IF�l4�j/zӹ�����)u+h	��z�X����� �`m��/�+���g�.�R%�]�H�������ۺ���ve�i��jӏ���loKὸ���"z�L�"���A������|�H��.��1�}��Y �yݙ,2݁���4̂tvK���� A"4���%y%��v�}|4ʗb&���Qh�o7�����~ỤJ
K��A"7��#D�_ju��h*�>kʤ��[� ���ci����ԤRM/���ա��Lȕ������s 9�a� ��6���f�Loۼ�*?�Dg	�c*�I���I�_3�6�Ղ�������s��m��h6=w���u ���܇V�a���X͝x>���B����@���ܢ�����B�5�2􈑜�:�y�?�43y�/�\��<����!	d��ϫ�Nc?PXĊR���)� �O������T�׳��ӌ���+���\RbƄk�"�"(˟��K��E����eQ��I�
i�?tq�C)B�;���uo����d�O�2���LSts��ؙ*Q�E��W�?��Tf;�W: ��q��Xl}=+={$˃*;Fȝ�*S"��x��.������XkH�픗�w&�J ��x���g���f)��a$�wG��>��A��^�}�|��"#��z>�LW%���$.H���S�cFӤ����]�1�on�p�9*ZJ��6�/7:��}��HO��Q�^o����R�l�[���v)��g��6d�0vO��F�[}y�;�F��C��A�s"�l����K�v�f���{v���h���K���v�C����\�}��F�bI���f%�:�{{�
�L%Ʊ>�{�C�}|R޽{�.�E�ͬ�=�Ī��Ē��e���u-��1��nX�Q��]�h�}�؛Y��|[v!����Q�ˊ���g��:�#jN.Z����ᣒi������^�����9(ం���\��4:'�0���,�~�{��@�m'GV����׹s���?d*���q)>�2
!	�e���ܳ���A��;��Ж[���!K���᥈B=���ez~�z2~.%�y���X�������	=	~g���k'�r(y��VLH����ݠg�����d�O <�Y~J�n��W(��h���v��=�ⶎ�+�p"C`+�G�vy�k

�dn>>�Ý?~�}��5M�[�|��ș���Xrh��$�-��6H�0�4��s||��]Ĝ�_6�|?�D��5G�DV�%��&}�S�D����ZtDY�*�ߤ�x��g�T��SXk�DL�6���9p���v6�������4�$��,�-�]���E,C�(��c�J��u9Taߓ�'H*o[$��P�f�`f�{�@�B�T��NT�j��:oN7Bk0�N�	=����S�ר��[�� �X.�.�:��r�f)K����G���p����ǖ�s���|�k-�ئ���P�_�ʀ	�
?�T�}��%���Gm#��^W4�j�e� u��=��5h��h.5].�条�df��������!@���RC�$�Chjv�
�o�>��P�n��s+��3D������²��Q��!y�2��sՙ�H�TYp��LΌ�g+e���;�+#�i䨕8=I~pBz�1���Y�}��tû���G��$��z���I{zv�:��&zE��h��$���-Ռ���x5��	����
���QQЉ&ҝ�x���W=0���nԝ�ݪ����,��Ʋ<��i�#��B�����[|^ԃ�����<ЈGi:P� ��q���{�$oܨ"��l��9������(^�nrO3�hyKRA��tc��W�w*�R"��@B�EY6�Ю�N��,n��H������A�/���(�r	if�r�P�X����Zw��6�p`�j�*#	a�S�3��N�ц��X/	��?d�CʒC�no�/G-/�"��"���Z�z�$q��+��~=yv+Q�&�=�9 -��s�C����wC��0��c?�Y1��Ձh�����i�c>^Պ\#�Ta3����"3��v|oCd,+�@D�����Tn^����n����Cw�CS���Uk?Gߴ������EN�@Z�ﹲ�(�z��:u:�� �NA�js�q�F�@ΐ����Y�E����8��0����y�UiJ&III}¢���իW�!䝯�}���m�#?�$�oA��	�F��z�̴���z��(����������&���N�s����M�5j^Ck�>��]�M��;���E�~}~��m�Yh?�#�7�%�;qU����g�է!h<d���N7��u��p��,�*mCł���	E�]���'j��{7胸0p�j��8�iEI��w�E�K��Y�7v	f%)��֟a�7o� �g��"�|��Y��7^�<./_h�%����L#p�_�Y�g0�lfG��l׌+�G�{�	"��u����q�-Є6�sr|�ZX�Ub[8*{,�~Be�� 
*֞�+x�N<�xL��Jx�@�����?ڭ�qZp{�D�籋�C���/\�����NY�掣�K��x���zү�X��Ú�u���%)y��[>?j,Y+|NԮ1c�.;��������j���y �9&|~���:wkѯ_�����z�0;�Uyu��4C����٥h&�9`��xAe4�m��/?�Z�C�����tm�]�J��i�mt��{�3� �o��h9׶�Z�9��H֪��l��s��#��"Q��B3w��2Y�xH����0J�K1�����׼�ѫ�F� e��1e�����W�����.RO���G���؞SRQ�k#M ���|�s|�s��p���jzSJ���0��T�����2��ow��H���?�(�1�.p>����KX�J�!�r��D��ۑ�r�?-�l�0K1�o�*t�[��|����&_����Fq�/.��k��g�U��Z�M�������H�r������A�m�=��� �x��$+�]�
�v���XQ$�
�xLSN2Of�b�|)g�����{���ljt�������d�YI�#[%`]�:��S�F��~��p��y=9��#�n��Wh~2��
$ag����hĭv&@^�"��g����b�&bd�͖q;2����0Y���%=H�v����|�G
�a��|W+���r�>�)3.s���{��_���>f����Ĺ�K����˨L5n�*X!�Sr���y���\�7����!���ͨ5�5��}��z|<ʍ��Â��E/٠��V�%����8��"�$$��{���x;8|�8�ݕ���-Z��c?�����V���K����e��\�����bh�X�b':n��{���@�C���=O�|�G[b�0�LM[�͉�u�"��缊>\��9�q��s�1��ZI������֤4\"
G��g����,�����&1-Qu��@���;�'MTy�g㗻��:�����/�k��qo� �p~�,��N�ҕ0�G�s��q����ˣa ����
�c���}���٦6��p��Ԫ춪�]k4b�"������sR+�0��c7�������}rX:��p�.ۓ�T�w����+����ml�3�CyRW��wZ{d�E���z�����RUUU7����N������j�5��ku��u����	���)|eR;�6��f�s�˅eS6���f�����
D��+`�+2�l6��-4�J˟
��fc���H�¿�i&��߳!�db���+�=Ey#����Ua`clO>O�.�)��M4+�X�*����`v�����E*�.;�����;�ئ^(���l��������5�pE����)I��pU�;n������lpne��%*�sxW�u|`�D��xh}0J��Q?~�y4"�a�m��<��e=��j31��?j��U���_�6�0C �o���~:������-�>Xai�h?� ���*�j���b:/ܻ����~]~AA���������08��Ԛ�w�ט7�1�|��ND���	���o��s��m9?h�ݔ]8��d��F�Q��4l��ND��~V�~���x+�8�>/����
�Y]	��V�֍x���Ǚ�~��,g䊗��8sN�r��F�����$:Cs��n���N�G��S�����r羱	��H�WWW�=�	����)�f�k	���Lr^Ц%U_1�F'���s[q5��P���|�O�һ[�xP�a�C��Bȵ0_#��Ȍ$^qm��S����o?�p2 ۮ^�[};�կa2m<��y�hi:�x%[��2RX+�}�`�`������e�a��/#V�be�Gk�^�	</�]����Y9�ؾ��{��;���DWc��B��E�C?��R�L	&�h��H��t='���РsE�PHP���4�`��8f����7��������[g�};��.����Lك��C�4�E�x��Q']D��^���lN7f)b@6s�Z�@��܎�/.kJi$x[�/&GR�@$����߭�#<�%ݭi�t�E�R��@��@�dĊґ�;/Q�S�����!L~�c�l�8N�z9� :"�R�-�W���I�ȷ�("��[��BBq6�A�@G���j~����~Z���-E�]��79�o��_��c
�t,
��fV�8�>�4���9��o"?�:Z5�l�������{\��?�"c��Z�I��6�ZS���R�ڃ��5�!-��O��;��T�Q�f��P��M���ڳ�拶��^P7�$H#����z�_�X�6�!c�ea"�H��A�w2QW��G )G3l݇(	�Z�X	��|��V��=��d��q��XP���gk���r�΄(�Z��?b4*�_��$�֮��U����I��-�8�#���:��N��u�=��}\4F ׬�Ѽ� ���П|���g$������/�:Uc��%���-���e�v���5Z�lJk�X'8r����^��Z;!�����N����l���42���1AQ-4�ט�\���O����d�h,����+��D��\'�#�����n���(�Rcx0l~b�1�6:׻x�0�Z&p�t�>-I����{���:^�Ȱ��JD9��5]�D�Xo���ײ��Ƽ�:b5����I��{�ܦy	��T�����������V<ؼ��$���3��rW;��ɔ��̥���R���5w�4�hDz�gGCI|�m'��[[{�b�+��22�q��?����n�O>>�Q��3��G�;5$�z�ދ:��WyZ��8�lA{�M���ɏy�w�����-]/� 'h�/�[�o^����4F$ �^Gn��`�u#�ZkS���_��Ϩ=�Qjڞ��mGVh�f�]6?�kI�N5����l�E�M�����=ڏD~%G�H��3*�ݺӤ�"�I`��'k�����GݾM[kC$�]����??�#�����ǚ%�rR}��)2���i��۫'0�r���q�ޟv���#{<������C��FC�돣�d�;��|��7P���oV�X�f�A��#Y�ץ�rD�-L�?y�PT���7F����7���R��/�x*R՜[��O�0��g9HY������*������"�9)����T����כ���BI��ͨǄ���F�'vɿ���04�m���:h#F�d��"�O)$`b�MI1��*�/L�0l]�������w=����]��*R�A����e;����Va*�@�`n�!\��%S�l o���0~�'�\ �v�n���	M6��t�U1}�қ�7OR3�S�4�v3��?a�c�y;{~�B��j{�Wn��ã��s�{H�u���PAm�_���ٽ����8�Yrd�ng��ApwJ~���fsZidܲy�)��\�E�a��dl0�4R�tE,�4ƚ�0�x�E>�>��wK*)5�-���K1w}���EҚV�k���LK~rzo��,f�[��9�Vd�ћ�☆\��G;�?$Pj���hT����R�c�z�D��a�u|����M u��=�]����?�0 $U�h��N���~�%�[KU'���L^Q��% ����+�ϯ+`��pho֚��_��fG#L�luv�sc-P�+H�Σ���g��ϫ��	
�#��4aUKWD"O��ޛ<m��3�U��	��Af���2P���Ғ��E�~��Z ����hī�xω����=/3��6X�WO_ެ�� ��Q�8�e/�F�D8�=��c�J��N��TOꆞ''(�D}��R��"��r� ��w儜�F��Z���mRC��/��t�2��T@�`��˻e�9��@N^��K�.z:�V�Fj>�6w>5x8�S�k�Ba�t��G�2FD#��Za�>�L����s-qF�sa�?H�%K�wM�6�Y������	���.-t��>=�iR�C,f��wc���wt�UO��9M�t)LR̓m3����+l/S	�<6�s��)>������{�\���Aq�_�7EAS;ܱ���WL$ztC�?���ID�+��!�+�bHV��N!�LdIp��Ǭ1j T���#ԯ���6����_.g4[��4}#i�v�ߞ=�&%+t�Aώ�I	�2N����'�[����R+���;���h�X��;�[^5���Z	�M�mMM��P�Z������� ��9 ����������Q%���|}�ǀ�c?i����lNg:�ɳ*�~��0bc��lVE�l��l �B�[�'H+_5�'�.��B�����[7�kEH����K�}�t����؝��Ȥ Qc`~�7�E?��IYy�� �ֻ�5ZaCK�t��i�`�gv�N}kkk]Ss�N���{�Zu��N�*+^5f�Msh�g�|8����M�2��_=e!�;���ɸlv�7��_��v��M�(|�6k�X�2����n/*� #���eT:k�"�wp�p�'VM�6����0�J���۵�]%2/�&�^�:E6��E��T�#�]F�{�1fi�@:����>�vU9������jqϲZ�/���<������h�qq����n��%rM�j�۪ ������88-S���C�D��j���T@��sJ�7�O���,0҇��!����zP���rр�٤{��l�ھ�T;�T�!:��/�<J��&��i��-T�r*?~�W;RoN�Z۞^`�4fd�[�N#����1H��/�g�qթ�9Ȥ� �L�&ZP�\������#����5�:�o.�&��4�$�ioQT�X��B�¤��~=\2cgO.�*^�X��I!����S������+��ܹ�y� �ޟ/4b�n(�$š�?рiL#�ؤ���RG� pQ�8���ı/"��KG76���"l �	z�g��Эq�UV��?dX3�%��
>�>�,_c�)�}�
t����D�4)2��7zN��X���?�N&��s.!�����'���
bx'oH��6,��N��G8�(�&)��q�)~4r���qO:j�PB�i�&�L_���?���. ��d5+���t�Z���o�Qٵ�����/;��ݴoo�GG7,I��L@K�S)�֫���r�>�����������V7�\�[1R�c�z�A<mS�k��~��א8��,�,P-�7p�T|Ƕ5W]k)������PΣ�ū���\)��`��Q��=(�cNZR���p����p��! ���~L2��/��M�������Z����QjUgV�@��ٟ��"q�U�U�^�ۮ�m����B�f���|��=�-����	�M}	�.x1�{O9��L����y>ZB�R��Ô��F'�B{�
Z�v�NP�s�t������_���.ȩ�� P��#>���_�]����>��ʿ�q����/Oy@��x�4��="��_	BK5p��v#��,���h��4������=�F��S�Aۿ�p�*,�������'��p��#�H%AowS>�r5B��L������z�W����gg�e 
��s{���r��Kk�����HV՞K:>�Iz\�������wYY�c.��G�������]��)&���T�9N8!��/R?�H��17tK�+�1�5�.�Oc�E�Yr-�',��Ts�����C`���nl��C�~]Sk&p��c?�Z:Dp���U!��ۇ�8H9��x�c����%i7F��d�<�ڹ�Y|�0迎D7hu���,},�@�_����%�!l(A,zz�(Tm�b ��5@��Y2�bx��4�"fMi����)�,B������`�|��ޞ���(��� z�8m�F�{̭��vOi;z�����Z�.:�z!��R#����o�������JO�s-�n0�Թ�C��}�y��9!�g8�+������dwVmuꯜ�q��jsq�qs����X2�{8@�5z��Ub8.J�!1W�B��"z=-R"+}�]Г�V���q��A QVv��ڪM�@
VH6��,*�KO�8䴳(�^
��XU�r`}4��ϫK�__��Ъ�ӿJ�:���^�p���:�
�?g.
�}��þ�~�)�_�	�V�QٰcG V�*� ���T�2�F$,�>H�h�Ӏ`v W�]��l�]�
��m@r��m��hzJm��#\�����S<g��/z��[��H������ɺ�LE_J����|�g��ƌ�A7�ھ��V�g�Nו��� �ˬ�t�WЦm�3l&�)]�h���t�3�D+}���%�gM�f�]q���j?�~�ދȣ�cX��8��w�n�PfPt�|��%�sy�:�N	����"ܻ�L�S�#pԜ��އ5�,�O�O� FH����T�[��
����	P��I����$��T���x@嚕����ӧ���z�'�Z�&��~�z0a��t@�9[�%G��Q���r���b!��D�-[Q`���'4~ld�S}_��L`��<�����[��a�W�Ŧ��Οģ/ځNh��Z�p(X|1��8s�Zx �-�A�x�ʝ1o�t�ʿ[��\C�ҩ�\� r�K�hPuu�������eĩFDB��R	N����,� �\�}O@���������"�F����O��.E3��pG��)��s��Ȅ��P��Or�\�3ۀ�g	d�[�Ag���U�hE�����R|I>�~ŵ	�߸��ٲ��7n�5���fd��X���O���D{���5\�G �klBp��Mv ���r��? ��C��(�J����)d����BP)�U�y�C 7F(�����g(ݨBN��=�ѹK{�5�7S�g6�_7��~�rp�J�f� ATj��
%7,IK����Veh�r�a��<�p����d{�d{���/�M��c��m�~ ; tE�tp�돣N[�p�u���a,ep��	��t~Z|������I1�s��������\d,�N�HZ��W6묆d&r�HhѤX�|T�/��vPk'lS�?���	l�K�"�X$P�c�%RtM�&��c�W�8�ٔA��$Z�Y%����4��	[^�]L����Ԇ��џ�vw_sQ�����y'{���^�.fp�Ŕ�"6�}�liX���j���v�+����8H]͂Y��>����ĢTiJ��	���g)6)}�B+�߿ �04-^ı,BO#I�PPP��ugUh����r�t�y�/-���h���l�ٸ������3�3ᵅ�a�d۷��h�;:�2Z}��aq<sXq��귌�?��Je�`���M�vI�B%�M./;L�mM��7`3������5~������f�͚0�g="��4ʧ\Dr[��Y�[��O�ݹ�˴�P;����_��>��RO�ٔ�bX�� �*�=��p��p|��'�k�'P���̾{ �6����ݻw�0��U�[;��{�㘋~وA܆����m���ǽl.cT�c�@��.ES��9wk��g�2K�d���J��Q�z��!,jR�_GA��;��;UJ
 
��ƈR.]��?�g��/S���A��C�#Nd�Olx v���a�h$�����_�H«(*���Ř�K���D�-L��{�b�[>D�ӝN��a=��F"���^&$���C,0�կ�����[���/��V5��T_o�����FĿ�8�� &�@��bPw[�������i��eh�A�4�N���T������}[�tS��Ѩ��x�Ъ�e!�<rؒ����E��'3����ǧ<�%�/>�p��]iz��7M�1~v{r΢���И��Ŕ\�����lU�����B#9fn���s+������tz?(���p��`�3�n^�]�Oүç��=L��?�خ!(`�=\j�I����A��)�ޚA !�X�eZȾt��1aͰb�S�ܠ�3�zI(�ԓ�仢���:5h���J�$�(H9G����HX�g�434�A�,lk�*�5|?�"��<ʬQP�y{���$��45���3Yvf X2����Z]B>��~l}��p�	J��-Κ�'P@
B$�rn�y���Y��~[;�����~���y�̃׬��rJ"gb��D�9+����KY�_(��V��ڔ�.R].�.�Z!8���ݘ��`C�S�z)���>��ٽ�%?��jn8AD���״���-]�ZX���~. *m�NS*��,za�O.��&h���W ̣������R˚�L�u��oA�Nc�� �K�M�/�O����64yL���n�.[�D2ڬ�͈���S�j� ��y<w���)��}�.������=҄$D�Rd�ԉ"߼L6����c���|!��\�費A�4�rڎ-�Ct,�ct�y �k���R!cT�|��蟶��E���XR$��@R
�#έw�.���E\#���4gbv*.z�Rc�T7홏��I�د#nt�����?h�=�,b3NN�l����c	6�׼M>������Q�	.���SK��x	�a<B�E.�Z�]s�Z���߈��� 1��֐�D�=S������T����V2Zf����H[���ZE��\�"ԕ�F\{��}�E�-���е�_o�����N������|�����B�T�����Z��KS���<�?�3���%K�V�A���+z�Ϥ�q.Q��':��?�ُ�=�׿��84>ZA�.&�
��Lw�!\=�3�=��'Xc�$AЙ�%����1�ָ����^���7.w�d���C�),��I.qʐ����{߯�c ��p��ҝ dj|�a�� ��B����Ʒ#��~��}gy�oqg7�C�ڌa�m͡�ÁB^y����dv�;��i4�5��]�\~!��Q����<p]žEc��>���P���c৞���4�8��̸�-����L2����f�;t+󉦔��F��l�dK����,�ݡ�c�pg�E�iR���#T�/��ۑ���fQ�)�߈g�����^6�3����!�bE~�&��ş��X�ؼOkג?�����73>�����
Z���u��{�旆!�������oP�ܦ�j��0���|)l��S'`S�P��?�S_s�p��J���9����d[�T��,�Y�Е�{�QW����<�G\��,4�i8l�A��͢��Tm4�C��3�P�$���g�CE28}��З}�tZ,�L_%�~�Qټ��]�F�cv"T_�:
5�օ٬0j��S��m( ���1���61���2�)�৮@>|�	X�[51��;XSwy�QG��\a�u�?ſà���Gg��& �f�Z�% �Sg	�`B������9Ȇ�Ш�X���7��x�d�	�n���!��o&�P.��.�ڮ���e��
��K���G�	�~V��}2*c�UC|Z��Y�����B��$��F�5 ����7x�jEct��݀�l�U$]��{���"]5�~���B]#4��acN:V��OZ֊L���ts�Fi����5���	z8�N���4��2RLD����1�u��~�����{��f���,;w������Y.��aX���bE��������F+��n]�/5�����>y�[G�z�J��f�!6/|5iv���h��Ȇhሃ�;4�#�}�������������Fb��%;��DI9��,��ڧ��v��]�,�z�)s�97 2����DLQ�dKl�U��9!HoI��ܓ��J�.����E��ܜ�[���T��{�E9�c�����W��k&�/�CշEA���=�%W����_.I�s%��~�7 \�:x\�|d�U���W����c�ey����'K�._����B���/b�����E�^O�F���"ԗ�"�� ������>��h��
]. ��ؕX�H�9�E~)z�ցb��0��&�LŹ����_2����\y*������W��������JQ��dpvr��S$�,I!���r��띾�h�&`D���&�;�i�J3����F2jcû;��Žėc	�>g�c�ZZ9��O�Ζ���5Ł(���T�|����`B�`*9�D��7
h�������1�/I�e��4(�$b2�6�k�]���:�y��@wN���B�f�ϒ�>�(a���>W�=��x����R�A�{8�3�����/�C~�4:
�8�^ӈ���}��:c3����>�"�-��ZhKЉ8+r=fj3b C3}�_����b��c�ae�Q'w�2�BefJGcP�c�m��Pz�q.t��`�%׼c_;��?�]���q���{"�wHE3�VO~(�|3�~�j����.���g�x�*��*,G7���3��q	/�Z�:� �uh9fA�Yb����@*S>F���>:<�i�X�I�-���W�����/��>׸Ys�S��7�7Ug@����h�SrJ���袅����!���>�&��M(�7>����l�^�H3z��sj��g������;��,4_p�DW'g��;Vfl�t��|_[.%�m?/d�?���8J7Tor=8@:�2(~�(�R�W� u(	���W	�Ǯ����`n\<p��B�
�-��~[㪙��s�`���]o��$7��O�v�G�<;h0��^���S�_)1���>�u����&�+��e,�R4�:�Eȓ��W
��O��$���̠,D$x|3~�~+�/ ���ac��$R.�:�
p�7�ǲn*�:�����i4Zjb��k��rJ�:�>o��R�U��hdl"�P� h= 5�k_�f��A�6TJ��	��R:4�s��ZvO���M����K��5��O��3`�X�y�y��	��I9"^�E�Կ��x�g��@,(L:��,*�n��s�$���O��$ʓ/��
���2O���=S=�BmBr�a�!Q�?�n	�٨h���������<(�x�~G��0)a���bXu1��p���"g���R '��������E#����=���**aE��O�����~6ό���׀�u&�=�и�<`�գ1����_;�)Bc�}���Э�~W�)I�O�a�,5*�*,1�1��a���_��'�I!N�Ms�f���ޙO�;v�-�p�?SL � t���U��H����\�e'O��%�H�E7��#E��H#�+�>��ܿ�cH�j4��cȴ1(�
�°�t�)z��;P@5=�H�?0y�$b>�)&�S 29��`t��`K�T�bqhss�}���F����|{N��p��r��L����L��f�:;��sB���u�����,�E����+���z,5Z�m�Q7��\��}�e�B&�0'���p��-N&�(�l����?&��āl<Q���5��c����i��w*��iSrf�wMxI��UN���W>�s��� .�"
O�d8w��er+����rJ�R)�����1¶I>�D�8�<X���:�_5IIո@����1sS|I;6�RDq�: )�,�3m�p9'x14�#���ƑOY'��!�9t�5z��5"F�!�����;����c�9M�wt�����8F��;Y6~����J9� �BY7t�+����lY�m^8�p�,��E��X�d����x�u[4�7�8�
h���"���� �{��w,,�;���r#�S61$*c��IP�

��И��q%��Q�$���`__��X��a
�M�ad&$��ᑃUd4�c��9��A���{I�;�����ѐ��$+��@������v�.����&?đ0�@�e= kj_m�����xX"t��$���bݑ^�"��������@�+%�Z�/�?mѨ�֝�&;u⡦�͔�{�=9CE ��
�Ñ�K�@�@ɻn��X��R�t4��L�zG`�ba��D�S��w!���^vݤcoBW�(3tX������Rʬ���Î�^���JGޞ<Q��s��e�9��$1I���PRTU�{d�����7�[�˷�y?Փ�|�I�XF�޹j\m!H1x_8R����&��N4��U�"`�>%�Et4X&��G����{�w[���}z�
k{]�[�{�0^/��u�[-L~B�:1�;m�\�IkO��^��@s�"�p=�*@u��'��M�˙F���C��d\�]L7	qp�}|�{��1/��'�G�CtF�ߪ�L-w�}���l��%���^J^�ey��z,N\\��|N�i�WT��Β;����B�T�e���k
���!"�P	r��vbV�yu�_�]h�%��K�m�f�����Lx\xZZR}m63`|�J-9�r�N����l�{^�9:��U����i©�'�<�c��"i�<�,`�oѦ��ﲗ�y���Nw�Hɾ�9:��}ΊH��p�H6&��54ۦ�_9"����+����t�l�x�ĭ9pp�J{�}�p^�{���J_2������/P÷�
������ ���5�!s�:!��l��'�L6s8�*=bʬh(��ur)��$O/�H[z���C�>X+�Q��gX?�E�z�^櫳���`:�38�(�r ���T4����?�P4���3a�!�K�e_��m��2ƅ\Q`{����wq#�o�������T���w���WS��(�h�QqoT�@K(1J ��&Fp���`8I[�I;i�8
L�K��~ʀj��ݻ�\WJ|�V�/����}����K� �"oh�SH����_%�Ţ�B�v����w��7��c��6�ׯ�c�F��۝"01�b���"���B���Ξ������.txoj\3��ãz�O�hB���qYG���{��(��d__�$�����ih�F�l60���U�8׸�F�!/N�PM�����G����@�o�2�<	=ᾙt�6|�8G��z8�v5&���(�ިq�⥠���N߹�&�&J����:;!����Q[7�)���(��y��

&������A��]�3@W�Og0����
���J�-$v�B3~b�2b�|��i�N����,j��ǩ�����w��0����&��L^$;��
ੑr��D���dQ�S�+ާzUu��S^�?��]�@?�Ky��*���4H�L�8�	f8[jp�B�/~������.>���b����|"���q�.�5{������^�'��	���m`��jz=���-�x�*z���۟gd?q,��#�X��(|$�p0U?��-�g���E{����er1h�?%*�H�?B�-�GS����]Q�/_�GU܆nA*����;W���Ls���!$���C9ڱ_������"O�U�H�& �?�=�_
���\�zd�A�)��㗝	��7Oz�:��׍��3�vjJ�w�z���ئ?F��kl504�e��{�W�sK%AӉ�F�ŝ��w���ûζ.�����D6[�!C)�^�1"S���L�#�`���hm�荛�Z
1bv38��B��>n�}�(q�TQaoc�+t'<��ߣy������/����:텒�Tg)h޽�p�� w�=�K��7ۗk8e�@J�"�$,�&���=�u�{�tc�7fzG?���ֱ��j٠�w���j{�Y�kO����%8*w����<GR�n��hc�n���T�/�W�^U�A�h·3�*T �TK����W?��J5���D��� _�E�{�'8v����	��&���dI9:'��As���^���(�Sm��]q	H�#�]����!�
��_���ip�B���ÝUA�v��,��~$��aa������9����_8����/ۧ�������_?�o:�|���ၽ��2?8�C����	�}x�i:[��y���0;�$��'���GSߥ�Ε�����/�w����<C)�g�*Vy�����c�gy��ˢ��dgUSc9� dB�2�۫��R�ˀ?��(E����m�V�st�uZڝ�P4������_X�N��(z�MY�sM� ]�,����$���$�����:{;�UC؞�s��e�Q)$��.�8K�7
��=47Ϡ�憊t��|��E�=?�����KZ*�=	�ޠ�s�:��l1���R����bj��T�>��C����ZJ!����]o���(��"�_�|B�ك�����G!�+f@T9�l����A��� C"��N@���9x� ����l,�����J�0��������$������w������H�{l�,�e%�L꽯8LR__ߨʈ�̚\a`9�Z���c<DBkk~����=Ѓ��s�%�=��=��M�U$�W��/�^���-��2�v��u�)�)��?�Ru^"�Ǭ'��#[�:;M]�Z��kh��������7������Z9��ٗ�De����N�'x�*��^�~a�����f~|V�+��řw]������Sg�ST�vZͬA�&әq�*�%��T�vxx�a�֏~���D���v�S�`�ꂆ=��6���_?�����W����H�h�Ba�����!���4{"ۊ�i�4~J��+en2��Ěf͋>�S3�� �j����iF�	�hP�H��-j�oZ2���1\#���N�M��l�]X���$̘���u��7����&o��]��n�^f\(~q��֘?�����ؚ��������)�UiQJ2Qq{O�0'C_�X�NO8j��1����A!
O0��A[Z�\Z͔`V�>Kj�/��(�E��bȖ����MD�S���K�Ey���b���VE~v1q���歳`�*w�oZ��Y��߼m�Pv�P"_�x�n/j�=N+�5����ϟ༸q�Gc��pt�z^�lR�,:99i����tdk'l?AA���Q{��wТ� �F�.��>t��^Ԅ0#��h�I�`���r��7F2���G����[MM\����#Y�d���|p�4t:�5P[8%�'�P&U�vC[�B�N�)&o|��&&&B�@��GB�<��Y��;�iM'$��,bo���MXCa�t�!X���0
WuA��s|L�G��Ci���^8v���Q����4���5�i�`/2���	<��SE;t�C��D�@����4�U=l��z��Аe!)Ŕ�"C���P��@��s~]M8Z��qw���o$���0a��go�׏#�s~��N$��"N�b�uH�x��CӦ�/�F�j�У-EEE���<�U��ΉY�R��;��c�����
߉���_OXoŻ��(~j��5#x���;CΜ��;¢P�9ă�2����_P��X]]���}�뇡V�o���D܍ T��|�����ih��0-��
�6ι@7��5�!Q�#5�~x���w�l��y�꟏����ە����(__��������j�%q�y,4��nTO(Yh��o���/�㷭���f��{�>ڛ*}��l^↝�h1�|���O�K_��]#))R�Ss�����}7O��,�j�/[/6p�P1;w�s�1⛶Q;��lS6޵0�?�}o`p�>�F�����N��88^>�-�[Oh��+)�k,��MD�ׇ�I�S
`�,�T��nJ��+��|yMM��DJ��j����� J������ǀ��� �O7Wr��!�8�69C�?ws��~�����&�Uό����3�/�Mĕ �i2�m�p�z��2�3�A�J�F
+�B��D)�ǿgS�e!���$�L���Ϧ�{���R�d�7p�Q��LM1M�]�:���k��#����[�܉��V��K/(�ry��`V�F�l����ki�Έ� և�D�zf��!��GM���}�!��'/��K�<�˚�A=�q�i��ё�H�:���h�14�7?m�,2/�_Z"W8���X4Λ��Ѥ�ݺ,�;�u���$��=U�L���N����7�I���V���o��af�,*H��m��q�\��ntM)c��#˕�L���w�gk�J9"�p���g�m���$Hީ�y6�  e��W^_��ӆ���*R/o�7���LS�J队���T��_�A���*�|�>e��yۗ�cT�X�
�f�o]�N��N>V֮��˗G��Iզр������(u�2*i�w�|
�R��s���P2
�f���̑Y�8��KY֛�
;}ӫ���_u%r�H#v7�-|��1���V�1��T���3�&S����-��~����[4o�zz�n�rwwO�����ո0�Omqx����~�Z;��:�Ȃϻ�ƅ�;�����I���[���5�1�R{<�9���~¬�0,<q�{� ���jd��W"F��t�2�z���^���7�*AF�k��zt赙	5I�� 
�M��'-,|h���,B�\iԱ��nuR#�͂Ỵ�-�#��8
Mu�'?�:kk?Yr���P>;�I��U��� ���a��Io>G�ڙW�5��՜�6� �N�k�h,��W�m������	xإ�2���7%��D�+a�"Qd/�;�x�3��O�c�7�O�GAՐWP��"���ق_�/�^�)�g^��!�OL4ϯ�Ȟ8��%ti�"�t�c�f��&mn�Es{�b� bK<S=� IG��jהOm֗�KZS�20���<{�:�h��(R�~��1�N.f<u=��b���)�W���_mFpݩk{��B���ua�~Gm?��n��K�t��A�I�������림j��&8�"8R�;�[�n_�L*ICS�%��~?<|������0���6���R:���qN�Hd��`�� �}�y�Gt7������D,5Y�8(�2�_[�B�W3�8���}8��|��#h�Y g����`d:KA���p��N˦��0�ε�~�6��jm1ֲ)�[k.�%Ś!�fJ��3c���tC�FFF��m� ���B�N��Rf?rd��TG����)�����M�D�H�.�s����A�qXx�Z"��ن��Q�w�ɐ~4�`�G�n�ӑ��1�~�<��Z9�|��37B���b@(;�Y��x��;������mL&��k]U��\�媦�F��s�20�����g-N�x����6�;�p��`���D���D�n������L�h6[7�Ά3�l��q>8�g�c*��J��ۚw�$>)���?������}�"�h�O��0�ą�
��N�cy�L�ΕH�� ���?@+K�|c�|�2<A���Z�G�тn�ZKu|�ds��E$�U�a��8]C+�2���p�����5���������E�sqX���7��!5��g%�{>|�.���#<��A��*-vzEO%~n|��w��i%��&���T�:�'_�A#5
Ŷ�{�����m�[.���������{�y A;�׃4�V��`�0�C�m-u��z1&rf*v�|k4?�zGcp��]����@�4��zg�\�������6�{DN�v,I�^Ki�aV�G�Ld������S^�� 5Qvt�o���+4%}=f�K�g�������7�൪p{v�%�瞱Ǭq�8�&���\o�UR����~���QƗe�[f�����RQJۺ	��S�a�JŏVIۯo4�$�)[vg����6?�Z�s�y�޿}L�!k:����o,]Vg�����<���q��ӬϰDlm~�m�J�Xm)��Q"���+w��9x�Q2��xskk/�壍huv�t0X��R�[
�>����-�a7�Q��ϴ#�h�� �k|�M�WSS�WǽX���'%���_&�.^��+���kk���>���g�d�~�鹸�FKٔ{�8�[�L��l{���47����5�yB���V�ꟗ���D�;�$t���/n7�+����9xvѩl��(�����2+��%L�џ�J�K�A�*�ڤ�_��6���=����[O�b�&��ws�m���"��M�� ��#��n	�d�:2~fN]�фh	��P���p!����j\B)���!��B���9]������O�ɚ-o����_go�Ā�	H�J�P�>I�/�q4�Q���!����Ё���ul�FU)jس��q~#�[��]�'���<mV|a��/����eW4z5���(�n٧V��T��ߴ��^�i�/�^�EG]��G���޹N�~�b�K���M�5��n�o ��7�_Mp�E$�6�c!ͅ][�n���JW��^�P�B.@9���e\� �A�6��Z�K�x���b�MsGqx�:���k����ƒ��h��
n_��`���qr�PwL�m��R�Cy
�tJS�"�ym7?r{d�t�ٻ.-@�:�����������,�7B���$��9�u����X�X�Jyn,�ߚ�1|������5#N������5KLϥ�e'�mb�t��^��Sm�۰�[���[���]�����U/�BSc<*߄��T����om�s��\dd��D�����R��=m��#�q�Z�����n+�����e�L�_�Q����dk�b��+�-����H��X�ۙ2�����ȭ�yU%����t��Qz��*��],� ?ou���^���Bn]��1h9��T��D����I׆��wC�Dlv������s��sن/J��0�fz�I�=��Ԫ��G���(TH1��)Zh#kt�R�`�4� qxtѩ���#��2��=�E<���s� `tE�>	���fӞ�y��'�΄\z�&��Z~t�+�ўX�|Q�/��l��D_Vh��X�S�i<;��l���l]��97?P���r:�C�_j@�Ve��ȅ��o��ثu���R�ᯚ6~�6=�җޫT�U��af8�����~_!.n� ѤN�S���w�8�y�m=� �rۮ�YS��:W� ��-��F�$��D�]��7N"n������`��M,�Y6Wۻ�Ԣ���sEI3����oztˆ��ԕ@����g��6��h�>�n\BiZ@}|���
����vvBs��w�#�`B�v� 4-���7%Ƣ`�����{,��V�{��rW��}2<@$o����:Ԁ�����"X���z���\�CYF�+TI:�Դ��O�����G�M�2��u8�v�|j�H��!���?�d��}�O0Fl����=:�G�}�C�){���ѐa�,MJ�Q����2�v��P=����R�����ϗ"}�L������!4��`oME�S�a�[��y*��G긮}.Fh���^桇��&���W�աz:;���K|9���#��1�k����Ҥl�>K���=����j'n���|q�/�bX�ܛ�l�QQ�۷/������tR����1�+��ܪ"��r󡎀��|�����*��٧��	�I�k=�V:��!���]p�kN a��$<�-:��r��#R(e-�gI�
�AIiiO��qO��"�:���x�!߸�ܱmm�'�˔F0�yw+(����~fy������[kZ���n�5�_:��]<<�i���哪L��.�v���\�����[*&Ĕ[���{g�An��Tp?A��W4�g�Ζ0r̋\J\B�����|���7���7����_n���O^�Z��\�L�.J
3��N���aI�;!0in�Va���{��&�����K(�0gd4��|�h:��k�K@�O�d�m��J���h����ʎ�3�l��ZӃ��WV��P5��xئ@ڙ��*v\��gN�g��1 x&�F��'��aE�Vyj�{���>5%�3�vٻ����{`�-N�)d���}꣬m]��P�i�V��<p;�񿴟|������b��usrz�3'�զZ�xH���&�ێ����V����H�����V6�w��x���S��S{j�?�ȼ�_�}Ɣ{��a��yf�M:d)v-:ￛx�Q���*Pp#J��������Q!��V���w��9O�4ϖ���1�>D�S/�����]�������H�%�>]���b��J�[Y�ۥ�sN1�����ݨ�/&0L�sy����/�^�	����*����֪}t�5�]㯉��ޱ��Ah\���ݶf+�3'�bemYEr�� ci�^tdѕ7l0D;o��vi��w��&�T��t!�p5k�K$�د���4ߕ�Ȇ��x�/*���/�����!sDg���~|���ƍ�/f�	a��^j��SiD�J��p+�^�		W��(��Pk��Ly���+[`#{6I���%U�r���R�/o�%vQ��Z/lv1��Q�`�Qv�J�hsrNj�Ϟ2�ц����y�W�c�և2,�K�;F+nʔ{�2J

��3�Hc	�R��$G�BF�n��ϓ	�AO?��.��N\ӶT�y"z?a�м���ߊo�@������~m��a&�b�����[+t�:����@���8�3�����@�#����{8��n�TJ��XbxR���?!�+nIl��1�����wG5�@��uTT��4P_��Q��r~�	�qq[����F4��Q\��ص���ke�������Ҳ!��d�6�:���1kݶu�X1�1����m�v�X��(Q��\U�p���������+Q3���y[�[V�>^HLז�.͛���֚�r�<E�F���i�=v�B|�5��k"���w�����L���Y�ؒ�z��3�{ ^��.��k(S�9O����6�S�([��,�`�]��wN�%����H>�?����|�r����6�L�R4��_h�Ҁ�DG����ǖ���C/�B��j���!���󹓓�r��/&���g�V��e@Ơ\۝�߭�{��Q���=�� �
fo�6��VL�)����K
�WU�-�d���Z��z짶���A'�-���im�#N�h��ݛl�49�`[�����0��=i2
���8z�pk����"�U%�#�d��������5��b�3�@9�V���Bm���N�e���Ύ�'ۣ�1-��=�����l��	�5�;�$5��=���c\�BSH;2�v�1&D-sz�:!Y�]�m�+)ϡ��O���ʚ�w�R����'S�U���~�sh#oߠ6�;7`����ߗ2ͤ<^8����t��H�lL��M�=�����+g���({{�ܱ�k}��3��!ʹ�΁k5�~a4}��!��₭�	d�^�_��:ў�n�$���!j�Y��#��8W��/y=��HKK;��%R�KC�]s��R��C�\�.��9�ݢ���te|/��J���=���8[ xff���X1
7_X�EL:kQ�]#$xS`�l[j�M������*べ��u�������ܱ����;&���lgV���**'C�S�_�O{~�@}eP�3QU]}6�]��v�����ѽ�I��]Z�<�'ݨ<@�`tD��KJ],�̩EO��mʕ_H�D��1U��?NG�hM]�ϱ��\�iK�Z�k��ы�ł�'�W7Co���:�`O�Ng0vvu���Zym��^�;;9U:�d�.V}�H��������d�%Q�����/�ɚX/��Y��8�W{�@�s]�K��5�8��!z���r!]	^w򍍤�Wv����O�a�������<�$�8\�=66�r�Ն�iwW`�fi��v�^�/�����iY�Js�X[g�8�������S����j�Vs�������������h(�^�Q@g/oР���e��� }=��X���й�a=���p-K�����l�z�F)��T�4?ĲdX��O��<k�r�J��>�7����o�=���0���P������J��ö�]j��?C�lM�̩�6��u�PҚR딗��d�n�91���
��eϮ���t-��?R3�S��4����G�YTm8c�N�[�)J�ν������#U�uuuМ|�guqE����b$�-	4����9�jJ2V��Crn���f4+6��>��GP`jjj��õU��?�_�h�>��㙪��k�F���p9�:�����_�ɘ���P�Q�Z��yP���N�S�hjc�ۋM^��t����맇��ˋ�/�,��c��y�,���s6��lv�9����tS�����
`e�]��(]�P����QQlH��� �U/}6ܘ�h��R�9mĘ�d��f�$���4�[i_�]_��)�tw��)��������/x%�߅��T*_O�b�V���}J�س�j@9��1�����#�2��μ��sԎ�l��4��TR �~j5hju�d���|��O4�\`�4���W����0P333#��J���eftv꽯7a�C�&4������@�QhR�6Bj2�~R�i%.&����m�p��N[��[���.���u���� p��sSRO��	`Z]�������tG�?i�����>H&zTKxn���p6(!o�_u��d���:��3���5~ȕ���P��d�i �2d�k8�~Q\]/;���iy��D��_]]��g����� ��ۗ������f���<q8��?�j^'{wgN}}#T���	4s�sV_�\�{Rô$�4Q��{���~�q=�mJ(QU��-���7>�p�a�jUԅ�Zf9=j\؟^ϻ�sK�Q�"f�\k�[���_����ƍV�L������J]G.q(ΰc�^��b�@��D�|�׹\�ܭlI剉�@!��a���gΜ��033�sT�*�� ~/�2�ATWww��pCn.�����yc�����������Y:��glH ��+*)�?{v���,�R,���L&���H�3�b�^l����zzzofX-X�̡�4��dB��v<3���(�>=5777��i��-X��ǂ�%��� �0�2c0|�~Sߓ�t����O�r����ϓ/�Fd��K�`�c��s���z@B?��z����($�A��x#G��nF�:d.� �b��J����V<��Hv&����lgCj�i`���Q˻�űB�m�#Ma��r�TjKu�\�ˍ^��s�$+�Z�A�	��ŕ�/,��1�*��xM9M��G�d��d�A�W,�5�M*��þt������8�\�З'�ي�;׶�|�������(��� tv��ܼ�����&-��?��?5��LWW��/eۮ��/�er�G�:��:- %��y/�<Ew?��j�R����ِWZZ����K��}����ǳGmI�VZ[[�Ԋ~����^=�?��Q'���={����q��{��@����su�N�]����h�$������{N�-��'R����[��ͱ'��q��<Q����Q�B���A��%����n%u��z����͹�v���\~�&ό��o���j���gS`)-��"��	�����9b>�
�OX/�Rh�UBq���3}��J'�����0���'�*  ����^��b/rC���;��/n�L��S�cf`=��Ҍ�-�M�nħ֦�~�c���O��Q }�����H����e(��q	�x��E"��R�|�
᭫���:���߫s�\���y9������(�]��*�S�+=�9�N��瀱��������a�I��{�6~�Ħ�-��Qi���� ��&8���db���p�唕�?~� =ǹ�����Z+/$�O}ȳOT�� yDvnI�Q�X���Yu
f�]���V�5^A5@�u�Β��-3Ù'��@� q�T��g";;� `���v��b��Uy�����.�H,7�ua�[�4��ұ�þ�$��ϋ�a`��P����j�q���[
=#�L��3YJ5Ⱦ(����o���{�x���}�Q��;�Z�K������/ġV�ΥБ���phMΞ�q4�ąTbk����ƛZ�M�� p� ���wOO�l|��ZM�B��!�%ڷ�=�Ll~���5 ��� ��3h߸�֗�h<� ����鹨Cj�t}/zf���̀t4#~���P�!UB�X��6	��K����=���&��,�v���-;�e	�r
��uF�e����`�|���o�O�����P�9�6�W�RI��Q_�m���C�:
�������2ٶ��Z�U��S��\SR��#<L�EJ��y�yM�蟹�}��M�{�4i�2�>�|V4��].�B�y˜[e����"t�q�_W|ȅ!u�U���8��Lmm%55)�_���������Q�D^ޟK��T!���8Y5�����@6����
=���g'�{W57��5U��vil|{��-����/~ �&��⁢Ǐ_��>��T=�����Z"����5��#��>���o�1�J�[Q���|7n��>N�_�	�f�]�Zm��� .�'�$`����!X�Q ���n��5���X�t�z4T?"�T���,��2$��K@g^������h
���X ���r����a�aLH�e��АÓ��p�r�8�rnccc�u$Z9��$�Ӕu؄7� vf``xY+����a��[?��ɇ�V��� `�$a��ڀ�{({�b�����UFɔ����І��Ng����������[)�p;"����ҷkg���|�slM���-�!�a]e��>>�@!��mU�^���0�+�Qs h`����X�J<��c�0�}�]^.@���tfSvi��j���/�Å�[7u�;�GB�WM^@ɿ��Z)8<�7�r�5��8�����,s5��ҷ��,���M�@����;�œt�:���Ҳ�����pN�tT&�}�~mt�(X?[������j�¤k��M���#����+�^~�F\i�]eGj���ߙ�,j�8�|ȍ �իW������d_(q��xω�@���F�~]�^L��������{MK���><-�&�4��4��K�苖٢QQ8���%�cOJ0C��g�12r58����텇��,�pa�o#��絛lJ"�n�>�tF� ����JS>��O�@�2Ny#=�׮#�!�y2eM~�(�,*(�x�?�uU+�=\�������Fȥ;8�{�ahO�'��痖,""�O��Q���'�T �E����h@�^����p5��H&�TV�q�r���\MG�y4w��V�R[�=�b��a�I����qC�U������lH���}�|!�뒂Z�t�6�Ԑ�U�_̢cZ� �����S;�n��.����j�CVҚ'"̊�1RHT�b��죄����Zs��س�I:�R�%U�%�E��섄���)p�;v���g�H��������2��Ѵ�Q��� ߛHUn����@|��(��6�C�Er�^/_uQ`C�7��Y&0p�_��p���P��*dR���u���!>�^������	��k�,�^yM0QΦ��RCbЩۉ:?��6g�Nܱ��򍃜��_�Ϭ���[�93lcE���%^����	�܊�S�ڗ���Ԓ��#-�dX.�j��ȡ8״M�Pj�{��� 9����YYZ:��t����5m���7�&B�B���ˠګ���y�ܚ���*~1�O���j�`*�F��Onz�,sZ
�%A9V�6�,�E�+~��#`�r�6a){�������^,���
(K���f�~���. \���,��ڼUUgۚW8O�z�?���X$�c�B7?~� >��e�5Q�驏yB��Df��I�<�KĎC^��.n�C[�U�xC���g��l�`϶����a��{k@t�	Fxxd��_��h���u�
v���rHc(��z��̣���4����Vm��E�մR�B�02�s
֣�߰��C�lWn�\�S���#H��s�{�>�M6(�B Y8�;�y�>e#�>}��l�(�v��	`�g�%1�y�Kp�T����<Û#'���A���a�!�7~M���o�zj`mt������+t�����X/̞�x��%_Dkjqkj=�y�IJ�Λ�+ŭ���u^�5Slp��mwww�����{�](��G�wG5�m_QP�*
*M�WA�tD)�"�z��Wi��@��Co�ti�w�Z���x�{���;#��:��{���<g��.�H��7���Ձ�'�㇛^G&v�G�z��mV�u���X�A�C>sraX$����f��"*Ɍ/@N�8+����3i�Z}� w�j����g�m����$��;�Ȋ�i�	���˂��l��:�y����0S5��ͅ�Ψx�D��-99y ���M/.5
&H+mDx���y �@^?J � H�p��٩��1�tM5�9�����>�/W\�0���t�ޣ���vu j����>��8$K���A�%�DtC=�&�>Ѡ�?ծ?d=�o��W<_	�P�5!� /����̄�����Q�A� ��ҶṺ�����k�U%L�=$�g1��؏>ܨu���M�}��@�y��
Xxtm#�s=�H�!���&~�r1��=mξ�)S�ֺ��H��a����/�dn*����x����GL6޲X&��ȪC�f��j6p�����FjD�ڜ'�t��S��JJ��O�`_i�kul���5\u&{u���Qo����1Rg�0mVO�� F�sO��6��WQ�jW�^c[(Y�6˱4!����̺�}���WkNM(�
^���<x� �q�$1`��@�;��d��8�.E��;[���t��7:��*��'��#vD+�XEE���u���o�ݲ]��H���'%x�:$�p�m�06��gYh�o����y�Ԫ��Ґ��(]�΄�.gܖ;������ׅ��zd����]�!�`hr2����}˒0X����cڠ>(����U������0������8����%%gr7'CT�� D�:�M`�n���B���W%>��SM�Z��"�[8����Ĭ�ri�ٴo�����^�a�}Խ�*лt�`ƕ���m.:S@��(>*�D!�/�\��ƻ��TB�oo\��^���/�*��Č�2��´_0�����#��&�rUm�r=�X�mOZ��.�a�G���:��Q��Z��獰����6��Q�d�鱩��:��&�Ǐ���WH�~�-�r�z��H�%�&g��5����Tݒ�����*��c����缐z܀Mn����r�@@xʗ�d��2<.r��9˱������mf�!�Ɂx��]��͈s�9�0�]1��"� d0aL�k
&���J��(�U�H `����K���g�� 0j��jmm��~9��t�]�~���a3~&0p�N���o#��P/��H|��4��O��tu�,G�X�����R�PC��i1��p��4"�3��$%�CC,��ׯ�]�s��������C���-�PC��Nn�#ڻ��%�Y��7�.�M��:A���sċ-�>}�/���T_�u���k"�C�<�g\o������ram��5��C�/����o�Ex�nkhh�|�:02�[:ܠ����uh1Wo�b��j�� ׬1bn� p�F �B)h.T�܉�xA�@@,aA?2�Nw�5�%���^�>N�`����8Ghh�j�� ��!�]`�(S�3S9���w�׏����fq�R"�)�:�_	##o?�ց��mYI�1��Lr���0ĬH����	+]��0���O�H�&�~���H��ӻ�}��y!�����@W�������ۿ�ۜk����ȑ����yyK�,�U�;�Z�2��/d�)�$#0���@�X��Je^lF�d���� ��z�.� p,-��D�����e����Y$�6 ހ��w'��A����ېSYY�05LE/����u�.��_�|�~�������0)�N2����RB�"���Xw1q�Sօ��=i��K�3O�JlQ�S��)��-셓���3Ņ2#�;�=@~�R�2��{�qVL}Οh�8��ɿlW���h\�5���["��=x���zl|�9%$56:��d�@�Y�	bl��� y�Z��1����>�[q�����~~���#U�+Z�K�:�:B���TI_���1��rRz� �d<,"�#��ҟ�8A���x� ��J��m�	�� ��k6�2V����D%6!�?p��8�����G4�-]1gC]q��0Pޠ���Kݵ�f-���0�a^2� ��5��v�H�
��Z�n���g�֎�)���/W�h�n#� A:�Q�7���p%wO��i�i��W�e�'��w	s������^#�������hL9`��W�>a�!%~n���_���N���'���k_�C� �P��[G{I������`OU���� ����0�W�*�v�Oy�m�.�.�����$�����A�փ���t�m��ʣ+Cx�%���H�M����Y;���Y{o��������?�����jJ-��U���M)�^��,�n����܄<��FH@��������|�Zr����?�����1�Cx\0l��[� ߸Tݯ�������U!����kxnz-�%V)'V5/�)k��;X�� �ѵ���~�Bj�h�5�F�D�'AE./[g��&�5��@ٍH���D��{N{��`�����"Z�Z�i���h>��	��ar��������f�Cg��Cɉ4�r6D�S.��������i�H�'�o��q�B�D���^����1=;��`,Zjb��(P1��Δ
��w���A�*�����)�i�}O!@mJj�uU�3�у ���O ]]�d�:ұ�~_��Q��Чť%!�#)o�hE�ħ���M�D*�M)����o�~�z��y�P7ˮ�a-�ccЕ����P:|u�B�/~'��|��ˉ.��a�6E�r��::��Smdr��N��ۻ$��?b\p���Kx�LY���H��}Eհ��gFq��9�t�H�È�U��>�C�90�P�&���ob�`�cE�����r������4S�����c�*���l������#�=�=���n]Ā�JO�<���h;b^K4��M��n���E�~�JK�;rr�[bd��Z�I*�:�@59s�iH04���#�_�?t
�����_E_9F��q^W�����ǫF=bcW�Фl��/(Z[/��Z?��Xf^��Dc�g�Z�l�ix��3��L97_^Y[R���٨h<�����SO=���C��[�~WG`��<����6K��tP%ǁ�ʻ�⦧���f)�:&�p�%�1'��� ���А@y�3( 4��1qj�~�\�6kP\�¼c�\���@^A���̃�B�x�I`XbI|Z1�ڴsaK�ƭ�#F�;�7� ���{�_�A�:zR�	�ql Sn��+[�%F��c)��,ĉ�"�I��ib�5�QHz@�^�����O����Ǹ�h��l�=�&�|#�#ZQm��a?�b���ǽ[���h����[f (t�2�P���`��Ʋ�:jH�6�-���?�T�/Xr�9:�51������ˤzڂ7-@���K�䮑,p���"ZP_1�5L~qt�v�~�`��A�ݘ�U0�bg��g��@��}(AQ6 �uz���x�ϩ�)�leK$��^.'��h������%��Ռ��1C	����X�	4����I�B�=�߯/tm�"���P6��wy�Y��բ�D��5H�JLLLZ�o���hUa���&�
��3���Đ�W�o�h�+�G����n��)-8���@��-��7T���y Y_h��w�{��~O�QdpB��S�+Y�آ^??���h6�p�D*]J ~�Do��CgѠM�8µ�����!�=��ߠ����f�x���e{�"$���צ�ѷ��S��r�_Lv"��%�+�7;�oh�m��t�xc�ֽo� ���� |�����@6�K*����hi��m<๧�?���^I�^�j�����v'Hfm���D����Nfff��(�/ο�@`-hN�_�N��F�(�&�/W��p^E1�pQVL>��DT�� R;O)�P�x��
A��'��BD D�O��g+�v��DFxu�"+�?EG���C�4~���BXa!�e*�C{�TU_���&^i,v}�8Bg�4"�U~�<�ژ�J}OKpWB�<&il�8�h8�ڮȚ��jNd�������U�~��1E�3a&$F�"᪭���19�"M�3��	3���+.��ц���옗v	�c3�*<��U�����{���#�jL��%�%�C6�����6��j��+D�2a�}T#-�]-dj1M����Y|�����!�zkfڄlҩ�����bNB����Iָ.��Z��ۮ��<����d�]�1�/��ȯn�C����6���kʋ��|�\RNlQ>�H��W���0�B$����8I�O�w=:�!C���S��#0�j����w<!vހ/��ob/zxgb6��<��L4=a0;�8��|뢙�7h�ǖv�þ~��sO,*_�l`�ZiMI>C�^V<Zb�HI	�{J���uR�o��� lJ��bTN��������C��YZB
/��'L��o��� (K�1Q����'|FE)�|38l8PHj|x�8$.Ņ1~�H�#��x_��o��7����n?�oS�����_�����4,ͼ�&'5mC��j��I�ג��8k��C
 �4�K�I�+*�Q@b�͑�<�%���0JlS6�/~#�g`׵ ($$Cm�]/������aC�,���\zt�(�>*5�
>��|P�H� }?�A4F�;,S��T�p��շ��r̵����U��ۉ��n��dg?���K��@F<i�'	cdt��q2 ���H8Q�K�lF��~���Z�A�a����[��<���lZ�՟*�;]�;���
���̩��+:��ɮ�)������h�/R�?���po<T6H��܎j+�Sb9D��p�z �r\� <$F.�C90��f��}�A*�G�Y��ܘx�H�V�8%o#u��~I��ΗeiQ$L>˳�L�<����")U�ٹol��D � >�~+�;���2�\ ��܄��7x.3�sF�@�6'����Ջ�'�een���Q�ɩ���Lo�*#���C��a�ÍZ��M�!��+����<��D�֣� Ji���|�x�]г����Ӵ����GF\ٮ��g�7Գ\/������Ѧ�<�ĕ,�T
�7
2�+���j���r�!?����A�a�Ļ��Ff��!]�y[$�_@Uv���󒏄W��dhi-^ B�Е�j�X�����p���˲�ϩV(g�{��r�������ld���p3�l�C��R3�h�&�5���u�L���K��Z�Y�w����k�$D���F:���1R��-W ��tFCC�]�7Q��: [�]��^�])?�߀<6>ؕ4[��R��:`D��� �w��}r��T�g�)�{9�6tB�M�9���b�!Կc��<G����@7��*<��\0��9��u�P�?v)�;p*`M|���+������4P��'�����O��6A�7A����<& ��l /�PSg���:͋q��T"f�dvZ�7�^<�f�B�}��N�h��-���&W@Bn���,?<G�T����f���N�i<ف7��%t�o�n)c��G�aVYW�P#:�j<	]Jy��F�Z=� �M��� ���ݨ1Q�`0�1�i��"\\*ܙIR���M�^�HJI$(B�f¨����"�)�S����E�O� ���8�բ
q��  ��t�ˊ��;b��G f����	���2
�O�`�X�s3тt�r2�.�֢G�ՏZ66@UVMU��%��\-�+���&,��![�b�vll��k�r��25���:{�芥�Bv�y��w ��M�y����^�]���4@}���#/��d vO�Ӑmྲྀ7����nnn���^?�g��d7 �����������7��s1�B}b��Ș���i6LB
j�C�� ��1�f��")�F�9T���1ZG�K�ٝ�b�t��������H}��cz��
{�d��f�{�%Ȇ���,�%����ᅊ>���.��� �ʹ,Ɵ�{��f!9O��]����pD\~1�#�q�hG�� ���>)1X�p� =�C�3����L].2�d�b����{�+�w ��m�"��/3��Q�������p���"�n�{�Q��w�s]�����DK/�Fb��B����)�b�p~�W�ϳ?��=.�����$r)�3p���q0ρ��H�O���.��lDmy���1}�)7B6D�R^�=7�G��s ƫH�&i�&x�0���Jv���y��[���E���2mT�F�i������gpY7���Y�C3=U�3��|3�%&:�v�ڪ'�7�STڑPi��ũ� �d~�-�=��[D/� �n�-���:��ބG!�\~��
���#��w���堁<ؗx�sa �-⓳�&q�X[ԭwI���@Ä���ld1�� !���dr4.�ԏiD[ ��)��g�Si_<=ۈ~��i�Zb�q�Ч��I���B<o��9�4d�Ү<%�M4Oi}���̞L1���ڑ�"���R�K�W�}\�yt����c���'Rw�t��<�Ҷ�M���zr��SSW��@Lj�8Y(֝����)���o�N�>��s��BH=˩-�o�L6$�+w߯�獴��٩�$j�~�!c��2��`���?��V�0�*"�'��� ��<s��U%�2��b�2
�AZ�Ԛ9�]2��eh+Y��f��)P�UZ������HHS��Vcv��8���� Oz�J�)��h�����-=ν�����nB.ń	����\�@=ٯQX����!��eL�iJp��;M�$$$�猛
���d� ��oȭ�^�h9>Wf�ۡl����L5�ݏG�)�25#�q�C�6��+��f#u��-�K?�(i��(���گǹ�Y?7O�q?���~�L�x��aw�	��dc�?@a0��C7VSs�F!�w1�����Zm%IH1k7���k��♏L[�؞\o{�Ԧ�Sџ��(�~���ȟ#:o���Xʭɛ�FO"��ҥK�?�0z��}\Q�����-�U!�����+?O����O�#f�9�Nȩ�"�pYcK�)p��c"��q�G	��tP8+++%w��p���s����@�X[[+5\��z9���*z��P6c�;-OPE���9�N�����d��H����>�����˝\Eu������ +��1�6�멹D7�O�@�BM߻�"�U��}����=g�/�ꛨII��gAg�s�h��ʼ��X�([ *��ny����f�U��Ǽ/�r+���2��_��2{n��!�=!��3�.��31{U�����sz�����'�����2\����$Mv���M��$��-�ꀿ��-�|F���D�)��V��X&��A��?�0K>B+0KrcH�=.����oX�B�ܟf���:�E�����1j��'�<uD:�^���P	�+��.����G�?񳶠R�A�րD
&�6�a�>]���Gd<iry��U2�ʻ��u}A}�fȵV��!׆so�@T|���n|]��)���lFkk�Q�����B��
E�ǫ��w�g������R=ryt�����ޱ� �I��ы�ܧ�C]�0�5n��:�f݊Y���mǾ��}ll4��- ��{9��ѓ��Ӗ�F�u�`���d��1 6d��
� �ۄӼ���g����e7��Rm74�F�.A��&p�U$�9����g-x�(�w&���N�E����`�TG{������x_��"���p0��]���G�r�D�ݵ�p�>y���A�om���s�N�[ԊX'\i�\?rTS�կv�2H@�X��.�f���k�����#�l�3������^
%	���E�����>�D��Sr�F��g��� ,����(��������O�"K�A�ӵ�V@�>Cں���?�-��Q�'!;��@���#��5:hM��	�}��g��,'Jd~��c�������_
tC&�.'�)���	�����e33JJ�G�㍏�_r��;��p�]c�?e{m3 JS �p����D���J� a��@�_3F֢��6v�6��������Ϝ >%桫�U�xKe�#G�V;ٯ�b�I<k�D7}qz��q��sj%���������X�+W�dH޻��Μ{� hɍ^��0�R�1[U�ͧ��q�P���'���b`��3>g͂�z�oɓx{�E}}�Ҁ�;}�[�.j9��}�km����w�f���&6�����V's�G]�xP��D���<\��o;U��]��!9����Lv��v����[e�+�o4���}�!�S�\��lE����g(�d
6%�?~,��+C)���'��-��󵩮��]Ko3�A���S��DT��Q������bѦ�"2�	wO��ē��a,���3a�#f�)J9���&�����A�f��΅�ׯ_�?'X"�bxB�K���y�Z�7PnK��5����+s1Y��X]���{)`�<^'0�qp/��_0r����=�(�V���ݟ�i��q=���7(I��c����pw-ޠ3�k�v����>~� s�d�BNT�K���4�{=#�3E���TWdP�)^�w��w[�C��K��X���I|�;�Aҭ@O�X~��vݿ��r���s�6bR�]�a��F���:�#&X�'����qG�RXҬ#Rr1��Q���(he�));i�5��q�kޖ�R���h����[A�]���� ~jqڸ���Z|5#�[?T�HO3w*�l�V��6By���3�)o:[BW�om俼ə�܄�	�U&�j%J��.�bTg��un���R2�=��۷oY���l:��[R�Eﮍ=�ä�u���96!�}��(��}q^����{�k�{ON��b,�&-wl���7���e����{���y��D*��x����M���V�լ�F�5H�Q(�����"�V�����T3�"[!)W�ZZ���K�G�D���@��~�B�n��T6��CRR���p�ѡ(����(|���/pa^��0e���mxEo4�H��j������Y���+g�ҼId������Q�����,��W���9S�,��-��g�3�T��J�)��*]}����!Apq�s����Ϳ�c���Z�|)�|i�(����&:�s�,��²�7J=��eW���ݎ����}��߱W�6�����A �&h�6����X�!*<l��.�'�S>���rc��܏�lB��IO�=����D����a<�z@������ӑ��&�H+@�ThӇ���[&�RD�8J}$YG�<Оy~������=��J��/��qy�q���J���6]}#�u1�|�$�T���	5�'&ބ�`<ˊ��Mx���ڜ�G�!�T	,�����O$���7�1hΐ�_��T��*=a9���+x�� �2vȈ~����Z�Rut�8��B���E������'��}lP�N懺S��G�؎pL�;�u�Ol|�����A��7���v	hh��(]��c`�	6$����9���%NjrU7���B^��7OU~��qN�'hOftƀ�̪>����]h�N�;�6���F<�e�rf��*���0ʌfh)�w�R\�¢RH�$�q.�Qʸ!-'�|z{(��3���6A���F��'��Oz���z)5���K � '�YJ-��;8\U$`�?��Ml����ZR�K�<}D MN�i(lxX�`S�y��`�`̀���Qu;�f�i<��Z�H������~7"<|r���]�3�E#�}TK�`��[��⁷pt��4�b��i�H��.q�����(Qڥ�0 ��r��1��C�����:Gf�'������S����R��O13e�/Hf�����+��/u�G�%8��xυ27f�@�tmrU�7{Xh!��0�,T������<��Vǅ�����Ȏ\(�zC���`e�y�O|���V�矶)ڲ3ߵ�k�Kwؾ`T�/�#��H��}�3����� �F�0x�>�:Ǚ�u}x�G-nM�Y�8G���c���|@�D#�In�/�zT/�*�R�DW��:'�_9�fڗ"d{?�n�S��tݟ�-=�R��������J����(T�aL�q<��r�� ��`*.�b��(F�-Ne�������Z�~������)���T���_&��i]�ϔ]��t� ���]�(
�����Ng�S��<f�Ԗˉ��o�̊�<�����T���rd������>���|��4ہ)l,�1T:��P2d�Lp�}8̧���'�)��Dm����`a�m�s=?N`;��V?��tCSE`=��K��2��Z�-\/�`�GZZX��U�{��%4���Mx75���G���eB��_���a�Ӎ"*ė�,�MR9�{�=�ɇ�_�f�����=��� ��p�?�s䨇}���׬�\��Q]Bm���A���J�W�c	�(��p��wa�Ú�8�-�L�bצC��W�\^�
ag�ߋ]���ͽ�D\�[��{���#���o�ǩC����7�8�tN��k*k/ m�d�H��dPs�*mH�B�H�6�χ�߯�uK�=��Xiz[��c-�6-���o�O���n�G�E����Pl���؅ �f���c��<|/��Ҥ�=��&;��͆����yl<j�뽵�������۵3���{B�03#���3��h�rhĵ=HA��f��)n�޻���b�uo2._���n>�_�5H�QW��C4v՚�8U�wQ/�9EΫA�_2Gsd��~l�_a V}%���8���#w����@t3�^��7�]%�5;�H^�b��3����'�y`~>s�l��FF���#�HǑ'F���p;��5c��o*�1Psˊ|� ͅ� �+c��'�@EtØ%�n��Y_�ڭ�Eaa�R!]��Y72�/ad��aέֺI��1��T�����o��^�i���x�%BY�s4��b�*�q�*$��A����jQ�|�;����'�0V~�!:��s�����)4Y��հ�6�Kgv5��_����c2N�WW�c���S7�d���}񹔆��\M��*�I�Zq�w8%�=&iߧ�?�&�w`��R�e���XA�|Sx������|�]c]o|��/�.��ϜP��ߢП�gԌ��~�m�=��߶�R��]���ӟ���"��x�:��|<����'iy�(48������]��������7��&����
�AbUX1��Y`�=���!�^3�v]�SB�?bD(�&a(�uf!���Vc�+j��a3�H5���U	P��l�p��7�'���|VXHڃc._ׄT��_;y��	��[�%�c-
�}Hۈ	�/HwN%d%�N���0�q�`�y��NK%�e��v����N���<{�����#2q�?�-Fsb@U��(�#�@����}���l����ۜ�n�O�	x*���%yfk�֬�Z���Ϩ�� �*78�Îb�<Z��i_Ȩ��h������k���8�Fq��3`��=Y���p�����R0��갚�ḃy
�ˌ�]W�UT��'!�F$�.��.�!D��U�9.��R�@ڗ����|��
�|����Ӽ��_�>��{_6�nk���j���	�����:A�1���N��_ nK��=����9y����F`;�^`��Ⴔ�B���L�o���՗�4�$�O�s@q�뒵���ꍂZ�%±�0���K) t��WY���R�F��'����������,�t�f�gL��}ڬ��6�6�Є�)��E��
��U�6�8WE�}���au�����y��fMě�l4����/ƙ���QZ??QD��, 
���]���{�L�q�����>?���4v9X�ɝ9������SK��+n�x�a
�d�嫯)�`�r��4�2����˶�ҙ�@R�J����:���������~Bk��(��<��洮����ɯq7�%�vR	�3K4E�c��N��؃�<�U�!�=��M�/���U>9��w���:�|_瑟Y�J�y��l��pw�x���ȓw�M��&�q�~�k�B�����Z�^�m�T�3K�*2H���Z��N�9��u�;a0YN���8���s�s��¢n��J�ez4>}�q��ٿ9*N�xP���*��s�{wAe�byܾt��w��r�bk;m�G����wZ����/���Ο��R�_8x�V��V�q��Z|�N�K���=U�����/�S�oWEF�'"�X������̞Lw��|*ӥ)u�/2+Fq�ǫ!��}�ǽ�z�]�c��AU˺qK����ɒ��3ݱ��нR�u�}�π�7/���]���d�mՁq�c��-��=k��J�٫�5h� ���Y��r$TM+헿ךlƨ��=:����=U�"�n��Pem�p�
1B~�x#��Ke29齙�'��~�H,�V�Ԉ�m�D�	��e�_���Q��5��)�%���;�0�� (��d+����줯�K4E�0��S)�Ǜ���Sw��h����PoI�v��2��#{oI�ԫ���*�;����mh,'�;�S�n�F���lM����՝�ӖC�pVpPj}/Ų���$|a��(}C/'B�؈��OH�jﺾJ������G=0�3��Q��$�zz�]��,nN���R��f�Og������DLC�a��A�ԓ��̡�aȡ��&]����C�� R�����}^��#�����Vg��~Tw��W__K�V�`'�?�>�*r�%���n�M<���p[$��w2?`�7E�zb��`�|�������5P�	��l���bu׷A9���/�$�?cʡ�u�^(~%m-o��6��������%Ѫ�8F$p��*$�|18)h�_�g�Jav��C�Vi~J.vR��7f*_�G�su��ڻ`����s��/��
�|1���*���Q���@�k�T؍��TW�p�W��g����?mP>�`z�y�Gڐ@B�_巣`4���Qۃ�Z�;�-:�1/z1��p�S����JPK%�$�!�������������>���M�W �F߸�����ӡYS���%���":7]�~���>�f찥��3D,����ٰ,p�,@s��`��_/�Vc��%����U��a���Bs��Էa�r�d�c��絭�#�F��L�ۧ��G�2F���
-� u�}a��<�P|g,|AH�!�Ɣij���6��ĉ��V$��]��<6�.7 *��N>��k[�c5,"�u�n`��<5�!5�o�����<d���z�R����P|��8�Ɲ�0���N��$��Q>��z�&.�o/߈�Rئ�'�d,�u�>H+���бƮ$�����^>cC�m̔k��p������U-�,x�L��b��q���o�A?g�������юh���,=3�'`��<��O�ϝ+E��J�,�+[{|�������V��xNF����Gm@����`u�X��o�)�m�����&�P_�,���`�9/C�=�g|ݸN^C�������*�-9.,9$��,������W��OE0Vc��n��k��4 �ԓ/��	&��X,�W�*�r���뻗8�oYG랉A��UBB��V-�#����˜��S_Ɠ��oS�)AH'���Ig�b���O�������`�l���;r�7Ի�:����m�m�:V�jQ@"�ٌ���j��UJ?>n<\Q�wy�X9�|�&��)4�!��2!mw����fO�G��}�����UC��Coķh��Q�mhj���[��s��)`��N�tӗż� �s��OFE�9p�:(�������l_{=�F�?{���_�<�s=s����j��&���R,�#��s��6�ثAM�FEk���"(��*p�p�1��~0�7+d\a���u���������p���*kڂ(5��m��J�3�#"~��?~o�k���ŹXP�Kŀ�Vc���V�fm@���'���Մ�u�@LK��R>�XԻ<*�$Zm��pX�5T��ߢ'm��y��w�B�1�k��²��⓲�ǯE$DN�f���7K
˸���{[/���6�ɝ�����om5��6tⵌ�Dm��*'�K�ޮ���jA�0�P�Ju7�,��;Nq����P�a7,��ȖA�Oٻ�啘�i�32.�����;z��E1U���]X	��������0~7u��N��2�*��{���A1�?o7d���z������v�/�;�h+���-DՌ�"�ޡ�\IG�Ϙ�)�O�j�U7<�j��@K�R!������T'�R�-�������X%�D��][�����ӭX�T4��Y�/�M误u䏓Q�>o^�U��X��vS��h��~���I�`Rt�w�g�͈���Y�����/#�3ƿ��wMx�1Z�����nCF�U�9p	k�=���Zc�Qܺ���ZtR��v�:}Cl��d��4��^_]�Ή����D��2��?s*���֭�Q��9{;l(R��Y�����#L~��P�\��1���%}���c��+�c;:	����/�vm�<d|vC�(O�8�t��˪�&���!���(��B���>�"���;$8흩X��Ŕh�缉޳�C�;�Y�g�p�D���G��V�������O�uy嘘�:,i�׼�䓊�bAz��6�ڿ;84����6�=�*��D>~�c��d&��p�.��P��a���r�U�!~�eͫOi���5Kb������CY0P+�[I��B������_=�U���*i��o�|�pV$���º�L�b5)�Z8Q�4�Vu�z�f�8]u�*�q\JP��J�*�}�0�\K�O0�~��P�����O �qY����o�W+��i_�ܜ���:{ ��mүуL�P�Tx�>�]�0�s�Uf�P9��;�����=��SS�|����r�Λ_�&����&�۞�]�]�l���,�z��C��ɒ��� �͐g��C[_����X��{�J���k��rwN�&�6ė	*��n��A"J�Z#��os7���jy���\�t�:�c��_d���U�-���Qo��fjLP����U�XA4+[�q�Y��b~�����qa��'2h�Ġ�ܻg�e���lY=EA�2����F-{�lZ��l���������w�_R�1�3��>%!�6SE�"��ƹ1���ua�>�xːü�_�3�-;��s%4w͑��1������P�n�}�CJ#~�1���R�E�;�>5Ξ�n}��q��"eK˄�eF�͛�Q~���bU�^���/�:ho�u�p|�w��zk�E���q�a'qO���ɬIcnQ?����"��q]3��R�)l�U�׈%�hD�����V��L�z5�ŧ� ����WC�pZN�gN�М�g���R��ɭ(Y��ΗP�_Z\%.�|"ehV�ST�t8׭��5���~��\��GI�����:�_���Lk'�-�LP>z\ɖ�9ob�D`��/ף2�T��9�:�h�=��ـp���e�z�n������h�T�G��T6�q�̞HY@���jo\���}�����Cv��d�x�.�d%1��S/OK54�$�����G��3�\����.x��y��ͽA�Y��w ��ֲ��US.�D��s�f�?���X�;=����o�0��	��׈&��F�����N�T����@�2�NRt����͡����/)��9s�
��&��Q�u�ǽ��(��l�8��t|��k7��������]��_���ؚɂ%�b/�z?�x���5�'9ƞ��w�N��6n֬;�FZ�Dd��\,�)���ʠeP�O�����^%��SCbڜZ�`m~���r\Q�(.��l`�b�91�8���P<$%q*fz����G���>��QB�*D^q,�M��<�$~���ɇ��R�D&��t_�ת l�2�����mQT)ۅ�u�K�e`AUtQ��б�χ�M���wR<}������u�tZ�[+��
��s�JJ��D"�r�?�0s��{�>^�/���|���,^��(�{y�?���F�H�M������I!���������\�i�h����*��;����N���(Rk�'��a��_��0ń�Ft��t|�8��gz�V)����(�aa^3��mt�L�����]��B��U?1�-���#��%�PoY}�{��6�cOQ�/�41�f�Ǧ�ecg��l�>2j�Z;i?��WqǓx���'ٵL<� �U�e+�1J�K�T���R�;D�Ƞ)-��wF�Z+U\,eMd֏4�_8MV�)o��o�m��� |��!2��ߒ)C;eP�®�k�[m,�T�)3�V�6�?>�y6�3vA���;���܅�ѥ��*�8�^�5V���{�;��K�	zП�n��u��y025���/V6HvƿQYu�����C弟�`N����1K������,I<9���|�z�����w�a�(1�ŭ���vy�d����]o�'R�`�k]X%V��%�JQgn	�#��U����N�l�����ܢ�ء�<�JfE����,��L��"�h�EW��@���9�pNe�.Z�j65�ٖ����:�I�R�����b�ȱ�����[���O�ڤ��y�L���E�~���,�h�N�N���PR�{��Ĉ�`������Y���7��qUV��{w
b~jr�
���u��-�i�:�9d�.)��+����eۈNt���Vqvtnw��V�3F�u�=m`N���Z#��|�7\�[��`�X>͇yWMl��0V�9l����t�M�g�r��ʨ��O���0'�)W�j��v��\��M���V�/�(��<ȃ$M�Мq�ʥr�%�U'�s@�%��ѣ݀�elˏn��,9.V7�z�S~L*��O�_ �N׌vo^+5Aw1�k���#yS���wh6���	�9_�ԕ\�u�$��o 7��I5���GQ����+ 9�QrO��ڟ	hH�}��/��\��x��2o�� ��i	��j?d�u���X��%!ɚ��c�p���>s���En�0��$8N�=�M��k�[��T��>�쥈��×
��m]�)~�H��ȑ�~�b1O��:˱�����>X��8����������lf ���{ϰ(� \E�EPTT�
"�!LdQ���$�!��dA@�"   9*I�HF���3[���{���{w/�9g`���ꪷު���\&�ڦ��������~��˹��
�'���W8�O�RE�ei�tI�ı��]��g��ʝ��^e�g)ݫr��+��gq�d��%@�C-����5���n:�|�+W�MC�BSV~hI��+6B��@���%���A��Ky�'�+||��~ϟ�^�ksJd�d{z�D%z{�'O����[�-y/L'Vx��2�P�-�y�}��,Ǵߵ���6�4H5Tb���L�$ne���b�Z$�{3R+I!�z�����'�m��UV������ Ý���u��S3�nʞܬGq��Z5�M܏U�5����%��W|�`�v��<n�����薈k���}_��W�3S��<P6����d�VVi� ���m��.��=����h,�����S��W�B�OP;�`lmCU����뫻W�i���lJM�5�уC�ɿ5�y��gR3|�����+�f�����3\[�?ݳ�=r�}���������']/)���[�fh���Ҩ�M���SO���[��h�W��� ���a%٥lǕKvo�V�P}|������k��n<2�U��S?W��s�����V����'Nd�o> ��(��[g��K�9�L_�2���-H$���S�e��i�J�9nm��F���<��%�W^��\���\z֢z��}�=�IA�{雗��!��
�6����Q�z(7��5Z2\�bR���M����w���X��	�Hާr>��+c�ƭ��L >t��FM�`�E��^�k���_G���J��zs�rd �7��-�Z�Oj�4[�<�yJ�����V�Xu�n��m��ʢ��ql�-"����FW����7�טZ�,�5�,�FƖ���g(��nm�z��=9*}C��<��'�i��mO���di�Bj�q,%т9o	��v��_}�"�JhD}`�_��t0�|S�"[��&� �>�+��W�S歼�C�s��2ç=���q��h�+;!�m�����r�����I6�����X��Ӣ�OE���|`����͂ڝ�RKL3$���O�
��Szn�ޓ!�ם"��[�[S~O��%H�ɋc��'�N
_�M��Y�t�|U~N�]�߉j��;3Gy�;�Rۑ�� [�K�7�6�A�%eu?���h	���^n�:'�5���#�3��+j�4x�F���GG ń��+�5�O8.���������k�o��D2�{�E|g���{wi���,4~����y ��� ��:��/χ L7\�7����J���3|K�D�5ǹ�Ж�gT|�z���x��hZy^�0�Ǚ�u�=��o��~�n@p�͎fhd�j�56�h}�r(���7��}�fRʂ�Ck��e~o�++,}o���vxqP;��U�����ǹgߙ�O,׷����������N�;V%:n����8�asنr׾0���ë�[vd8�����.vd��u�E�K���1y��RH��.�ĩ���*��7<si������wr�I0��ZQ�ڼ���Ϲq���� ��[�4:�}N�[/z/��s�Ӊ�It�dN�*�n/�̻0�f�{O�]ɍ�����
��D��-[6f�F��2��?�>V��'��NX��$�(s�ߥLz�=l�<�6f��#~׾/����zG<|4b�\=�E
]��Ќ���<|�b����Sz������a�ƽ��_9�}����bQ�ѦS7�͟�S�h�;e7I��v��;�O���^J����o�K���͙'�]X��+���?���S.�����H�:�w%��;4J8Q�?y�|���ע�!�&X�Lh�o[!?P�lq�C�Oݏӹ�'�D�}J�9=��</}e���w���}O�};rY�e]�3��l0��Q����}�ޘךϔ�KZkr���Nq2�_z�p,�߲���,�������	'�H��>�]s}��9��[����W��W��On��sU�n&m�������:�g�K.�,VtF{�*01�-Ŝ^C�Z�ރ��5�oH���O�V��t�|�ؒ�woU�>�c��?]J&�=��d��|q�pCV��v������_�z�L�U����l7��&�]�!%ٝ~_�������+�ϾԴ[5�mE5`���뗛��ľo?�m��Ή�į�*?����۱:xF�髯��"����Jc�e���ON�#�������}ږMۙ<n�\:yl#��MΒ�y�?]�,f�1��ʱ͗_��sYS��_1��s�(�۶���fP�N~�4L5��V]�RH,�7,<�����F�&���I��w���AJ�geVӺ:�퇍i½F
�%
Dw$�7��(��c�"M�;�%
��sVT�Z,pqCyKsó�;�N�J�Q�
��J&1�<m�*QN����#�t�~Z������[ڛl��Ժ�R��9���3�c�����LVsg���5�=V���:h|"��zL<I�?X7H�~JpLs�̴\hg>4d�h��3Y����K	��{(a�E���M�6�#��b��	�ܶ��_�����J��H�*�����[2�.�ʝZ�d\�M��,�pƑr,����ˮ�+#�������{��������]|���A@E�5�F�hOE�81qo�b,�.>�k4�G9f��{�ݗC�
��R�:��D��S�i�GJ�56m9�1E�x�tT������7SRJ�x9��hIF����S'f����9T����b|�j�S������ܙ�./�/���O�s?8á��c�N��n͍r?����~����S"@a��]���ゃ��*�^`6���
�S�5\���F�sg�<�l�ݶ�j��
5)s�ۖ�z>��d��n�8��c��@���޸����.�d�"��9�C9��?��fi����J�Y8�{�&�J����9	�iŜ���#�&�<-�8���^����,��Plq�>�lyZ�~�H��Z�-�cm�6+�3�q�z1er��Q�Q�������D���T��kdJ�vf�>X��<�T/T)6\ju	��d*&���L9�;�30��ޮf�MC���mU]Z�!�J��}�-������Z��à�Z'�A�e��n�!1N�)�������� /L�9{�!!�^��3l�Y���.'ǩji��2�ތ��v����X�<�9�:��n����Ie7)�����Ws6H(�f����MY�Vs�¸���a�3�}�G���˴^�t�՚�/w����۟�2�,�qϲޜ�&�����|E��vYtC�n˔�)A��M-�-�5����H���]��`�i)~Gmqt7���;��2y��Ȼ�ߕe�Q�dO�u�p�гTt7����	�B�吗�����К������6*4&
W0u̴j��|籤��(I*u���>Q���+vw�^�u�mlc6�� �M�F)�������em݆��w�#��i�M�F��H��U����e�����FB~	^�����NL���j-�`Z����c���c&���6$��3L�LԪ���h/;LFv��z�}9}���g����$z7�*�פ���
�+��O������7�?�4r@�5e��m��N˦a2���]�?M���1�'�u@J���8Q#x�;[�}~�5�V뇅���WW��R����$u�:yTװ°yOot��^��-hL�<�n��M�Gh*��d��-n�[�Qy�o����>
�b0�ْ+4�B���@q.p�e�g�=����[�lI:����c��;9�i�bI�N;�l���������P�tQ4҃i��$oF��_'��~�uS�}���`&���Mf(��{;���P���gϲ߾��}�t��g�6?\X�L%=%Vkx�e��Ȝb2��r$W�s�G?H�ّ�2��W��'M��i`y����!�o?��3"��?������$��Ӣ"�5�R��]Ф��]-�nl�J=�k��̍�M��d3�:[�4�<�����Б$�7_���������<cf��V܆��P��3���C7Zw5��j�(`�f�d#�N�0{�Շ��֎�*��\��%�J�zu�GD�TFp2�Ns�VG\ԃ��־�c,e�������^�`������6�Qy��u	�_��Qޫ ����{��y�"y��*S�p	Ec��g����7������(�?!�yg�-�����ݯ�����+ct3[H-�Nw�>����^Pʗ��H\"MńgK3zn#<g��$�#��ډ�훇�=��2�6�����!\o��f����*+�����;]/^p�1L���53:���4Ϛ�:MZX�$�D�����	�C5�	�Ő�6�)I�_�A�~��&�~������;Z������I�؃j,#�:D����saN�V:9����ī��J��_�d�|Wj�2�>��mԈ�E]�~5�g��J�ͭ� E���j�ڷ��Bݐ�V�@�|�u�P�nv�k4�:H�)U��G�)�vɐ}��L�M��k�!)8�����st�;Ty����=)�3� �Q/�'V��^���gk��q�B�L����P������|�iG6l��oQZ&�~a����{����w��3Z��;��fw*�i�Kp�Շ�˯��ߋEI_����M��F-�]�v�)�mF*�Z���.�0�T����g��E;�?j���|cMgǴ�ˡ_�5��>E������o��Ye�33�H??���l�i��5�xp �)����?_�F��g*�g��rMp�;�Ln�d�2�MQ��z�&��|��Z8��ģ��ޟ���	;�w����ۆ|`�ܞ�J�d����E�]�_��N��o�������]^�.�O��'h�z��X��u��"�E��\�.r]��U�+Uq���|�xjP�g��G�{~�����O��?�Z���i�����O��?�Z���i�����_rjLL���Y8�q�s{���[g�Pܣ,xGⱑ��wS��iՅ�މ��ֺqqI&{k*=��:��w��S��������T����x�ߒ��~����,��������u����\�.p]��u������U�G�	�#�b��ȓ>~��ӄ�F���1S6	�o�"�����y�>��t?��(&�md��]����2�8,���L4,Mx��Г�ݽ83S��}Bȫ��S�P�|7�͓��V�D�i�H�Ȭ�Z�xTEO��e��,6MU6J����2U�`J��l��ϯ�eU�.p]��,0�?��]6��5��3��RV�%�Wv�;,�\�������̛%�/�g�_�5�1]֤>�g��1�ǉy�B�sU��|��ݨ��v�8���#}�������Y�����br����ݪ|�̌q��k\�.r]��u��"�E��\�.r]��u��"������ �o��gb���Lmm����Jm]�%{������a[��Xm}}����B�b��*�鮮����\	�� .��� .JJ���>~�~�7B�g���.Z�k^����7 i�E�8w�N�g��[{<<<�~~�/�����+./_3�0??��cPa���Ϙ�(� TTT���虐�p��A75����t0��9�����c�߬�����ի��������ׯ���	��(��������S��TWW��:p��0Hx1x0Ix|~��k�g��h��ٟ�;��6 ����64�c�>��~JN�dkk�)�>~M}�%�RU�16߫�||fff�x|���,�4)O/hβ�A�@����`{��A�F�mҮ`�dɻ���X��U����xCMMm�×l��zz.h13m�LG;[��LgG6fZ����[�.�|����Naئ.�677���:WVV����4J;r��\uһ�����V77�y	�_s��(l˶�
4�qiʹ,N�(ަJz������6G+�%�oJDC��i�_�	���6h�52���mc�\�|�zC�J���0�Iǹ78˸^�ձ�E�8�=�N�Ŵ�P�z�ko_�K�Y�~a=q߫����9Ϝ�S���f$l�^$��*���F2���;������LNM]266V6-�wI��XwE ���Ru{;�NU���쯗ҝ1�9��˳�֤�������bѠ��jN��ąߎ�/�"*{3<3���ٕ���Ƒ3{Tda0�1�XVJ-LzI��A��(4K�o%iK~������c��Yk�E�Qk2Zi�%n�p����%i��;���'t�PʹZ�M��W�+Oҳ{�f�:]�;Ǌ�T2�[���������E�|we7ڣ3]����08����}�+�|�����HfOz��8�aw/�ypL�I���;���8�v��0r�`�綱�Wf�~v�|(������ܯ�cs=���C?��O��_}xT{X/V.J,Vh�Q���Mu�~�Myy*��8p�?5�;�F#�+9�����9b0V#����{R���J��A�R����;ev	d�SS����`w�s�����
ܙ�ƽ�lmm����000�6��Ps�I�#��->w9��ʪ�3���B�.IKKM��'��}�9���Z���M���y(�Z�uHPa�����M��1�XĦ}�&�)5�F��^�����lPs�<����N�3u���D�#�@�g�/^����l�cӕ���_/���r���$�R�ӥ��m��$iW�N4���S�u�x��2�\!

���ݢ�q$u�)_��:|����:Щ��S��[�8Um��hU��
�ۼ{�K��D�U�@��/O����XJ-��9x������0�Ϋ���p�̞is�M�/�Y}z�����@~~�i�$�>aR�y�����:E�C�<�B+����-a=y�5�>� >���f̥*x�aa/B�ͷ���vGQ�F� r�h����;�[Y�e�������9@R��?������W�up�r��������E���B�-����Ѐ��{��"�6�܌A��3��%�%��m�l��K�Sc݁�E<����09M�c�8�T'I��{�޹P����~j�����n�t��]O�I)��;�S��F�!ŹRX5���l��v�v{�j���6��h> ����۪h��w���?^WSCe�=u��0��mߩ�.��.Dʫy')+/3������a�f�,((�D��(L/W�cojty�]����׵�/f���$�L��E�~��m׽`Gr��gQ�܌e�ٶ薍ۙ�xf"�>�bͅ2��M�g�n*�,��aQ�U�/�� ��5ި�}/��\/��լ)�<��}%ZN�%JS���{�^-YY��'{����yfݞU"FE=�^%Peq�����~lz}f�UKz��U�I�<bo�J*I֔���i2�S���/w�ªu@Տ���^�����ʤ4���["(��d���0ĩ_�~���ɉ�*�;��<����[�@���U��l7;
_��C��i7d��v�1�֚�TΠM�)T�!�S[�o����H�L�n��lsC����vUH�fnN�Ѓ�O��M�T�����Ӹ�t_��J�����/؛��h��S��~�	KN��ne~��}�>U}�1��u��ϋ�/���ܯ�<�����:��-���E�~��=�2zʗ�Ҟ@���:��J&q͵��܁L%��k������A���wg��g�s��ͮ�Io��.�ğ�*��2�4����e#s���}r����eذ����.�P����GJ�7��I�
�lŷ�$��N�|H�d��@��[�K�DO
���:��{�awF��fy�WY�#2��^�mMK�b�>=h䬔���s.J���fө:E���Ϣ�T}1�3�m���O[��
��i�%�?��D����A)��1��]<��ͷr.������k
�݇��-���ݰY��~]<��(�L����8����Л�n=�[2 �w��st��9JcnaQ1�q��݁)� 0S	SR&X��!6&&�H�k�>}�$����tT�[�y������8�{�bǁ��+��x�F;f��r�U,nd�~��D�N����%D�_�CM�rvn̰0@�l�˫�JZ��Jh����� ��>UZ\jJJѷЋ��e9�Z���g�W�e��/]sS;��h�X!���������xR�COy�PP��|C�H��t�����奅�.���0؍~nL3�+�B����Tc������T ������_s���|M-���2u��v�3�ť�{����_׼�	s-+%v�/��+Y<h��8�c���pQ[�WL0�*�R<_{���tg½���+���v{qU�3U�F��gZ�4`B.O*F��8� S��������������0����{m��������� �3#UR���B��Ϯ| R��A� LT��J	�Ef���^�S�7i!R��2�a֨�▆{�5�ű[i&������3t+o�A%�7gy*��������N#>x��T����S ��Jݠl&ini�g�m�.Q�E�mA���75�:tȴ�`Y�'��;""�F-V�GV�ԁS�kW�������$��eO7ϖ*�xH!)�5�NO	��Τ���(A���3��n4�K3:=��[v@�ޔ���˪}���v5�bl�
�H`�≛q��v-Do���]�[��Ew�!�
r�����ٹ*G��ed]������N���u��ҿ�{�8�HU!$4~����X����%����o������
^�n2����:ؒΕ3�a\PH�F�,+x%.��N!~���*q�hk��X�,���9�KDx�xx�bX�g{�)���O����R@zh7b��v�#�Bc0"�x�|H`��m��I)m�:�A�e��:,��?M���N�x�������w�oލ�9����Y�,�3�M$��Un}x�G_��hG���EE��*-�u�}hT������b@�^J������q.��/Q�8��)���W{�oOň�瑟�A��񘋴X��}�<]Qg�[ס+	l���=>��ZG,���5#��k�E���<-5I��w�\��;s��M�ԇ��vghR⒳��Ei!5*�d}K�YE�.��*v6�WT����wZ�8M��vק��������J�����d����-�=q���~)k�~�m�ɛ���� X�|mꢽV!{��JA�7s�� c����e��vl= ɢ9~��]�N���(m�;�l��2�@>R�#5{Ȱ�vu�QZ@�sWv�%c�|��𸡶lfٖ9��u�MY�Bf+:_���z2ι���.2NŬ��Ӽ�� �M��I(
�D��.Ͽ��tu��Mo�l`�\�d��m�:�%=N�g�}u��+�\*�.�HIkf��Tٌ��7���yN�bQV����1���-������b�W��TLuM�K��_��;�+/�V����VU���J9I\���`fG��ҫ��4�fm��0<R�h��0�N\�BL�lc�H��(T{�]�i[񯒗0�w����|����"M�h��-�&ʹ�X-t:\�J$m��7��!t*C&;�w�}Vܮ�^R��O38��P���D5�'c �A��#������h-�ތ)�]��[xȲ��Gc�����%��<rC"�������ۗc�o��pRU��$�~yJm�'geiD'�~��P���!�6qo�򸼔���egl!�F� ��WIJ���Lt��b3�*����0��r|�u��`f ��`�9 *��w��)��4�R�� '�;
;��Y�"ӻ��R�"WE��g�۲��"`���T,[����K�<���Q��^��y���N���P�R@����=��J;��`�s��~a����{��Q�f��kF�����6\:��[�Nh��>9�����s��JP%��������^�u��寉!22�t���B�Q�M<	U-@<�
���|�e�㭳c]]����$y;&^���ug��� �q���s�A^M��V:ƹ��t������kz�y�v�;�9�^�u~��{,8����B���޾��+<���4@�$��`��.>��� ��Dۇ�� ��J5�~�WV^���*:?����]�\0�{i3؎*�M�Q�ɞ���f�7���X���o�%q�y0vW�SE�NI�>�cjEح\{<��00~�#�E�4�W��N!'[���Z�N$uQe������
�Ri7��^Q���/*�N@�8����Rǵ+��I�B��1��Z����dM�����J��������:��eI��d���,���{R��T��a�1*�%r��3��8z���/h��g���l�%�m��ݹQ��q�0�1�bL]�@#W�L�Vd�i�j��i����P&j��	��({���B!�Xz�=�~�m�U� .�"H��P������`,,1U4'h�}�D���v$�02XS'R��a�\����91'Ǘ͊;"{K��f�H�@u��2wA/�;��z�6	�d���혧`�{]c���I&?��J5ė�E��I>��.���r����΍ahq����Cy�E'̱�xGP̉����>i����!cG[��Uq!rB!0��*戹�*���Ҳʐ�V��رr�*Mj#�I���W1��:�iy�`Rl�UK�by��֐I��fMF�I�r���7�m�թ���Ԣ@�:Ss����:��%��?Q��jɣC6�,�b��)�b��<d6Q�WiA׶�W��[��"c���Rx�Ĺ�?�{R欗��-;�WU�,-���W����@{��t"f�V�7]��Ѿn����2依=��ږ�� w��pKz�VV�M n~�������>V�6[ħͼ*��/lYo�ԡ30�Ŏ-M[}Z�!�'rm���)z/�f�������TȀ ;t͏<����`7,
��e�ܹmܜ�1߭�����<�2x�|;���~U���V,�j�P�����3�$ˤX�c��!4ю�jev��*�����4.��� :u}��*���;.̂�6䦂��/ʞ�6H���>�|皟
$Ȧ/�bn�:ʜ��:��L��2��k�Ɛ`�~�'���O �*{���|+�����h~�Z~���A¸��!�^x�N�}�, pX3�?1�>ɀ|�t/`�vz��s����W���	d��@�"ޡ�]�UYH���[OHR��I��⡂8��THJ���!R �{�.PE����hs�%�t�K�X�y��!�VP�ؗ� U.q��Vu۩�=�
ZP��)~��%�kc5��ܸ�3\��X��G����s8�}�w���Pk&_�%�E�~I���NNN�T���Sa�FaV�)��>�Kj�@���:����H����8A�8��_%0�������˶ ���R���\��?��S����}2igU��	��?��K�uvX�/�y�'j�Ĩ�|��H�;K���+��҈�A�����&���VL��Q|��ҡ���]��o�b�,D:�j���`�T�?���W��rQ����d����mY�_�ì6�S���)���0�0SW��뫫_�ri��5�|�i};r�z*QIO�������v�+֬J���Pq�|U6pv����[�+Y
�0�����P�g"~�#�v�0Þ�fX4m5iO1�`^��[���n�Xd�)�x=#����L���_/��*@`��ǻa�Ϊ���ޞ�a^�:
�f�3��[$l����\�Ji^��,]���dMt��{�˫J��g`��%:�����:��8�@�gF]7"��c��xh�n"W��� ��}�G��^ù+˫��"�Y��p	�J��9�^ ��y������}��$o�
A�3�QYe��A𓸴NW��_u�d�`'_�s����� �
=��ӟ@\������9J�/�*�D�sdϴ�9�P1=?r1�k�rAA�D��׃E����ag(r�#����!�Xܥ�Оc�ը��_�iE�9�ҢJxF��:�vlQ_dp��l�C[�T,)$���F�,����[	GsH>�/�T�R2��%���a�79��A���.&�d\��ᩞ��=O�I��:qC�_!2�F��(�I2�qV�q��zZ������ TW)�e3-G<1+�V�d�ikֿ�n4:�fړ#�8���0Hp2��O����P��6��|.�}�ɜ�zs ��+�#+�#��rK�P(#�c5���%Q}G��F��Rs1���3�h�JZ��,;��̫W����Yє�M{�D�u��ϪE>��\�3]+�щP��+�'Nlt˟q䥅}a�Μ�a7T�]�GJUHuG�X ��Mz�Z�&Z��E��`��m�#���섩�I�K�*�Q􍓮K3��S��o��*�ܤ����I�Q�$X8��uG�y�w,���ϴPi���rR5[Y�Ꜭ���x�TwTd���A> �|ƪ���Ӯ�B�w���?b�d�;P��;Z��
˃�zy�*�X
��]�����`V	���,��皶�9.�a<nu^���}� �� 6Ѝj�qqq�;zy�vxAz"�e<�N#{���2
�H�����Ӱ��P	j�+�<CګM���T(`p	����n_ �a)��|"��VT�ƒ?�\��x��B����� ��Taʫ<dV�	q�f�/2�*�!V%�e��d}�Y/��� *��ɒJ��3�ˋ0#~й}��o5��]à_P�3Bx��1��j�]��=K+;�����X@"��!�J�	���k9��,t��`F�g���W��SIh��m �92�"���������Ǖ%��R��'+U	��m[`}H�*p[Ѣ�*�S�����T�JƄ�A�GT���G�"��^��}��M��]}�y`���@=�Ѕ#��G��"5�ei@�a�A���d�o�BbP�Y����,�	\C�HW�����'�AQgM"O�.�`N���(��\��D �+]~.�~w�_0ѯ|��d�`{��X
����aT�����Ɯ��
f��zG.�)5�oZgzW�3R�Yv����4-�#m����b@��\Ǖ|F�x
���v�=�l�?�H�NÈ>s;):$S��e�D��j�fO��\�D���@m��Y\GG�j6��JBL'AgMەW��emT��*�����t0 �i�����Ge�y/`֍�m��Pe+'�^Ǫa�{h�G��	!`[_6���%Z��@��N/�������-��kpGR��lU��`�n�lx�Z���/��W��*԰d;�μ��3(E"f�a������"Ff,>�E�a�o[�QصZ�.`���gF�	���qz����S��D>�#Яt�ݯ0=���U���j��o�M4Lg��@��☌�շ{5�=+*;�P�����9��o��K@i�Dl�rxNl����~uq~`��ZRM>Zc�L��9�ꅮ�0_�+��ܬ^�N������"��^C+��"��BEn�% �`�n���4X���YM\-!9]T�KF��?Q�D�j�.~#u��A# 䁴�\TrP�����RI�����`��2A.Dd�ΘCyN!*#,,�KKT6�3�w\���]�- gi��5"ՐW�Rk��o%j^!��6���������m�6�>�b�+���3Wj�l�@�۱�뭵?��^?� ,B��h���Q��tb~q3*��ٲ�
\�4&{��h���X)�H�t�JT�-u�h�$�����vt|~���ݹ�AWH91a�>n$��~�@\�����o��X�m"
��DſI+��}��;�aO��^x�`��U@?�I��ۧԚl��W���/7&h�Q��Lvzq�S�{�pZ�l�j9�]�)��zdSwQ��B(�	7R����":����W�*�	/��
��APS=�`)�P�Yl4]�cA�%�T��"���yZ���f���l�\j7�V��'�l��A���>���BZZ�A�0��K��w0SwC*P;��Lf;8��dMO�5DuzJXWx��~2��%1l ��~���=�b�(b��E�N���^�������PӏN�P�]�Θ]&�������#�k׮�r⮓π��c�$.~1���K�.�w�4p�#��O�f�l�Y��$�Q,��ɨ3�f��$�J?	��Ѩed��c8�]�k{{{���v=&�k�Ζ��?����>�p�T��J�/���;׃J��o{��� �Bd��լ�q�v1�Cd���Iim�J�6[�eY�<�Q<��-�b�N�}��s���аi����*&ƧP}����B2L�CI���ݺ�{��D�9! ��τD�����3E��	��fT�k�u����}WX���3RX6�'�H�~2�#������s�:���  KK����]��$.B�&�t`	��?l�8*PP�!D	=C1�S��t��D7���Vn�;)׽��"ĽeZ�<����>�����顐��^>��}��t�&� .mx���p���a�Lm�,iG6�F6j����;*����SJ�����' ���	��tU��o�b��˨'�/�m���k�>z���ն�U�]��Q���+!��f�C,ot<��{螘�G� ^� R;��@�n�yq
�
O�{�8}-��!����1C������fj��U�Ċ+q��-�����C�V�$`|�THxV���G_��h����V:�N)�ݲ��|��x>`�%��љ^�L�ӝ@/�<$ȍ5�҃`� QvȬ���5p�����y �9�VW�K\g��u��8]Xe��j^�o��S��@ǆ͟w�&�ο{����gZ�V34��Ds�6� z�;wrK����P_-��Rq>���p�b�२���R:��XQ�J���m�RQ������F����`Gb]B�����T>S{�Q��h��ÏpZ\0����R����L��O7��x��?}8�#�8�b�����N���C8�����D���c
��j܁���?u"���kѥ��.%<U:�/m$��y������o��?�M��<�ǠP���B��Tx2��蚘#���_d�RY�A=�� ��L���g�3L���}���T(_�t����~�5�����܈UJȈ�N��㶼rt���pSfXt�c��r5F�s��7~��~ ���j�4��Lf?V�##2���E���P�Ox渲ܴ��p��[���Rr?O�E@��S��Vߐ�sC[?BE|f��͖�a�^���_eA��Q��O5�o-]�z@�+IaB�X���.��n��Lo������(E��8��(ۍ��h�'��t�^LQ�e��'N��)q2b��C�ܟ�K���X�;+��디��M���>(�4�+��j�UtDP��6v$Q�l^���b�s�zo`���u��n�tJT�e �p����c��� �Fg���͍X@[�Ȇx�=<�y�l�3��.�^�b�9u2��K3���%��,���yc���ym�%NH|�(�+�ؙOB�,���x��:V6w��:��dc�LW��Hd�c���
Ԕ)�ho�G�IЭ���1�U��##�e�8�|������2lQ籨*�jX�ܦ�X�M��B�� <����{�N�9�Wو!�c�o����AF$�!~9��1�1!���vz3.e�4o���N�6���EPU�3x#�#�����cJ�	�rD�����S��E�$_���d�>���߉�3��k7�(��uэ��D��b�9�4?�*�:���d���! U���'��b̏����`���
�%d,--O�I9�5^�F���v�ޓH( ���o�>T�n�����TYZ����h;�32o�����aM�j���{�S���,�&��3{�p�%��� �l�����O͙�m�j���=�c�t����5�a=�,�Ļ27s$)@߉(����E��ag0.�@�������بc糬;ZX���mo�W%li�D.��s��[�C�Cݱ/�$�;ܳm�l�U����q`J����W��������UR�HC�Q����/�e+�}q<� �W��m�Q~N�U��X����P�9"*;^�Z�c���#��OU��6�ӨC*ܶ�N���¼l�f�2����6�; P��A�PC��`77�����%�@�L�IÖ��@ �z�ԡ�.�xk�M�c�Jm�K}X����CҀ�a�>���7~	��b%�q[��&�m����bv�F��;��vgq�&u�<��+�0�L�J� 9��e��i��o�C䨙�an�I��ڹX�.��:���E��N��,��6:A��'�k	96�9b�:>�ժ��g�8M;wX]B݄8����*gM����3��t|8_axLuR1��JbC~H<�Î[��S�&�=������7�I.��~E�M�O�Kҩ��qQ��C�m�Qi��_���]ѡ�i���#�`l���|�.����V�P"�3�̛�z��^7d� ���$ v�f�m�~�\W�~�e�3��]!�հ�]K#@U�U�>g��N͏�� �o��v�p$"m .��q#�76G���A�g6(_�l_�4�.X�֕��Nv]�JBuC���?�N0�^}+���V��9�ٗ��g�u1��oXO0A��W�s�?U0���(B�u(*%5U���&ԡOܢ����f���:�Z�A��u�C�(2��K��x+,�5�&�>�Z;�|L�X?0��_���U�v!F�X�\H���8.�qj��-�B�B9.�HZ��.tq��S�ڂv�k_���'�?;G[vĬ8d=��ܹ
c ���$w/��O�zN�>�l���y�LP��+BJV��ٶ���Hݎ���d洚��#��6�x��6�m���^����3��!v2��P��EW;�D侳�x[�x���9��)�j/=��h����'4�a4qy�-|��nk��ßSCO�3��1�8#q(Q���{��0�`��D�B�Q�^R�b'u�|md"�*�n��6���A1M@�O |�#AC�Ųݞ䫇�4U��{�_�ӧO��Z4h�Ȩ�ԉ���џ�I�t�ۇ'Z�uʉԞ!�b@���Η�������h$���O+%F�j��M��F�'q�D�F��򀗄��;Z��~���ܬ�: h��w��Ϳ#i:��F��5�F�+�u�j�,��ǌ�q�^<��	Gp��b����:Z�>j��C�S$#���q��>~�Y{���~����-�=��;w`y7څdo^{u����`fF�o��tbJ�Ψs�V?��R��R�Fi����yԞ�A!�)��%���E෡��"k����iw $���
�pd ����w{*	��+�<<w��^Β�Ld2�_�L��e���y�L�v�/�Y]��	˖�R ���hy+�m�J*�3ˎ�N��o��5콳�E��m\��:����K�7
�>V�6("�d� �J_�U)o^�f}��ia�.'�~��(�;w��91Y��ڧ팑c��6��T�-,���~ZV�|�h�9�F��S���D��*u7L�~���o�NI-�iP~I��B���G`�Xs�2���_w�x[CK���X*
?"A�#L��r��%S+�.@���@����+��M�<@aޠ���"�w�(v3�Өٙ�)��}�[.��$޳�3�
�tՀ��s%҉\�QK��T�4���U��d��TJE������X����Xq���:OA�q�A>#��a}'�����n�rN돎�5�7�S�t��K�`�����9yO�ׄsވ�`�)ٴt�q�lQ׮:��b��O4�m
9�������l�U�Aw�р*��t �����N���7`�Z����,�
NyO��u<���`f�۵��~��'d#�ws�w;<'�P�
��8�o����-�d�8��K������޽��������� .�/�ϘtTΆ1�Z���5Ң�,e����젎h ��>������(�p����F���zh��~t�i �"����������p�xU�����ml>DA`2�D0A��C��m�;���0ӯ��^كZ��W%��R����Z��OqOzZ�׿V�|�J\���Z���<�m�#�vK�?�N:8揎0kD�^�A*��!�%Q�?LN���{�1pN��.&� ��Y��j��,[L���B|��+S��Αu�d~y��1r,���z -	xdc��4L���H8�]�Ī(�&���k�m&�E�!K1���ذv�O���|?R�a\�x�l}jξ�;K�Xw�[�{�3툧�D�.?L5���������}���"����c*~j��r|C��E)9v����M�
����q��MmQ���[����!����ne-�������-��SAqea��站��<��ۙы�����P���4d\���_�ol<�y1Z�������b"�%]=�
وnƿ�K����x�Nf�u�~$�,3:���e�9�X:҄�{�J)��yC�z8�ͺ�K�XO�[=�^�������/2�;�:�D�1g��!Y��a�8<�j˿ՔM��Kxy��1m֋Ԋ����-���N%�'��S/�)������@�w�nǹA����sU��6L��6��~ԃ��m�/x��ۣ���@m�N��S���/U�����la,�'F1~5���nA�X����.Q�������{� �KA�U�sd��;�܅��@���xDM�q$�7o�*1��yᾛ�O��`bo��d�`s�I�ܥi�o���[��k{��]F7��,�g+&��?R�+���� ������� �A�X�a�7)&Ǯ,N���a5k�$<�6wu�q�3�3�����Vvz-�z��;�t�>���n�c�0ٴ��c'ԛ?�a�,��(�����G�tT�z�AB�ɸ���%L�'��R���%S���C�%�ǜ1�i�(���������6�����c��p����]@=>�Ÿ冲cE�T�Ie�7t�?(��0LEy���[#j��zN+k�K���[q'�MC(����?��������]�Y��Qx���S�j����<��p�梕9�f�� B� ���K���4.C� ؾ�	�2��{c&T^�{�kyaR(��'$]GW�)�)%Ȋ�C�d�`bY���c�$��}`�R,-��������Zv!?��^D/� ��-�r�ڣ���-��"���q���X|%j�.!H͂lzt��/je�o��400�����:$'GdU]ǯ�B��XS�:Z������"t�h�=��aqv��2�*x���3�Ti%�[��]
�z��UWn^^mfS�-֧��G;,WTT4m��;���S��sP����}D���
|���K�{_�s����X����2m��D��5�]B�)IѦU+c���l�B�U���	-%�G{J��}_�uݟ���u�;��:���<��x>�z��u�o�(v;쫌NH�s����A%0�x���)����t>Rń%0�B����	��������o�uvLo�����v@�����!b�]-�,9�6;����`��d�Js�n��k�u5%�e�3}W=fg��Jص�w*u���N�9�9�軿�x�@��� �k�,絳i�%VV�Y���=Qe#��0ծ�X���J�^�BG�|��ϯ�0�(ɛ]��>=1f�/0�d�V�G�gǕ�N��6Ɓ<V�}���p�,^�f��YM���Xcw�ga�Ի�=::t1Ci�j�y�cRX>:5զ�G����<�Hu���T	'D��8W�|sr$�Ư��bS$y"�P2���V,����f4<fG=�H
��-��m���T(ۄ݂#�����
K:ĚG<=g�'�V��a�6���� �F�s_x�['�wI�}m�8?�2^�+>`
��]�5t0嚖��sp ��_����%�q���j��N}�]O����0@o�h*,�9m^+�aA^��Gs'�� o߀�c�ܛ/\?Fȇ��o>YvZH������?��D��Z�����+ ��ڴ��BERI4�xP�)+�tù�9/���U�K����&�6ݭ3��d`݀E-?�@H�k�"������ةkiF�b�+��"�Q'�랞�=����d�[�(�[��U\�kT�ho?�}��}6�x�Q���?L��@���%aͿIMj}���p�����43.L��C�����>�h�-���RL'�i�����T�MӼ{�z]³E��5�v��2*
��@�)@̒��[X���֏�'y�F8�T��<8��=�)����hp�I��7
��]{n7�N�2�䊠#�`�bՇ|�,�5�k��lf�\���9�ۖ�sc=?��$-e4�H��e{����e6_
vj).��Df;�r:66�fo�lo��QtwEo�>���Gp	ƚ�i<���	�nEc[� ��a���S����7ÒKTE��xv�eَ�Z��
-�w�y���(���Lo�PZ�5�`����ɒ��%�-�#������-���c����J�d�'G������T`T��>o�u��I�Y�/?)cb��B;�VN�n���^��%=.�=�TC�����u�Bc
�w�D�.�������t	*A��PR��(=�;;M3�M��
����iV<x�߻���Y���	+�{,��2�϶���;l��k�.T�*��C/�tf2����8��[��GY�X��<rN�[�V �t�6�d4$xs�.�ݱs�\�85��м��DlĜ-X��ku��Ңb,}р����+�1���/O�����X^�M˗��}������~%U"�����8��!����[b��b�7w�ĐP�h�ƸNw����,sk���ak��s�-w����du1hg	0�$��)&En��W���Y�����]K�VaP��2�YЋ#�UL��<��l�p�O1��[���^�?Tpa�iRqHE���4+{���߇�]ad��]��O�����(0Eg��� �ws��?��H6��Ec�K���J�����p��.����.]��bq��e���w��X���{��b�
��S@Z�.r�o�n��m 8y�/ɍ?C�/ ����l*Bh��u�5�Sv����?/:GE$a���� ���JhT#,��]IQ�;�G���������-'U�`���c��PCׅ���d�'��/AF�
Y�F��\�q�3��v^�ӏ (g�
����^�zjR|{�Ý;=E��:=-~=�6�[6r�X�
�aAᩞ�t�;`K �G��g��*
�������n���ŏ��3��!-H�y.ͭ�\[:&���1�6����w�ӹٜɞbF���[�E��|��>1��g��5�L��Z�0��Gj&�4�P�N@�_Ϳ��?�s	�5�!����|�Zʳ��	G���O��Fv  f���R�^JII�u�V|�,�>,��������ʭ�u�A��LW����A��h)���?�}���ݗ;�N�����"\EY�����2�O��4Â�jT��$̑%_H���Ę+FK�o,����wqq�h�.�5GU��~�|�m��S��/�w���n苙L��~�?�ﵢ_�cX����j�`�#�S!�yE�#��1�>Ăn�h��U�ww����u��π[�r*�"�շ�a�]&�"�����Y������e�������o�
 =����Xה5XR\�h/��
'���: �R~�q����A3�D�L=וX�T
���_u6�N/�r�zޗ�q`� �yay%��)4��yHfN��+��"��n�$�jTѥ��M���4d����D�����2����n�l�6�>]��s� %
W�)-��w&����;g��ՍE�a�H��BP_/_�� )k� �n����������/SB`|�ܩF�R�1bDy�ݿ�鮫�o@�>˴�J�HW7�t�R��g���)���pv���^&IQ�J����̛�0���++W�֞=���T��YEĨ�8�P��٬s&Y�x%;� <��/\�1fk2�h>�ȹ�;S��*�>�:��~n�~nD���c�����*b�5�U�V\G���b�j��|�y�`fn^����J�y��aO��]��D�'�ݦ���(u���)0�
�F{��bf���\���D����R���K [�b��K��h�#��k�5Co��s����������؂�v�-^9̉����	����8���d/&��i��D	��Zc�;:hTvq)�`B���ue�����65�N�-�j���OƉ5)]޻��?���ij�'X4��'��F��a�����;C��w/�Rb���/G���>�ҳ����_1s^y=��9�ȁ�+��d�C8���qFs���h%����_Q����������4�6�<� E�@��K�ZOVc�̏R1����NRY�b^l8�H2f�Q� �fB�v�E0�]����F���G�	41Μ�*��~ z���{$i�y��Ɲ1E0�g�D�x�u
.+�IY@�rd��ځ�����gX��"��%+�Н9�ҍ��rr\i����(��kZ���p2z{��h�=X�$ɀ��[\��D�B�<<F4Y�b��r�P	��1v�6v�kLJ
����_䤝�M%�=P���cYN6��[3맅 SoB�-��8$d��6�����UQ�o��+i�GH�2 
���%2��e5i6�S�����[O�z�IQ��-��������F������Æ���y>$�Yc=��c�;��;d�tH��C��],OvI���~+�.o�`h
uE���4�'á,4���X����S�爋�ѷ�� /�F 0G���3�u��^|y㏠V�Y�Oi��4c�H)k�9^�;��|�͊�`f�- H6�RH��W� ��E�\��M��`|n��K��ɺ�?�I�5��O;�Dq�g��_[+{�P�54�l�}��ŵ5����mѶ�q		~$�*@�wV�!��j�!+�~��Ѱ�|v�6C'܆�����p�2CG��J�4Ao�ƽ-&�kƸ���u�?�)��w� �V�8�;s�n�#����@��M���ٕ�u@����#��i;w�,�&�ob�f�����$!��M�(V���֨)�j�ȥ{r��b�b�vh����ѫ��v�5�*��c�c  TA��L��Uű����"gZ��1^�/����ƣI���%C��<ͮ�ʏ����E���S5����B򅞙z��͇_�!w`��b�#�4y����B��AAAԨ'����9�f^:��@���h���_qS�Z�[�1N�1�AB�Qh���)=��
��W�}�Ġ������F������2胎ֻX!j 	�>�D��ִvW�e;���s�Fr���#p=Iʹ��X���߹w�0��ޗǩ���w���t����L͑UG\̦�����Ȫu�#@ʘ���`�:�
/�jnf&R�����ո�{����v�f9IP�Bө:�4s��]��z8��
,WA �[.|����diV���"�xkt�s�u� ���i�k8���ze�:	]/�(�K]Ĺ!��p�zna�Y<�ӌ�1A ��B���/�o311ѕ��
��ɿ�]8=� �w��c2HH�4�� ��}�A��Z�%,���:s�(�Ȋǭ����f��	�ˬ�]6x�h�����P@�J�h�g�1 �����.��$�HU���߯�����,8�����\V;9�͇�j@Q�0���BT��w���D�.Rq�lj(R��4��������p��{ ����k�����D�
:�96����#���&J2�4ﶶ��7*`��i>9�(�s�)`�&q&�r��+z5n�Z�n���o.�������=�kb��ps�&q8�W�8�����x�(�Bȭ��]�����U"R���;@�|G�ʇm���T���Xh8����U�!�X"�a�'%q�7��G�{�������s3-�C�Nz�����VJ'�����~�,emG���@*!A�ZE۬=F�LXqN:�Y��c!2HOD��c�&k��	������*��e����.>���	M,�G���+�fU��C��M]�j�N�>e��_�͉��0o��n�0ֈ2�ѥ��v�D�w^��؁�`��ڴl��z�SÔ1��.�4SS���ڬ��>�X�GK��@�ڵ��#>2����@�t�X��) > �m^]�����$�L�q� ;^?Sϸ��&�hk��bx���8�v�\�����	=��$ʋ�>�d8����$�R�FRJ.	|�a�:�ũ��:ߓb5��<�o�ϐ��@9���@�T�C�)��v�I�?r��7�9�{�m�sㅅ$��{��z�"�&Y�\E����_����G�N��Z��L�߹�tUq�#Mjj^�2�C�Ejr؜��.��zk��:�eO�MC4(���͟i
@̄bRq�&�.���&X�F���ن�q�xX4��g�#��bf�t���.֑7Z�)�쓔iɃ��Q%���saL� )b�^SPdl��4��U���
Lҏ��;�gW���W;k��]��C��f-5�R�Mox�ڪ*^�lsް��";b���ܢ�B�n�������*^�o@p����k�LP��^%%%R��>j�v`��&hR�CM�qE˹pP��4����2�ۚdj��E~*EjZ&14��Yg3������%oT�kIi-[�y��
�|������ϋ(���))$��E�ԧ��c_t	C?f��9���$Ji�&E/)Q
㻓�O���Xl�{a�ʹ +"I?V@������&�N4�|�O�.�A��@ ���IrR����D�^꤂A*� ���(^��T~X�|#D��:��L��rD�U%�`[)�$�0g�諽<R�a��`��M�������mF=���r;Ek*;�:ͦ9IBԀ$2=$���Ø��ν'�P�X�<}�zIp	��$��0��S7qyψ
�~�
��D� ���}XՈ�G���Z��{a�'��fVV~��НY�����(��e|M�nx�.t;��)X���@6�v���9K�Hp�J�{����J�U�:Ds���(/��̣�	w�o�־3�QThYm����GMR��#���Qdm��;	$�s���_(X�z�X3��dz[0B��Dm7���Q��H��}^��,P��od��"F�{�5C��@$C�(ap�}I� W�vJ�U��&�} �ۜe+c�7��P �H���Z��h\�1s�N��5�f����朱&r��/��*��Q]��JL��/~�>A��̇1 ����@w=;���$����a��:H�gz�P��߇Z���,�*�$+�ڈմ���)6,������D��O��'*v���A��N0�w��׺_� �K�`5�*-ޯ��o��l$כ�.���=��
U".}���}ٲeT�a8TUM}e����̮$�h�`D������;�UЉ��Ō>eZF-tl��G��OG5ͽ����.0>�z�J�#4��T��������1.6�K�Q'���a#O��ы�����tĳJLL����ğ/�K�sz� � ��}��M�v�����vf]��*yg�����1}�t��Km�<�(��A\��F��,-�H2���>}:�]�"���L{�ɾ�?���忘Qn�Ҹ��NH�Y���,�U��t�-����*5�E8��vw�:�?$�`�-+�DQ�B�⊁�!I�\��$�>�n�tޢīV�AT.$}�����??�|y}�`Ѩ NC���)�I%{��m�	�U{{8l K���o� .���b�G|�/vZPU�+&}�		��?��m%]K�9L�~R�b��� ���R�X�O����dT'�}��bi�+7������$��X�^H�Xk�,��H��R�V���M����������L�ъ�0,���^��U`J5����FL��R��Q�a=��N?���N�oO!0��� ����-@pr&}6Q�#vӣ�x`$uv�)k0���� Zؖd��d�H�<���ݔ@��Lğp-J/��B~;aR�q����+���I�oٜl��g�ja����ߔ���Gн�>qi�M}6$�?�;�Zj��1��\Q��k�9 �/I9s��&U�+�coM�fh��^d��Dl�����f��ڍi�g�4�E�4w��F0�����Ԍ_��T���L��8C�M2.˃FB�}�}����gb�ňTa1x����������5w�EH��R����\⴩��~'�Ay��Wz�&�d?Au�����ƴ�xP�x��:��iJ���������X��JJT6�F�fn%��/���؈�t�4�~|,\����ǊL���Γ�P��?��c�Y��5���;bb��s/����?]x9��_�:ijw�X�_�5_�d���>w+x��Hf�5B.!@�ҿ0[�d�
�ӓW�,�+�<�]�p�%(��;�f=)��~ɫ��`��/�Sy�ޯ �aA8�7IM�n	a��0�k�^]a�T�J��#��D@�	n�ձ8�G늆��NR�.#���,q�r\ϭ�s�";O���� ��k&��N�����a�+��,�d��e�Iu�qS�?���ڀ��Ɇ���g���%� �T�`�!�T.�:�n� l�4�-��е�
��OO�t�)�<��ĊV�Bq���F��f݉YDL��痗0s�ki�Ϡ��y9�8�`�6��no��|r����c'ô�n��u�q��2�eZ�H]��k���N���8��Zj�H��Aatd�*��;@���5�V����I^^+���R�{�	�Q�bt���Q	�V��� V����V������ټ������k+���������b�6������a���AT��LUTBBB�c�pq�4���%�J�T?<ʸ�B�+
A���k����$ \��o���:���0Y�?�1[Lv]��cݭ �q���A� �aʝ��0�@RaR��1IA�"��NX߇�0X3;��I׿�0f�5	�ϓ��%�	~���c��T�NY�c/�C���W��N�Ǯ@SW�����)O�h��hc�j)�=��Eʽ����z���6�Kk�T�|||�x�-K��+1</@.!�h:	�JCJU�"��E�f�� �8��m���40Q��7!���1��S�ͯo�cҔ<y���]M��U��Yk[*O.�~����m�M�Ci�&9��$b��xGK�2�B$%%�B�� �r:�(�� �3z_�eJ��yI�|�M�C���������m��L�Qe�6�Y%�i�&p�@�N�LP��V��)�)g��"J(��666�p����^	��YY�nkJ���
}x��%�n��C_�[3�jk�a������134}�?w�	ӝ�Į�n`����`�ПEC�<��gB������x:I�F�)%��Y8_Q�@:i�tŰ�����|.3��9�8��̙��A��NI���C�-�gε����4��r>��y������l,��w41}�7X�4�܄Gp�k����]�[�"�W`tj���!([A�
�(�������!DXwjCp��J;bF
�`�l��8�9����%��XW���^@���\0�!��߮�o�œZ��:����с�o�oT�w���a�A��ra��𾎩ƑA�
�D���9��3mjS�=��ȿ��%�⽚>>~?KP��31�mn�����Q N���4����t�Lue�﫱	92��*1c��/�k-'�}~��_1ƴt��-x���ԛO�?D��&8�O���}�<���wfH]�6x6�I���Ys�y���?�9�e�w��9�Al��
�~�2}ss=}'�%�U8?7{)�A��)�PM�I�,3|e{^�R��*�=�!�vG� d`��^�cv�J��G��5@������88��rAGڗck�z��;%77�ٲV�,^�`t�gA[��;�Fp�`�A7b����&�;U�8��Q%��+�y^"�T|�@ Չ��7/�Boo�I|��G|f�F�i)/>�Z/��FyѢ//�V�Jje��'����\����s�7��n�1�4�h�x�}xo�m�GS��N5���s�(�߼?kWj���_Υ��K��V���������{0;tމ-d�VMM�D����2a_o֦FDl��VR~��a�
��'JH���	_p�����X>�TZ s�.��j�����/@���.~��̋�7(ʌ!�0;�]0��Q�J%�F-�	l�r��O'��GGDDD�����׬�i^F��Y��kD�6���c�J��M�U����-�� �[-�l���~�%�s�a�wL^�C_�u�l=�R�ǡ'U�L��\-%%�uS��]^���گDj��o��/���vy��x�̦����ێ 򳅮�d�LO���?����?�f�Ut����"`A7�ď&��	P�FW�U�PA��FԦDGG_ś@D4���&8-��"3/������Ǥ�~C������VWWk28�w�Ύ�)N�!l���]
!~ڱ��aW��F��	�ˀ�&c4;D�D���r���: ���%�����fj���W=�]�f>���NJ&D�AQ����R��F	��nJ|�:wơ����������1Sz�\|i����Ҥ���ZX��ط������kl���7�䝊4�f��x���m�Dh���t��p4>��tl`һ�­�`���*��g��	����oa[�;b
Fi���;�؁�����}7H�f���=747�9�0ݮ/�x6ô����1�Th��76�X�8�Gs��W�7�F�Op�wE|�o�x'SL�
�Q�Gk����S͂�%l����L׏�H���+;L�XfƝ�����v��3�}��捕?b����w�����=uJ�~A��@���_9H��&��J<A�27�J~���ÞaA����`~�4y�3/`N�`��X5��s�wK�hs�H'���{�K��-[���Q��x��R;t�X95��;
�U2>�֌�H�
#�ќ�1��������ӛO:�wjm<�W�/}���}�zL�jE���@���mX�/õ�]� ��k0����O�'���~�8�!�_s�Q���,��<¢��A7��Iw�����Ԫ[r'�-�ކ(���*��}�� ���Z�:A���+�u��d��J$ɽ
!j�C��f�j���� 4��E�{��{���-�L�I/��DV�)ǒ�YS��z]��̭�����ӯ���ZB_"#�n�AaV�>�}H;��ЧJT�����1�a{>���������7���|Wt;�%�7���2���&ø��%f���Xd��7�`nU�3/�m��`Gg>=��Z8G~{�����8��5&�FQ+!��;�ϙ"��� ���#�bW���r2��Z��}Eh]��paz�#e�7"D�2�/HaR�C��D����xx<i��iџ�B~�HK?2o���/鉝Ɨ\���L�An<A10��0;^�*�DM�����c��z��_�zj���??a��X�j�偣>h&�f��t(����;�
��������c��=���K���?�`Dn���J�z3oTY�sM�qU��7c�����#���x�{<��������~/E��<�y�a��2�ߌ!���덄�ob�>�<��Q�^��<C2��Uy�&'Km6Ⱥ+�{���0������L���;�v=��<�g��������X��i�) ����,�ۆ�}���Bǰ�w=�Q�֫��L�?�1���$#}�\l�����������%�F���-Rъ�JFK�_[�hjy�nJ?mFY�|i^��g��1y+�m>Ǝoզ��LbQ'tT���9�p�|�ҥ�U�zv(HW�L��ȧjA2R'K������C�ŗ���=E�s?�!�L��ʑ,�ڳ:$a� zh2�/��̴����񫊊Jo�=p>�=���Te��s�pz�un=�~<P���&f ���>VF!$�0��Rt=۪|d��Y�vu��N|^����!�d�ôq��K�k������0r�r�U�����ʹ(z(��+����cl�lB��=�C�VHS��l\��n�Up
N�+�
;�V�L���o�	5����"�p��X�4���$�	�tU������8�7��/�����t^�G$����~9�N�'e��o��-5��WTTDm��p��"K"���+�m�8�8.�7�\�U�*B�41a�`�?��1o�<|�Bd���O��U�8l���
a���TЭ�yn���+���g��k_�R���*
���[w��zKuM%��w�pRY��p����ş���3{��b���Q�ZB��X�w�]�g���p.����
ȫ�OS��k)u�o���cN�ܒ������������W"`���= 2$EhBj��~�} �����CRR�H�
��Yqm��`~Z�W�Wo��	C���w_�	�LLZ���`���1����mƃ���'i���Z^�k^b�ׯ��6���OL��?2yȄD��KKz�LA�
�P�7<<m+z~�/cw���p�^|iJ{0n53zeS��UR$1[�7�Y�p�]=�cP�����h$)Ju�L�}�7����L�p�ߴ�=��V9��_۷��ֶ���&���NL���,!i���D��Lw6GG+�p�5H|�8���qG�6�rN��	jf��Joo0�O�>}�Qp ��ŇA�q�z�"P��a|�)�w�������z�H�0�b �7-gWH[� I���]64̰��3��z,g������K!V?�� l|�~�ky��P���٨i�t=a�;�U+���o��n�pd~z�!ز�>|ϵ#����3��&�L���Ejd�zR��TYY��9©u�X�ZVV�`�n{o�ZP�8�鱎�j��*�OE� �l,��p'��D���5@�}��+f6kFrU�띊3͊�-� \�.N�[%����5S�%���QaM#5V~��H��!B)�8�&��C���=Ht~́�WQ�V�፫���mx%�/A/X�@3���^[�g3o����@��PaY�������in�I�	�
j�cυ1��E�]�a�6???I3�Y��'))��5Vo�k&��F?s���"��/?�j2�SWV^�)q��_A���LK}/_�l8nk��U/e�oƨ�.I�|��v
}����UO��=z3�-8 (//U��E�d]�o�m[h��ۺ�W����E�����1!��6�9���.��E*Ʉ���|�i��O���5fziֿ�+
�z�h�u'�>%"�� ��B`4��+�������7�B��#��>�ٷA��B��=~3�|�զ�m4_,!�&��t��Gz8f]�M��׊u�5q���I�?�G�~ML�/f�\�~aYe劺�:�6nw�:��Dp�W�N�(m�\�]�����ש�О�ύ(l�ٝ�ĕ����X��s#�FF"T(z�������U!�� V��oEEH~�R�k�W�Z����N�M�S��f0�l@�wv^���i���ъT՟}����'<�V��Y���a����A��qw�w��L���i�'�|i/����D��(ni���vM�q�`t��%a4T��-_���9�%�K@��V��ǿ�BJ� ��ޓ���z3��@��ں�>#u��{����#�˛]^�|{w��DȞ��}��$>�$��FS�_��*Jݪߕ;7.=��a�acQ�!��e��N��V��J�d���_����E�~{�P6�HĪ�
]�EL�����}�B��$aQ����d�����\�(��}��gO8�`�pҹJssw"�,S�TQ!�׳�s�A�"��>ԇ�ǎ[{���I�+��5�-�K�Q���`g�`ׁ7p*�d�*�sڂPD2�љ���"�3������[�� ����*���ӕe�?��bs�ͧ��6���7�h\�������=���_Ǚ
v��Y�eL0��zV
��鞘U-�ĩ���v ݧ-Ÿ���3�k�㏽9����jD��<���@c��{�_:��Gl䩛��Ӝ���$��0NN�+��!�B���eT�'臏�c_2�O�Q4����Rs�_a�c�E���l�O~,��Ϝ��w⌋�#5�����Ok֮�{'���f��짮U�ߴ���r��l8���Y_�|�,���i>uqA��#�,��X!�f�:J��WPQ@<g��ʨ��Y���~!�!L��ǀ�B[��P6x={���T�6����(;g��6�Ź	�ш)P�Pc��?D}��j	�%#0bg|�wͅ$#���p�(㙄����P�aأ;��,�|�'�<פ*�ƘP��؝��M�qףd@]�/��[��2?5������I	/�:���A"A�H ���`a~
�\���.F�L�<��ŅL���Z�փ$i�&cpmP�U�`ۋ����q{e�*p��6�������ͽ���}[�SӢf��Gd7��T�2"�s��bY��)�w*�������ǻw���qI"����^o�)FP�ŋN_#��V[�!do��$�.���Y�1\����I�����an�����Ltx�|���!߂9ɕ�X��Sya�B0-��`���=�����G�y��%�.&rc�� 5�����SV�"=ommeNK��@j�����h-���֟w!e��Z!�"V]�Bd�m�vV�wuyc>n��a�K~x�ٴ�`� ,��[Lv�D=^�wW'��Y��	�*�ӹA��i� �ga!ݰb�%t���iҴ���foX���>4�"K�_I����c����>��a�t�����hT	�>��_)*��o}}=���@j�-��A���
~�)�����r�T�,e��ѽ��E�'6�!�~o�k�yl�`łL,Ȳsp�(�!�����/������xˇO��#+�Y�h�b���`*z�u����$2�ϔc@��0�˰Ot�Ǐ⨣D�{��F����0�@%uw�~���EI��h������u��={��̿'a:'H�Ѽ0̋[� M ��T94_�8�X?u���pU���o$:���3�X��������ZB?��,�?^�!��U�W{�#�<E)�һ6��AR��������b�4C���z�j�����}q8��`���à4�0��9-�ĵ��x,��H
�nC7�%��Z�<���L�ʆ�.ED��	�Z�ti޳R��LUgN�Ɲ�;���D�:uꯠ]Y#է1��.��1H%?6.������_-�����F�+��ԘFVYE���J٧O���rPA�-���x(0�P`����1��ѱ�P<SL�����
ڶ�� 
����`����Qc�8&������B�ۀ6	j�H���Y�;L�`6�2�;�G�ӱl��L�cӈO��g�����rr���@��J������ѩ�Q2ߛEm���)ժ!�5����@$w�L@\!�q�o����]��򮇿$�L�c-���0��;����wj���Ԭ�d����*!:������Bh�c�����R��̦;��o��ݰ���;���k���RS��?�*U��x�Ԃ��Ʈr
�)�,��1&�����28�ڷ��'�� ��7�R�0|�]�r�����&?�(�t�6{5>�f8:���^*���K[I�5 'O8�|��u�믉�%y���24]�<�(��3�u� ����� ���k1��ly*s�/���G꺈��q��s�����q֧�OY��>e}��������)vU'�_r�xt�u	����;˃�b�X�����mb��w���j�Z���j�Z���j�Z���j�Ok�}���q]5c%*9b�?߇�X-V��b�X-V��b�X-V��b�X-V��b����2�����o3/V��b�~�t؈���y��׺o�x��X-V��b�X-V��b�X-V��b�X-V��b�X-V�rk�C7yL��uڰ���5���8Y-V��b�X-V��b�X-V��
����w� �m��j�Z���j�Z����J<]HЉ/N�E&�m����+�;~�)��j�Z���j�Z���j�Z���j�Z���j��lї������~_½5��Ĺ�������c.Z��׿.����;��)jm������������������b��5�����>~��?|��Y�d��5 k@ր�Y�d��5����kzz���م��5��*�ږ�Kt|��k��<�f?��+ެ���!��.N��]k����94���[}�缸(�ߒ�����������Xqa卤���lO�iK�y�+)Ŕ�Y�+gP�}z���g�{���I:�mZ02�E����u�.��f%ۧ�E�GJ��&KO�5~�a��I����O��Jac�0�۞�O�^F򎰓Om�έ�GW��|v~.s��ۤ0���r��&!8��z��:���-EI����coO��9���c�.r�8E�����e�ů?Q-��x9�����E�F�=��>s��&^"�����cs�������:�\�����l��u���x�H[k��F�f�V/N؋VT�z����1��_���X�7��0/�͉3=חYԴ�2���D��X�����j�������lΪ<X��8r����6_��r戡ai��O��ZTӂ�lmm_�)��w��,�z��tS�y.����̝��q�ec�=OՌ�o��>?�����N|�t�����%��$�a:�t��ٸy��~����>7�_���HW7�k�� M�;ǂg;>�R�Т��7�ו��46����̭8y�^�/�%i�Iod�@~�-�W��E�5nc�M��$o�Rt+�u�l��i�A����jV��:g�K|9V$�m��� R?~l�L�.��/��;�� �o���F�;g6��-�ӧ�'>~�������
�m��)�[��L�2�~�&==]&\�A���'=!>�U���Gt���yڸ�٣�����׀p���Όq��J#:3�;���ڿ}!,�f�y�\'�VK?����t>�a��3�ڕ��W�mH�5��[J��Ţ���O~�ٕ�
[��G�pv
�	�͖z�t���$�ky������b��}ʀ�{��v�G:�6���_��^�{�d��B��7)�m^����f?E����k)�ms<�olf&R�(��I7۫�*��x]m|H����N�뺉6����]/^��Ñ��Φ���،tU�Kv������K�����2��.J�x������	�T�Ġf_�G�^�G�3�}ԙq�������\ⴹE��k��+3kA�]/�P�V��Z����@��>����^J�nW�|���xk�ۄ�YSa7�>}S+9+�E=7#�]��	U?�[��;�u�6��{�+2��c^����;�-řF��11��H��;��J��QHk^���3#ͩ�Hn�=̦�6���nq�|F��p
͵�6C_��9֥ɇW�t��ON���4�O�q��N����}��6����@S�j:v�����+��efw�E�B�#l-�Ͼt	F�i?M�����fI8�kz������4ڞ����NjKuixCo!t�����ʫ�Gw9$�e�?��Q���o�Ro�dKB&��o�O�N�iJ���q��)zy�O�>m�y��ѫ�=,��,}��k���V���A�Ӎ��w�5���� ���କ��=fݍ��sMlF|s�-1��T�6ǒ��.�9��!��_Djɒ%�[����t�4Z�^�8��у**ð��IfJ��;zG'���
>b�O�n}zbRүbbbt{��c�k��-GYK4,����N�h������`[�Ao�#a#777zNK�e�ԇ�6_?��;'Z5�|J�2�1�jp�2F8���Mv8�^ͻZ�k/Gyy���	w���������Gdm,��T|#1���mw��}��;&��{�;̓��T@֯2�%''��p�wg_,
1��IIK{�x#�������Z%SSS��Zm�jj�������V���ݹȴZZZ0�����t̳_$��d��d�}a���Z���=���L+�k��G���?�`r4G�� ��ɑ�k��çj�)���4!�6g����F��2������8{5�󄄄��`���c���읾5�ւ/\�~hܓ����C��D|S���O��*�}��mm>4�T�L�>yy~��V�ϴ���oLA}KS��IB��o��j��WY�h��t��u@'��`�l�!ضQAQqv,ѸP���pL,M4&ԧ_����w�;�LL�>|xmӁ���4��/���6iUf�ո/ق/�L�U��_�:�[Z�,��u��o٧j����S
���1j�qۺ��Y�&��e�5�i� �<i�q���w��i�O��b��;�C�u��I��*�>*y>]k2�u�BBf��_}nx�lYm[[��sק�%��n��O���+�׺�u�#�`�wZ��y$����kv�f��#_36wd���I�ګOO�A��m�l���	ǵ/5��'w�^ �P�J_ۤO���)����͈�^AW�K�b&G?.&�g����C��S���x�Og��K��<���C�}��˫���W�g�ߢ��i��>�笞>}6I�k��t���>�L�������'���t�G�11��\h5>Y���m:��^%�c�jI{��:�[%&�2���c��;�7P�w���i�3�:~��#bbr���{
bm'�sN��q�
l-��ˑ8�86�Sth	�s]�p.�������e��b^F��}�˛��5�<	��Z%[�P�����G�6��}���c��=��r�Z�M�Kݥ@Z����-��
F<I�*�5�'�j���0[	�I��I��0���t+L��=��w���q{�/<�Y�jn��I������P�\��g��ٔ�ՠ�穕kV��r�2{����I�^�,�֞n��F�[��3�E�t5�Z�ͼ���N��/>�{t
�J�)����Ŷ��������I��2��O�4����Z�Lw�I_�*��76f�;�:�a��(�zy[��#T�g��~�v���h,��S�V��{ԇ�N>�7Շf���wG�Z�r��_cl��,CD�#��	�F���5���(\|v0o$�#aw�bq �.��!ɛ���tw�O���m0���E���������ޙ�gާtG���+V��EŖ�rӲ
��ތ����:��=5���d�nS��&]5�V���j�=�9p�[�-�� ��vg�x�4���ڷ�@iK	}�߱x��d/�#�3��ʄ�l���"�C��Go��JKJJ6����4�s�5������XT�����bZ,RŜ��=u���+��G>�~ASfC� Z��ԔU���8�9�~�T`+�Z�B��L����RP�ڕ�J{��N3�e<0bG�ӧ}��̒փ�'���"�B1k��Տ���#����&�<5�q~}z�e�0s^w��������&ؖs)g�;*��3�g��3��M�}];�ӳ)h�䞨N���>ڻ�%,bn�pB�"�Bސ͈�ğ����tv�ff%�)*�g%[�m_�#D�M���i�Spnɽ0/zc1�j8y�XV	O�X|�<RͰ��v0�(s�+��C���5�n������ӛb���%�ҵGN����s��@`��-�0l���ƭ�%R*����g�t�C��D&����m�>�e��צ�2�&6u��W��O��.�4|���qd���>�6�~7��\�S�3����Z�"�����|���ۧJ��hv穔<�1�?o��$�:�ڹ����4
�x���7G��i&��g��ݛtɮϖ=��=E�;���05��@6�K�E���RD�q6۲c� ��Y:���R�w�?���t����8k׭=y���᣷#�������G�f�R�j~���H���HM�R{�ܾ�,}�cǜ��c��}-�iv�q����ܻD���u��n=��uqo�^���)~vN(�b.-w��rI+��Wzߑ���3�x���k
��͢u.��!��^v�ҥK��@����ގ����T��}=�I�#�;'F}j~����?��y7(�m�ל��_k71���/l!���wH�]��լ�<=���	�GT���~���#G�d	)e�nDRb�z��j�H�w?�.�l�I���l?��m�[���I�=Rк�"�F&3�u\Nh ���'`�U�/0ia�����h�mi�#�z=�K7�6h�r�$ׇy��uh {�}�gdZ��^fg|f������L��������Sͭ�v�I���p�Z{����vC@�O�vdXrqH �ؒN
`:���5�96ԉ����2�ҮN��]688(Dּ�{<W~mSW�3׶ Ǐ`�߷MeΦk�EM|��l�ӧ�rH���A�lܴi��yĊT8>3���m-j*�N�4�yl#_Tn0�_KQѺ1����X�#a�h��5)j+��{�Њ����8��B�����QP��{��ro�����0���x�&�N%���,�	mN�8�m77�Y.�a����/7�>���Y�V��^�#�[,�}PpT��6��;�?�U��6��bY3{?b��o�Y�(�����Wi @�q�Y�,��m83p�þ\���^z�;D.e��*��rX{��ޞ�qg�����}��:�~\ץ�w�����-�)�-|uv�[@��\z\��=L&��N�Љ��p�`L�m�1���g�,��mrt��og�8�,G�v�C��ԏ����P�:�d�J���ه��0m+�z}�]E&��@8��-a�������W�tF�k�񖜣�v����g�� * Cq��h�#Ge�^��-��Ϯ!+=��P�U`P�<� P��y��-���v��(V-H&9��xl�Uԉ]]ghf����.h�;w<�`oГ-&��q���I���n�n����壷�{����	.y:M�}�����mHWϞ=7�i���P�Fi%7w�2��7&/î8�h�<�S~9�)���q׮]�N~��=����WWz����b:�~�:~�*t���ם&���2X0M1|��X�x����L�r]�&�Ӣf���˗V-��o�s~���Gh|�nP[���S�� #�U�uNՂ��ګ*F��N�w�0O����s39��,ԙ����\���^�=o��YM�`��d��:��w���#��i ��Ig%�=�+�	L�՘:�@ϔwd�ݧ�����:��E��&}D��':����6�17�-U��)�5ܰ�w��=�Ik��:�+��}����������4��֮mAR�^Г����:+��ڈsv�7�lG5���s8��ҲG�G x������CJ�1�I{�-�;2#^4V�j���B��%�nKV+������~P���W�ק[-�T�Y���wc�}̫+�L�Xԏޞ�����N�r=��{�����{�b��6�Ӌ�a��:0��G���.�B���엫�B�Adk4yӬ�/.d_>1=� ��Zq��/s���O��TVL��	!�pPf�h���]����v��7r���P�tn�ZH8�k����w[�;+�u��-�6+@�uD@!�G�*��[�K�>���T<�#D�q���'�g�߾{��,�\K��ಮ�.��x5�u���ޚS�cgA� 3ܴ�|E���8rğ����>7�����0'���m}zĴY�RG��=!�i2��Q��I��;.��M���z���ɲ.{kRN[Ը?�wf�]$t��:�� �����vefL̄)��~�4�Kwdl;Ƣ����(�s�:��
�6L8��?��q�Omm��sC��,��w�c{�/$ކ_5��ޖ�)5pq(��rF[�b�<�!D�!*��fE��A0+�E�����ή��0+��5���ka~h��bX�������e�`��l��+?do�9(QQ��n�����q�Ӟ��ys�9�6|2!�k[����)s�ɷ��S�n��W���]��OI�yl���M��ʙ����e�v�M����v�����y"�o�)о�J`z�~�+��E�ne�k�Lм�)�v�����b��3?��3��"ϝ�3n޼iL�^/ϦF�[�j��"sh�>���.����wM�\z?:2�����~k��&Єג;�������	���8P�������i�b�6O�^{{�� ��S.����ۧ���N,�?��i��D��4���v��?ƺ�٥sz?0j�-���r�~�����]�~wO��~k��|u�y*���>m�zfkZU_9m}_�z�ӟ\S#���}�L�uS`��C��K����t
�O���+'>8�[}��B����}4�F���^�c09�EN�ܪ|ߖ�{䕹��.u�G���I���{��3�%6�w�Kk9�T���^_���������{:��������^<=|�4]���ze��iͥŮ�5�K��ܖ+����~��݋�A��N�;'��ʾ�ǖoy�k��)qB���S�
~\�H#�_�n���}3�No�������}U�+-qu᪟u���]�����c��9���e��ү���z]I?W^���d�9`�;�H��v��f`�ڟ���J���?�_�SjYn)�(OW?�uN	M PK   ��!Y���� =< /   images/e0d827a2-ee8a-45f1-850c-b31b1c4188d2.png��;�q�>N
��D�JQ)��J*��Uʾd��*�,B��}���m�Q����[�1f�>�瞞�9������s��c���u]�u��u��G��<\"\,,,<z��<aa92��������q����3�^��/������o���"���a��lb�<�{����������K9gW�g�^�yz;fP5EXXΰ�ݹe��D|%6���m���Z�}��G�|	0>wW���^핟2R����d��6��ń6���7��h����l�j����8Qe嬆�y���'�%*�����D� ߭C�o�+��X�n���ʦ�6�3��G&����y߫z��|��`��@�_���in�fJFʀxYn��Ti3��T{R��9�?�0�Pz�i]�����+�_����{�z������c���S�V���f���R��+��^������mv���ž���/�����'tߧ��̋�%��� �������'��ԭ�ΐ��S�����=���� ��݈���Yo�����'*c��}6c��jiՋ[�<�DՏ�&oR�����W����WKw�������m�a�L���w/��7�Y�g{{�n�핯0�&P�X�I���EG������7�A�b���Y~�a?^2B�Ʈ�������W�=P�^�8/��J*����<�^6������#��A�N).�=�H�{�կ����c4z��ڀ{f1�p��{M=��S=^�����V�R'�R糹�.'� �� ����D�K�m	�Ʒ�㕦�Q3�R��X����0��?g�����˩x�X�K�a�y5��W8�B���m'��\�O��/��ʜ�Μ��ʰƒ|��Q6(������2�I����T�Z&3��@(R�j�M�]9��)�]���I5���!�%�����s���y9U�����'�{���zd|9�33^� ��D��?��5��f5j�Ʈ]��sl�e���f�.ltXP����s��Y�<��V���p�.P=oq]�n4�¥�.g#Oڧ���/y*6X��:�G)�z�^?)ӷ�ꩉ����zmq����瘉:���R*Xo\ߔ{��[�Ю�]>N"%S߀��
��;��|H4�=�_U�z��Yy���_��S�������Dr�܃µ��4��k�s�Q�����=�'���/2WU�f��sv��!�m�'���׷Zײܠ����&K%�~6O"�4�_Ihv�>s�]�ڟ���e�0������wp�k����}C�"��r��O���tτ���5o�+ұyݮ��,�Ʀ���s�l!���)CS*=�2�ai�4)�u����G+�~"�����.K��"�B��Q]�Ư��*:v$fj-�fv��M��F�#�;ČۣzM��vr�L�z�zYV��p���㶃��Xâ+���ޘ�Rw%�y^øl"������M��60@��-߬��p�|�i�2�Cc�hl�D�I�z��yrz`� ����ُ�VpnY���`a���m����i 4�⥒��7ɢ�T{b<�/ʈ�V!�r��U��w"����$+5(�Ь��`�g��7Y��b��zJ�{l�GnEST�Y�^b��Z��㡧��-L��i��H�+���%�	�bX5���Н��\�����E��������w�UdUQ�a�4���9�����Jܢ��,������<e;��ARO|�-#\	忻>^�5�h�kC�+�%?~C5@z�P�n&ن��7���Q�{������}������H'#�I��`���<�_t�E1���?�Lҳ��H�S��N]��r�xy%���� �q�
p��I<vFU���=���{� �������L����3�~,D�w;�F@�ս��5gI|?���1��%�ee�����c!����]���+���	_$,�{�\�R�*	�mL,Shܯ��?��������y!�jy
:$`˷�ؠ�1���s.QI�=�.��r$w�'k��/1R�O�&�/��㱣k���]�����3���^���&�*c|t����ᯙv��!f��ɳA��-����f�F*1Sj\/f��Q���R����|��ti{t�pN�O�|����2���/t,y���(�� ��#�+�6��O궖��х��X/�N/�_��9��P/+;�ڤjon�M&e��,3��B� ��\G���8�0'��N��k^uN%������f��[�@�|4���l2�FY�����BK�����
�H([��&c�,~oB�m��׉'k�}�(,�1��CG��~Br�m�'��{�}����.���<i%���١P�0�a���^�#ğ�X6�7G�E:ݱՒ3查p����}��9�:��U����e--�C�VQ[<�;�+��ؔ��@�Ϫ��7ೲ��O�$�4s>v�&��pq"��Z�-�}���~�lȣD���*h����ZWR۶�|D���ܫH�]�j=�Y�m	`�)�p1����S������ɷB��F�N��%�M5P�}|��i�W=ո���0��j�Ҏ3�0f��Fv��=Ī�v�O�_
MA��:�އK�מ�$?=T��WԳ�,z>�0~��`ԂB��W�� ��e�%6^`"����əY��D��	Yl�0� 5�\V'���T?��e'�5W�_�էP��i��y^r
�$�j���\���{6����6QA�7�������)�:.�
�㽟h=l�Zy�ܱ������P�5�ϸ�͆����L�ᐾ���(���,um[�9�ia�I���ä��q�o�Ҽ��=ꩆ�1/5�4Nԍ�������۰dl�`�����d�����@B�gd�V�q�������` ����tc}W�.:�1���L�-,��eg�>5r�dHnJ��]z��׬���z�kBc�K�����58��A=_~+nnq��!f�����@� � LC��-a��s�Tĳ��ї� �.g��d	�V<�1�wC�t>'5��٭�+�Ԫ���D�x�ms2cOJ2c�w�7���c�x���,������;��t����?ʲ��mu[���q�f���[WO��;f�qӏ�7\��>N����@��D�) ML�7��m�M�:Gb�C����w�/�p�θ*���@���t�&A~�9�	%�b"��1My?Q��A���[�;��"�R|�jE�W�\�BU7�B��A_�@ދ'�xLO����{s)+j\α+Ѻ[�ق���h�Bcӹ��T�u؅�TB�ހ�8�5?p��~�&�@x���p���4Bx4��&>����Fw�\������r� w8��-�_ڜ��P�J��[�@[D��z����?!bq����u�k|�y��x�\�iwH�8��!Fb��)���N�x~l��!�0���B�c��j����9���:QF���Y�^�fh����B��z#�b�hʩ�`��1�!h-�3��d'Bt��2a���K��d����?��%��x�-qk̪�N���,۫���ri��	K��n@��pp�ǚC�h��qV;KD�2Q�U��VdT(�5����a����������^��^U;�V�5�Ѵzۻ��,�'�Y��^.fĩ�u��mm͈�(���V�~�6����ɀb�7��}�r�_/'����q���'�*<ѣ�bѤ��a�<왖�-���Z�j��;h� sWJ��M���h�A�R.w옵� �SRLй&w-jB��7k\�<i6�gy�>7:w0����]��>�D��˖ I8��&Joa������ja�p:e`1��40T�#zc�w�U��l0���O1}O��K*p�7ݚݾ�W5��$%%�O���Y����s?V�z�S�8�g�'{��YU���ҊS �rJ��Þm@�[�p/���vWW;�2�Y������'>U�p@򔘇�k�aQ=Ȥ+^���A����R�7}���>���n�|�̑9��)�/��1��k62���[�sy��ľ#c;��� A$���o����w�o��~�ہ&\J�f����5��/n��Z]�zj�w�f�Ĵ��N��wk�����y/u�F��yC����4l;��!��__�'�f:�>����0�.^�'�.yYmE�̢sP)�\�C�oJWV+^�#6��V�<\��]*��\�S7�,��$E&��Qq
�:��uD ���R4��l��O�f˭���ya���hh>��}�g!9�`%���2���j#-�4��m_	����l<م�3i1�ta���53�#�\��Zy�R��ȆV���Q��Me����_[ZЗ����SYx ��n�yD��y�#���1�aK9vܥ�7�@PS:WQq�>O�R���;�|R���Uj�w��cC"��:�Ȫ��
��j�%�xu��SA�)��ۯY��Ǹ��.s���c<�ۭo-���]�_�ҷ���U@Ȉ�v��٫cKhrԋ�׋ ����m4�li)�r >X�u��2v���e��*e��l2}���{�E��}Y:������vO Q�,��" �D�
n��u�E��-b]2�?a����
f�]�k�4G_�b�S
���d�
��@��>�3	�J�lr���3&䲇m�����	��-��_W��_����e���q��ۭ�t�g�or��>�}�߰\Y��8�<����2���7�� �b�t�拫�K!�%�����b��?"qd��?��KS3)ϴ�$�����4W��X.d��&�[����溙 �+��
���1B��B�%�v���wB��ק�I�с�h*�\,�9v�9S���k/�h�$ۭ�vW���Ѷ1 <�QP�hY�۟��!
	b��Aމ3�g�y�Y���B��uE��8�4יm��H�ȰK����B'�Y�8c�wjR
c{x=��HY��i�RUC�Kr�G��'1�ۃ��yƤ���3�A�y;���>��H��ބ4S@�u���n�f̳����#�<�>e,<i�����[�~_9Ӱ��$K��e��@��!V=�'�c
��eۺ/�{*c)g����<o�ċ��g�]�P6�e
Z)/���l����8[�V�������:�}����u���n[y���Ҽ��}��6�M��
P_�J�����ӥH�F�֡��;e$<�jbn�:�lw�<@��I0�F��n`tU��P���uxq}�"ҼT_oݙ �����׼Q�$gV2����ɏ�Y�qO{�g�p� �F��}r
��~J���Rs���e�� ������lN��'�B�!@��v�3����u�O�P9��,7lJ����!l���ѣ�_��Ug˷^�=�?9���w�З��^Q!+_�����[ BZ¿�G�c����4�}��+�w�4�G�k������ڂ�ar���>Q0�h �PiY(�z$*�����{��[��U�H|S����{�#!9mb�����p����#e>)��oy��(�k_aVB�B}:a�3{���G�����z���=	�����t"z��aRͅϺN���X��3��!^|��9dl��䲩to�|"��Zm`�R^����q�՝���>#��2r4�炯��P��N�x����1����*å��5ס����y�-��'z]����F��\����e����gOQW��iIr�7�(>2���2څ}y�1q.dHV�99��\ZL/��Fwy+b�a+�Ϧ��]"4ҟb���$�X�$��ӯ��, $��I�a��ec(�w�G{���t{���yB3+p�$���7@�e�N��Фyf�U��~�Y0x^�D���� ��k}�I+��O�u�����  �U~��G@F�����Ә�$���Gܣ0	���}���Ʃ�7�yh��y����i��e�=����QI9�iu'��}=f�e5��&��D�ᗩwc7���a2��H��vdy��Od�ǀ�����3g�HeN�x���%�ҭ6�u�q������)�{d�Td�MށI��A�Rɖ���ٺR$/��/�Cl��< /��D��E>�6�Z(腊��\lD�X��;�6�{����V�k9>�6�'a�3��{���G�v�װ�K7)���m� e�gt��|�j���H�>�$r��^�=4��QM����D�ϱ ��^QA�wr����-b�ng�Y;�|��"\%��n��VB�ӓ���1�mad`D����vt��9@6x��(%�d>��ᦎ��XH��`��U��j�����kМ�H<��1��������������ػV���l�٬�~ {��)rً���������k@�[�o����J�����]:��XY�� �f=���zajȬ�sV3K@�Z`�m�F�H��3��{�K�;+�J.m0��r"`�L�{��u*"�|�^�>/e���B�q� id������;��S���W�fן�ǄVԘ�k�î�;"�*:%�}�ׅ9*3OW�T��dȐ���4��D�HB��ߑ,F�0/78ꭶ�����
o�#:Y�P�F^����5W ���+�ɧ|�j-{�(�_�k�(m����3�{9���Q*�S�Gr��k�E�><9��\&Ω�����C�)�#cadܓ�mǀd1'�G��G�PCf���%G�y���M��~l^��[��>�C�B5��~래��]��ت��.�EѼ4Eӡ'1_8	��1w	vWߥ�������}\`���I���	��;�2<\V71�y�qg+����c���"�hX�{����.`#�K��	Qw�udO��۴,���Å?ŗ*�=�1+�X��e~eliU#�C�5�����⇗���5RZ�6�Yo��Щ+1e,1M���3r#�N�H_���0�[7JJ���'�ڔ��/���I�"_���=dv�& l�>���	���qzo��l�A�������EZ�{�7D�xJ�]o��P�������iGz�?*0����Z������}CC�!�#,y���?Eg[�x��
--���_)7z�����>�9�2;�u�������k�jAV�1e����ƴ�o`?����9�a��8���8��^��˽�ܽ��W]j����/���f�&D�X���,je_���4�|'���'���v��(d+�'��z�z�G������yO��w[G!����2hHyOI�-f�?��GtJ@�9���s�+�#y;P/\��~��	`� ]\���{Hwѣ�4 �y
��gf��p��3g�� ��P�ɘ��'E�nk$�*n��[��ޔ?;~+?�z?e&�ScW�>�`>�/HIG.���[�?��N�O�b7ԙ	9
$�WFz��+W8 �����/��}ّ��-ٵ�Y�����rS��*�9d�:���~��~]�-k�Vs������3�qv�(���Y�IH玎�+���9�\F!�Xڐc^��1���h�|���sZ�����u�{����� {����e/��:0+>!�k�P��O��6�ߔ��Ȁ�T����B>.g��	 ���
hKW8��c�Ԙ��� Gc+<�j+c���|���d'�ۑ���9�b��5��'f�̬�z�	�>S{�9JvڟT9��^NK�g�㪨����ql����>�D��p�l�j�}Ms#7��p�OY��	���	K������C��0�r�ئE�/7��/��P�{aZ����Y�,,��^Kh�/�;p�6R˯T;�Tn$��=�E�$�t���V8��j��ݐ����a��௜q����yj���:җ���B��+^ ] =wb�D�.(�ޣ�Q��"Kd��I�)�Q��c+;�L��j��ӈ	��ss���J���������P��c0�8avq�S]���-_?(��p�Lk��K�qw'�S���^�4!SN;v"��=�ۋ�+J�>v*̶Ԇ/�Ҋ��,�i�6��H�}^�1eP�ϳ�@�^c���}k�}������Y�3\g�n �D�נ�����!meDlf�I�X�Y_p��� {V�������	{s`?�H[���^��;1��'�~}[����]���VV?SN)o�%�f�:�+ec��QE��tǄ�WO������b�V���h ��?����i���l]��G`boi D� 5��rA���o#0�5�֕��|�$"u�yl���Ybg΋p�`
{��z�p�����YW�.zv`!����Xn�1-[-����SJ�t�Q%(�f�ǟ˛uo��W�b�.��2$U�FKI^HNc��&w~b
�䖝�y5zR�3.V|��_�}�ȝ����S1;�?�B^[�𩱜apR�.�[�E
����r��k|�q��omC�P.��qquM:?�(���3"�*�GCkv0��IIʰպ��4�+�ܲ_'�]�IVV�Qn\��j�q��B]�.#893Ա�7�M����ߊ�:ۄR���1���&��B��z>��`�D%E�o�ŗ���l�}H����l�{����{�4
OX)��'蕕�Y��j��ٕ�]��,v�|�H��Ɂi�b�WRd��w��m.��t�������t�/�f���x;���0Y��&L�).rKX*X�Ȗ**���`�<��'m��\��\<u$+��<���y�I3U�B�c�TdݸА�-��[g���?::��xtD
>a�;���3:4|�$�e�_���8Q��E�e��E����Vno:�rc��r��ѷ=����S`k����P�`S��=�[b¬�C��϶EʤyP4���Za��<�s=� ��Ei��^%	!�E�7vDy�(>���絶����J�������Wx$,T�_()���r'���r�$�XS`U����O�X���d֧֌
{��}:�kɼ{���л2d��y��R�ݡ&eU��YƯE�W���+�Q;
w���@�g��3�q�+��.n{AU�"CE�%�JS�B-8���uv��7��~����uՀ�z�%n�̪B6s��\�zU��hgi������̢֫/s^�(7JP�����V��xg�k=�;ʹ�!|�i��-�&��^[�W��P1v!!�lJMSS�(;�6,�l�n��y���2s��PWuÏ2R�#���0H��r�uV:۫%[h��,��F/���M�W���Z�g\��ζpN\dբ����OL����	��Q�"T��S꾏e���D�	�Ks\_�#m�(^<��~�l�K����[B�8�հ������)E��W��Ɯq	u)Y�7���튨�\ ����b��K��ڞ.�О�|�����V^��4��^��w|��D��x����q��y�e� O�@Om.�~s�	1+4�1R����>�8p�����8u�\m��5@Jf׶�
+�Bpk�k��j�d��z�1�Kh�$.�&�n��?���ޒ޷t4�\>e�Ůe�.K���㦝E���{��M�?h�ǭ��X��v�z.���T������r���*�?�x"�7�c��[L�@����43##��V�_�R��;�	crߣ�]7I'���Cg���,�+.-�)	 3���T�ZN$v)0�4��P����`�h�'ʤ���4���9��&FH~�T�3��[X��3*|�7z���S{�N��y;�����t"�v��u���~��v�}�04 ɣ�;�^,}*�E=;.�b�댺����9�p`�$�"��lܴԡ�?Ѽ!����,�ux�ޒ�����e�J�A_���j�ֽ�v�&�O�4̦X���{�1�L5̖�U���W�0X}���[z�T��f5;��G���������0͘����%���s~z}�������!���*_�4�����f�#h�m��l^a�)Аn{����Ç�vHc����7f�WԀ	���[3�p�[&��	�LHk�����:�^�8�p��������-a��Kl���n �zo�q�4�my����=�o
"�wJ$��W��]p 0���V�I�*��y�����H�aV�vtA��>�&.�{�D(���@����Wn��ڐ�"�	��L�����8ɻ��ww�wzƼ���t`}�)���1I]��ǂ(u����Top�ʊk�%���WS��YY����V�'z��G�/�5�.���Qk�-�+*������;�Ǔ��-���;�:��T�~��)�.�I>�?�\��ؼ�0Ra�K�y�͐���;�ߟ��!9HAM:q�軮Y��؎O�в^����EKU�Ը��G�b�R��Y�Ԕ�}��٭��M��9���ɞ��"�������� 1�;�~�U��ɿJ*�G6nߪ�� :��-�n��\��V��;����wa�I6lu6�t�����`jo��常�=��ϩ��O��G�;���M�MT.f-S_�ON�Mwĩ�L�~E�/]a1�j@lR	pd�Y��B����J�6�������8����M�T__����mf����KUާʼ���@�̪2��Xp-ݸ�&:���1d�$Q����o��d��߾�?�O$�}�����[��3���Z��#,����n�Ľ�&��6�30�`|�f�S���Dy뾥w��O�1�k�⦤��nۺ/�K��K��n�'X���@��h"9K,8�J������"�)��S�X\>������
t%CL�
Q���Q�F���(� 1Z�F�(�
����e��y�dr��l�`�%�����n�QD�~�j��s��-Y5>��a��-��@p��e��!��U���}!�����MS��k啄�WA�4[�,,�y���n�/���N��~���*JI�KH�^pj��EB�*��[�Ӽ�eJ��#�%~G�hT�������
�A!sⴏ��`�l�O��#���(M*��o%H�6O�s���O��j�9��ezFG��#1r�x���f��>�����y�	�7-:�5ώ7�/��e&�ZB����������q���oB��w@C&m�b��^B	R!���{�V�y�1B�>�̂�ȹۻEʊ׿���+���N����b#���'�NL���
Gi�8:������Fh(�by��5�:������t�[��^`��wf��_֠P2 �/S'��ZxC�d�� E�"���<wB=S����~;�����}�}ʴ6|�-!��1Y"��J���^T\�$�Y'����)Q�������f��૒�����WUU:��p`��9(�|�Ǐt��UG���1��v޻��'��[�EqS�!�V��6�eL��rxAc㏞C7���v6Q�2Ƀ-��ս������`��R�Z��5�By]���gw�K���&��84�a��q�J �tBmg���^ԕ�¥`׻��_��>�P��^�\���G]-7gq����ǖ�7MzKΰv6S6⋽�p�h�~�(�GG��҂��J�Jy?U&�'�0�
\����d:/�:��5�H���Ǖ��^3�x^��ׇ��,hf�ŗ~_a\^�'��m�|�>)� I�q�T�~�����'���|x��{hZq�o��B���|���B� �i�a�rj���ؽ��".���Ѿ�A���Fqa��J�f��b9���j��.��u�dw��8� H����b�L��Ë;Ik�B |�;��Ã��l�q��f��B�+��= ��T��Cr(��5!-3sp�yS��7IϨ�('����J�$��_�b�E�0;H�[J����0��E�0;h�)
(#1*`�.��\}>�@�D�Y���mY�k֚R۲�v9�f�l���
˜	n����/���Q����iTj�ЂѲ`�+0I!�G�&�n��i�̾�+3隡�3HL�H�V^h�T��5��ڌ�M`���h�+�N]�RdcQ���6lW7ZE�t�:\�ҝ����onn�+<�t���	����fa|.�t��W[�hC�࣢ʕ*�O���s۵��g�/7\ t}�Bk]{�+]�0�x���J���^Û�a����vA|B��%�+#�2
*ҫ�I_�oG��Ȫ>�i�x��\�Q1m�Ob�ø��S�·v���ӊ$s�l~��S���b9�0��b=ZP*;�F�n�lw���ӈah�w�@�n��V/^�1�f/��}����3�˶7Q��J&�H�؀Ęh�r#�3;�%���cso5Ap�204Y5�Q1�6�]����
 �t�Iy�m��Y����=eՕx��Y��_ѯ�W����_{L��ቓ�D���������gWk�cÓ����A��rV�����X���6�u
���� �F�l�+�t��yw^��o�r�X�}��I6�� 1����\'9�ш�o���ؼՎ����	��נ��l�\5>�n�q͡�!$����������/ך�o7�?�h�$�<��qX����p�g��M�X��#�����f���T���v��Ym7}�`��Ri�L��潾e��:*��0tA'�ٓ@�)P]��_`%�Y�,a@W��D��P(�'��Y�6��n�1�`���&�E���D��vκ���ф2���q���'���s��%���l���Es��xY�����:Q��gk�78S���}����	�(���z���wố�6����u����6���f�����e��M�uݿ�\�Z�H3Y�� ,����evv�����q�T~�h�k�$qx��7ln�q����`�g�>o
�&Q�9)s����b@I�A��!3�j�ǔP������<պ	\�jN��d| �/MQ�T����^W�0Q8�Ygkf��T�w����4��Bh����ݭ�y�Эr9q��YL�~*"+��k?\X7�w��Q��|���	�w,ﱅ�V�����Y���|n�j����L�OW�ԪC�al1+����)��<����fP�	��w���'�W���Q���bL�,B6\���G`lŇ� ����6ʥы�o&:mi3�s�Ԏ^�m�Z�z��O��%~�}����m�IN;W����ݱ���oE4|~�lUN�Q��B��`���Y��=O���>��i����]�]!���r*-+���CۉN% ����^���{8j3,�UT�Nଯ�zyo��n�������[*W��A��:��Z��_y�C�A�_�H�#6{de��M>#蛨���6��h&��\�~Fj{��*ʬ�����x���R���:|byOL�/o��6�VJ��%HǺ�z\b��Ϥ���[ٻ#`tF���\��)P綢~��`��T���W�k=���0l��h���!���i�O�҂���1���f���l��B06Q5���	{\�&�qJt�C���~Vòݗ�WJfv�8�<.M���Ѝ�7���S�m����������+��?q�@n�^����&���M�m>�/k�&�,!HR���V��� �cR��`�T��������:��~Fԅ~|�ll���u�'����4���켵�y�Hs%bpj�c��*f+�����d���Bm�m>���ʠ��{lڻ�ަ����'*ފ����u���n�;�T3���n�舳�t�P���U&z���F�p=�:_��g�X��7
��o���{�+��'��qu�5y�7K��YMmh4��[��g��m�ThH�P��8.ַ���%+��K�����M2Z�Z�m=\�'�V(5�܉C�ʱWboo� �+r_ق���V��O6�����t��:��rϖmw��N���?�n���;�H���p�%��U��~�$#��H��Ęk�!{�b$*�8�G~f���W�V|Y@�Uɗ1�ǵ��߃� �m-���aT�ݽ����4�p��h�Z�9̹���p��;/���&o1��ZmFv}���=E�Q��_>���Sߜ|+B���@X��&0vv���ʊ�I�&�7_ѣ&�6o!tB!�d�5�3K�ܧ���K�����N�k��_�ɺs��>�8N[��/0�g��{ޞ\��w.�t�bs�p�u
��܃���I���MI\�ŋ� �t�R�Eg�v�m�5�bUꅠh��{[g��l�[i	�6A�q��yo9�Wvȹ��a3=��N�W�l7T4��Z��F��dO����[��O�A�������;������є��c0�1]��]}��I�Z�}�Z�;�/:�]_ij�pE�Zǻ�}�7 n������ךm���|���Ӏ?�)��;��n��bW*ǔ[��(�	��Q����]���vzƇ�[f��Ǘ��䜖ZXm�F{}W�畕U���KL�9�?E�k��~���dvv|��r�q���-M��Aza����I��Ɵ�o����h�~4\�~Ԣl���{X����5W���o9��O'_�A�\O�ș2��,�3R�}�>t�fđ~%�ȡ=�QK�R�-J��T�cc�R\��4~/��*���
NɎ�UZ������}o�c�a�Y�|m�M`��8jj}��*�"�>�|���g�L���_����� ��;XȆ�Fkc���aw �H8y愸.̅��)�^~��8J���=�\�����y���<������y��QSf�����1~F�7���;֋jS���[ ���7�<�
��$ܐn�k���*��X�|!�Db��)�=k<u�fc'�c�܁�j:pA�љ&�8B�}�V��Ǹ��/��=��p�����揗�C��ǩ����ܟ�,).�8ϴ�����o�q,��тt������u�������_o�F3�Z����'���_�\kl��YS�5}���̾u����#���EG�I��cE�A4P�~�V�W뽢����2���-*���r����s-�=jJW�j��PN���&m8�-���9��� ����쎝Yߤ���]��yW�޷���2+kwtS����?3*Wӊ�`�0rhh^�wɻv���o�	Ҍ\L5rA�>�j�2'G������(O��&Ų�n�ޝ�����-�h�|.2�v�{��}WY������{M��wË�Xn�IWBXw����F7��G>��ߡ��C����+-�V{��#���&�k�M�4�L��s����r�\�{K�"�7�����B~�gt����k���ϐ��J�T0��y��D�[�cTqq��B�_f�R�qƘ+U�Pp�Q��J��mh���ScW�9�Ⱦ���ږ�@A(p�Ŧ��z�爆�Y8��LPY�����K�뻍��d�9�T����Ҋ|���u��^�w������\1�1ʁ���2���p��|`���۷��������X	���ɱ8������P�eN	m�4P!m�j��nn^s��i�i��e���H�g Lm���xr��Ï�?��7f��� ��^�Y\�K"��y#�/���\�P-0J�9��T%0� �8d<�[Ü4tJ;ږ��m�-f�O���_[�뮳#��L��oy������0נ���d1;�w�	�ۥ���4�p�����w�(R6�U�s9��9nNߍ�Lh���=�cc;��к*�S!SGOs�X�������Z_�4��A/��&w�!���s�7}\7y���Iδ��%2���'˟�L��DD�<C���7m��`J��K����za�v�o`����2���}�n�]m{w��&��[/���7XU�t8jQ�mCqg�TKS�W�8��NP�,�,f��'j�n���0��ʘ�<�Ic�3p���	�W�5� �PGP�8s0l���A��>��ۦ_2=��� #�qk�V�L���
�5G�d>7Z�>���$��>��a�dil���^ �Ql�~�*�VbJ����
V�Z�+2��!�-�=�-�PĒ�O3c���;��~��a���A}ET�fp��_.z������/�$�ǈ��<ˈ�W�E3�����io��,����f�m��S�q��ݠd��#��G�6m�����������>�Ś�����WJ��"�e�����
�fj�{I��{�x�e�/ʄ}���%��籑��+;L(:��600 ��}���<�6h�I��ߒ͖��F F���+��k&�>��Q(L��P�	��US����� ��6є��T>���x���t��eh�jLg��St��rs�cb��a��wDo]:�a��N.��^W��cR���`~y͒�m���\��P����k�q����ܴw���ĉ�zX�M��Sx�/���I���r�I���3���7!��O�V��V��G�ҭ��x4�����o*!�k�}��nC�G�b�����*�X�[�B�j�6���j�Zڨ}}��Y�ju�������ǧ2�$�ַ��N�Cz L>nQW�f�I�ؔ+��A����+�{��9��ͧt5���	Y������{-�[���:4�3f~��Wߥ�]��]����`v�ٽI�a��F^!?�(u��뵾�f�B����Ux��N�Nv�þ"�mU6����m<vDl����u����Լ��Y�S� ��c*�'���4?�H�Z#k���\�����̽#ܖ~����y$�Y���q�R�-E��gݧ񧰝|Vpʵ���/���8y�f:�3�a_��'�1gKNO@��i��Pi5��g����'�-3�e�RᎳM�	/�`E=�Je���G�(7�O�p����z�?���J'��H/����Y2*�-�H�����~i��zuU:��0���F�n�E+v���8󘀡��7�}�~^�B���W��k[~����n�s�'�߮��q;���,�%Ô���
FA�WY=��3ߎ�ܒj6]f=JpQ�����eO3�W�:�܍�Р?��PN��G˖a ]fsY▯�½���[�5po�
*�t��tK���
�t3`� %9�t�H�������-��#%��h���������߮�<����<�	+}���鉼��
s��ҧ]����.�����y��ə����|�Y�|4�z�]�"9R����H��.�>������O>�G6x"�|}�f�7�"1TJ�u�TF>��)h�s{���8F#�b����#�.E�]���K�m�{��N�O��UҢ�o��N�'�7[���\�^�}|Z;N�/7��/!׿�-���'U���+�@�H��<c<|N)mrY	�豩�"�~��{)�j!g�!����?�Q���=\�2d��r	1wj��օ�s��\eKl�~��p~�6�^c�S��{лD�g���5��4���7�U���[��,p-Z���G�m��>����/���3n�TF������yך�m��3~0~���f�s��/��
�}��ȹ��!�#�"���!r�������wu�_��2߼$æ����Y�����Y/'LC��f�FF&�2�/�y�Y%��������$������S����q���=yK��?m��%�,��]pmv��^�jS��^Re���~�����Pj�y���1%g�ڢ+�c���0��GƐs�f�	���q�1�~'�:����{Ң����G?Q���=�ZtW�n*���q��҆�l��|�H�28 �8�4�3��}�#��
N5o�3�����@K<;#p�~�o��n���H��f�qA͖�+��j$9��@�`��8; Է�	������2;w�.J�A��)�p�s�	�ϽkB�ȫp����`���Ȍ^V����My/A7sYi�c�pa3��{*�-UJd��>��ڤ�������1��6n�WuފO�����(��ol�U�- �y�mْ��xn��W����<.9����m��.�)O���>�WIS�#���'&�8���)#x`s���4B~FGG�K�_���Y�����r����lio�Rj�o�y��=5(]٬>�,C�⟉����7C�Sm|�5S�A���������t���b��u��P�%��������"�=�h��K���ؾT�hˢq�_k��C�f��\y���}b�"��m��ZN��k6t��W��Q.ɘ�5��Å��Ε�j0�'= 	%>���H�+
������2[���u����x	8	�m�Sg��D�=D[���;���9�:�t����	.Pe�%���\?�ڞy�۳��Cy�Ev�u�OJ��G��a����F�i��<���"��iD�w�T��%�P�%�{���ƍ���R8_I�?5���BT�Q����@�yi'�/�7c�Q� �G�N3h�n��U��e� �+5�����~Θ�׾)zŝ�Q���M�������D������-L������[�����9�tvs�?V��!�<V2ω��6m\ykD�/����j�eI;�*,���h��怫��G��� �3.le�n����z�;�l�qd�Qw��-EML+R���l�5��Y�{r5P	����z������F�e�
��e�>�N4`���=��[,���(�R|lp�s�(������fa8�A���?E�f����5vqE��+}j���b'��$QJJ*����Q�N �W�O
^���=D����%���7�m_c�7�����0T�^�4	H������o�`�f��4;���O��v���K�-���셇��՞�M%y\H���5�\�l�`�ѝ�.9��ʍ����*��66]fB )��Ayi�./�!}���
��<��Ro�����!ʶ�Ӧ��ʼy�����}���};
w����|�(��n����zxRVi��A�x��W��<s�-��d!������ +a�eq.h�p�+�-�X�����UO9�1�\<�K��aENV�)�(U�2X��`�q]�k�����ܷ��ɪ�K����Jђ��xB(�h�:�9Rh;Tx�C�����u�������g�o�#�����<g�r���&6ө2ڐ����5E�dD�ٓ�bo�QGr��	� �A�;Y�i6����Qs�����Wa��*3V�y�����\�Z�t���Q} x%�*p��.���k�oM��1_6
A����C��!A�l�[��f	-
��w���km��	�D�"7��`�@�JN�EC^
�v/��6��9{' ����z�5��Ŕ����rQ��q	�;�$�vXh�Su�;�Q1y����H�jH��9�'>���xV��F�8�p����q�������ZSK>��粋>�zk蹽Њ��\0WkD[�/��ݯ��7���&7�F�qV��r�99���o��U�a�Y2@D�j�{G�Q^r3�J�]#���܆l�t?O�b�CG~���n$q �'(���ƥ`�l���1c3���
�;8���2k�G�S��)����X�����������W��[�.�q��8�^0�/.���쨅���#"��W��#;��R���R<j���*�%$X��0��~XW�z�jZ�-��!/�ə1��[�`�SrJ�H��n�ߏ��wsA�3�)�S<.���T|ϭ�G�_��$;���֥����e�׿�Xŵ�)W	?"-^�;�k2j�����X)ҁT{ɻ�b��,�0����^�;ݬ�Y��^%�pJ�ݚ�Ǒ�1 %Fr} ~3&Dȓ@�8���x��O��&���v�eĻ��ʺ���L�N�
��ؽ�7D��L��ˑ����L�7/9�b�S��9���1����9 �q��=1�������Zq��-Z
�Nt���f�H��`�ҧ��[�4Rk� �j�1{��~�[9��6�L߯�'����~��W��Fo.�����՝*?��Q�q@�?
B)q>7@�n�9��d�,ݘb��\�8��8D��c6m]�?q�cx�VLc�Nҏg\�� �eV�EE�Y3�'��y1R}3�F�m������qDu܁װAf���i�Κīmm�*x�����2����hڍ�4�[NY��m]�G��z�g[Y�!��`��R͋Q:G۽���\;��g�𫡰���h��Κ�����*�2^�U>�q)ς�\	�nN����
���	-����]�L��t޹���镄]_-]+��@�VVl`g�e3uN4V!�xW�R/�H���؞-�]屢*dVG����O��b�i�bD�yb">�+;̒��0vQ�
�A���^�2��j���nϔJ�$�����Ȯ��Ɗ����f)��oa&�SqhΪ�
���l�H3̖]�c3�ĭ���9;�[������b$��%z��CU���{"�)W����`��P'�N�s�����i�=����v�A�g0�V�ĕ~; f:��\+�Ȯ#eJ�Ҧ����N�B�?�D�md�vώ�e8�p#��0��n�=�r6o�?�kD$�&(�۫����ֱ��]��УF�����9���\؛,i��7��Wʹ孭l��c}Ѽ�Q=�@,���G���� jo�����C��7�n��x����D��ƛX�1��;����{�j�c"ū��	\[~-��:6=�.6�ܥ�F�������G����:�M��`�C8�R�r�����(i�Z܎�7�Y�3�ZH�ϝ+aRy=A�����>�F�)>�,Z��b� �q��}�]�����;���f���֝>b�+�P?iN?��L�J��~v�r��ǳ��S	��L;!�$�� �RNxBh,"Eꑄ\m�$��I��-�������o�H��B`z��������Ljޑ���R!��J �k�%U����BD�*���L�E�7�g�W'��.�5��i5����͵䡎�-KѤEz���GB�詟�SUUURM������=�q]��j�(�����t���M!���TORP)?Z�(�gz\Ay� ��醴�����})jC 
�e׫�����/�{K0&� J({0#��wB3&W<� ���d/ͥS�G��Q ���~�]��AAϟQIA..��z��]p�,�T�ߖQWW�8��l���Tp>>|7���Z/��u[ξ��5]ڍϖO���C�����!J��i=���[�2�P[���ޜ~��h���!1��y3/��������.���jb�TGb��lh!u�P��:�^�g�x���s��O.�:
������ZZ2�j���P^P��Ɩ��ycv���Z�� %��.������G���:�z*�����!�|-��I������8����G���Q�>K����H����Z���0�D&#�G���;��d���!�.�ݐ��%n	���o1�$�X�����O�@2/�Ã���2]x$g?Y���(o /�����7s��l�E����%;���wg�������:*���K�]/�ѹ�6�Tx�������O1���&�ʲ^�N��f�;�K%-���g]��k?8mpB�ÌW?g�"#�G/+��洇R��dW[�Ӻ�f�O^�+phrXu��i�cq_z"S�#�jdh��N����[�e�
�[j��ՙJ��㦳a�z��U�j��P���h��gݨ�s �N�����4H��_��w�����at��k�n��	&;-z��7���eȒq�M6�ld���LW�@��S��gJ�yo��\�V;Npg���ڭO��n�?����-���w����Hӭ��ʬ$��{s����uV&48z��[����N��0���V�x��j��L����p�[g��S���8��S������-C�Gɢ�c[�w8V�iۚsW9pW�8��}���(Ol��%'ʅPb��Q�{�~����>��Tʨ�h���?RZ�����J�)o[)MfPN�b3�\�ND<Z���p+Ln��8�;[3M�&ڲ�'E�	���!��ߊ�
B�'����$��9_^����WF�
�K/�	8���/$0�0D��{�2���7�w�R�XD��7X,��o�Xr�5�mp��l$��}}�j���ښ�{{'�����9�-l��_*;$��@�>	��`X�n�G�ݐX�����.I�W48l�vǻ�����o�
�֤�l۱Y��"���I������BR^�Aj�}DC�� t������zJ���`@�t(�2��E{�)����R����/�ʑ����#C�6�Ս�Fi�+o��K���iĒ��en�Y~#�׈$s�a��(�fZ�P�߯xmN�M�Ap�q�H
��2�J)����Ղq�ɧ10�;^;�<���������F���\FD��+���--���~|P�~־~&��2�޽;~�ϓi�޽��Z[MZ�	���K���`������:�L�̢����*&b$:1Lh+e�|@v�!Z{b�="��v�����v󘁟pQѧB�?�=����O�F�Y?pi��^�~��:y��;�����wc�gW��U���?���,7i�t���xq�	F��jd��������%��}�-U,�ho�`�������П��p��V�>M���1�?�|��j��F������;�|�L$��3�u���3#�,+�e��@�o���o{~&F� *�X./����J��:�!�a{�|��T�?���C�@�m��[���A�ߣ	����Sk�蕪���\#
���Py��o�2�O
*��	���C��z���oz�87��ےnL�X�6q�32Lts5 �M
��!�gݿ�)4�� L��Q��(7�y��>uT���Cj�r�F�D���clr�*sP��^�'�ı?����S=�M����f�׍4X���qAε�"�Â�Hf��i�JR�Ś���r�g��$��~���ڈ���S!���h2��QF�A�g�N�I��H���jb����<�0�t*�R�S�@L5p(z7tkd�m1�qWEw�g%���#="t��O������?�~�ƝZ��k�f�qMe����W��N�1�y����!���uƢJ��X�K���'�S.�����h!��R�A���S!Y�[�T�#Tf)tؕY�z���t��y�I�f�+ws��=���{��'+�i���;Խ)��/�jmI������Z�
����u�gm�$~ 9��ܢ�Pk؇4���<�Ζ��x��5����Ϧ���xIՏ�v�Ƹ�\�!�!EP�g��Zp��9���^���n��{p� |~[�=�J�Y��zIn��d��x�������N����mUX��h����S�(-�NYc(O�F��ҧ�?�b�%��`b s�h׺����vq�0=��g �5��U!��F,a�]/>���=*g�(�'�,K��Ls�Ў�����y;��z�_����>>��ܠ�����4���M� .�	�Uj�����߶3�=�S��vԉ��:���ǌ�Gx�b����d黙���	M�ԁ��s�a��gB���Y��C����OW��7fG��],1C���FU�h�5w�UV��z'��C�[�,�I��i�3c4�����Tx����[zp��{Ʌ'�|�!o�"#���;W����r�P�4v��I<�[���$$����m�*��ڤً{[��7���Oj���L*�u�,��g��v������-;�)"���z ݍm�nx�U1[���j�y����)[�,��~�^�8{E�+����,q�[
����8?�<�]f�l�n���F�p�1C�XG��K���p3
�)	�YC��_�w���>�В�IYܺ�M��,-ku@��0�(�o�c'W��0����6is+Zb��o_��߁t8�)��nü_'�YdP�!�~�gN�@�C��Jk�im���������3�W��V��kQ�$�d"�->;UA��i_�_�V�<��� Z��j�c� ��{�V�����m�V�t��_��v�}d�{�aV>�T�-�}�D��*�8�&H�u��	�ﾅT|�8�����)qH����"o��$#l��[�2o�qX�P��H�"��+g�b�]n�Ŗ��]�W;=���Wh��7oCa����qX�t�h�kI��C�GX;��γ8p�XU��&��#wL����}���s{��"d\u5)��WZT�"E�Dtꙧct�T�5�k�{�^��kj=��\����&�n!�-���$r���
��s����3�V?��yA5����c��?Q.��{�x8,���0m|q1�I�~\�����Mo*�ї�X~*1���.1"d3��9���8&	�:�5�O[���o�Gb� �t*קcY��M�p�N��1j�U2�N}�G>�&�NʎS��HE�,�� �m�a�>����g�TAs˦���ڙa��\��k�z�jGU����Ұ�
���$��&�����7a(T���ӽ�r�sa�8F�)����*���X�=�%���!��=�Hl�+��{��0JQ�����M�Y΢Eh�v"Y��NT��nϔ��o�*?����e�`�	O��%T�^l�ȋ	%�j�;��B�jk!MUr陱JJ7}t��<RՁ����KΖ���<��[���{KP�[�ɥ+9�b��K8�+>��&��8�SQ�ѡ�ɜ���uX���~v0(8"�Ű��*��2��I��/�4�e�\X�o��u \�]�ͥ�;�U�M�bs���
�Cx��c����\>����dH���l*\�8-�'�����&�,��y�]:J+@�hn�n֒�(1=qh �|(1�O�{_�5�h���>eИ�ݜ����aG���#&�w�MGx�QUI�|,���H3U�.jJ��R'��}Ú���%��Q�C/���Dޏ|	{?i�9-z�:(��m3S^�`@/9Goe${�1��шǽM��G�����>r�7�'��@8��~< {�E,��D�X���/s�z���@�qPr���[�>�t�7@{��4����qPt� �/-�z�V�l�/�;��H=�����s�BZ�d�y�e��S�֊m�8�]cL?;a���ȆE �F�A�Y�������]��M���a�ڞ��.#5�3:X�R�e:���eֱ�������OK�,��8���q�.OUxo��-�����������h��DB��ƵGSq+�u/�dɁ�L�WZ��W�V2�*�S�����Ӗ<f)\"(�۸����������N��,�'ȑl��Ź��eVG�yQ���e�Y�"��������PLe� ����E�ђ6�*�!k?�n�J���If)��pcdHꗧm2ϛN|��,��Rea���=�Zpˍ�q���6ߝ)z��q8"�ʫr��V�)������d�R�Δ�T�>��4���~�� ����ݝ_q^���lpjè��l4��v@��Xzt=�v����w�����@&0��f�e��?%4-�Uy�V�w9���mݘa#�=��(/����i1���nV.m�G��rA�g͠���n!ҝ�z	"���M�������$Aч�Y���l��4��QwJ0h�����|�g!R.)ݐ��yl@�{6����LI����
ʑ٢�����dsw�/��*M>q��ɞ�s��c����!`�7`�WT�j��X��O@��K����sv�?���F
|zU577���)((�S�Y]1z3/DY[�X< ܞ�*:��`�bCF\Qq��o�i=���~�?�!��[�x����Yl���mR@��{���k��9�6@EG���#4|��X�{Q��v�ս���/kg�4{� Ö;?/�mZ�Θ&��y��5��I`�L֏������	W?N�I@1TE_{-��:�����K��t��Z�&Ti��V_2�+rgS��{oh4�^��8 *'�o��&l�"ްb=����>�\��L�(��~!>:���l#�(����х^%t)�޷�����3?Ǖ�:{wG���jן�FTȾ�'�� AQqo/s�����T��p }��hO�F�����g:�6T= 'G����}��2�����t�|����:���;$���u�*���OG���yPcc����6�����.�Q�0e�C�u;g�e:�A��"�%I��ړ~�\@x���Ҏ��ɰ�xȨ�j|��ɼ�f������ �U�����hM�ῥ��ܼ=is��s�X��!�So��]�P�'gM�e��w�e�˟r{c/ɪ�*�#0P�O�)|��:�s��/���dTM����h���۰�?0i���)Ya$F.䎘U�j�� Ӿ龩mЙ}w�p�ёB�iQ���(�R�#�y�Z'�=Hy^�Y�ɮ9�j,�B%��<ֈ}%5~�2�b��)^_��i���*++�Ӿ���@ڮ�`ܢ�ϱ�~��P�H����9�,��v
7.�.B�d��<]�&>����к�3R��5��UI��ʸ��6���6���|M�7`Hg}���l�rn������&k6�y,���v|zʐ��g��I��H�2CD 7��B�6$]Y�n�B[7o|Sqԛ����`=��c� �پp�����(Iٕ�v&������O��G�Q:���]c��)��uF#�O��9;��Cm���~q'���+L��ȳf��n`�� ������ ]ʳh7�Ŕ���fi��a$�Ö�f��Ȗ"�o.+[*�E��~؏�,��j��:mA��[h�IT:f���2�2��������pLe)�����wq�eF6�5vGZIY�l����g��s4���	��8]��S�8�Pt����M�>�@��Deպj���(����[y����V�mJ�Vp�;�n��LD}E���Fv��V˵�ܫ���8/��*Hl�aNiJ��>�ln�y����n��o����j��e�����(�q���S¯GvI*nmu�K�63����?�����|�cJ:h�� _r��z恜=3R��k�;��H��I���ǌ�軕�^«���؜�-�#��V���J���2��C���H����)ö�\��[^	E���bj�.�ȼ���"� ��!�MƓ�K�W�G�oy��?�B m���x�~k ��_,.]��|��>��{7����S6��#���0(L�\�����8� d0x��uin�_���_]K�y3/�nޥPQv�n~��}#\,6Tl��c�g�?Β�p�kF���$�FB^/̀_�Bt:��$���?�v��BTH]�O��>�We�޷����2%(C�i��4pl�X�b���E7�̦��-�l� ��V!�$~u8����,7)ʐ�]~w�"�cY:��pM���l��83���-'��ZKC��Z������3��kw�%��a��Ht�vZ�p�E�l���l����f�y���<+*���8�2����a�Wb �m��K1��x#�vc;nH����׳WY�{�NC�U=�(s��UlC��U��gC4���4��\:���"��ޟ�oϼ���F�	.����w��������	������P��ӌ�;z$���|��'�5����'Z2����p���"����=��$�gpͦ~]rmW���GJ�]�X�=#��=���}���23�b�F0�2�Y����h�[�}�+!~������1�b�3���S�����˧��V��W@�P�\Foz��g�[O�(<���i"/��KD{����J�Do�w��C����Z)��?��2�J�3��͐+VE���r9��"�w����r�f����f>��;?$d�+N�k:�UQL$1]�E�wF���|�RR�)���N���v���궇��<��� ;�]eG��l���`��Hg���;v��J����=eF㬚��:�E7��bj+��3���̓x
&@�h�!5�Y��e��G��2�n�E�y
s�`�� �T*V�Ҷq&��>�C+���vk�,�V�����"�*�:߲�󥌃҃������0���b����٬Yt��- Ѫ�ཀྵ}��d�͉���O�6wp��۰	���5�@Ī��7�߶u��{fk�~uY����h��3)� GsR16^��'�QAs��4�IK����3}<wcp�q�ln!���N͐�5"��U3��[��|�= �<ӉMb�1�z1�Ф����4^R�x�]������2��8��ھ�A�ݲ� 
�Ϟ�3�-E9-m-����>��;�8�%�p:��' ���E^d�JX��mg�$,�6?�W4�j���(o��i5�?4��R�"��)>�Ŭ�iG��M=���6&�ew�'O����~Ÿ�8�\zo���E�k�qHyb�f��cP����"�4M���x�V��Ey���-ބ�aɱ@;L\�W���"C�֬�}1�w]�YI�W�$_q�3K�Ό��陃@
1/.�=Y�d���m���[�X/H�*g�0/1�??�>T\d��2����R�!� �ȟ޵P	8�hӭ$��E�oqn�a����c��a�z�|=_�$�wB�)�X�rZ��>򶈂�WT���ftR��
�3�w�j�8�@83$��&>��̆px�����b��4F����1����{�=	Jr˺8�4�g�o��]�IzO����.*ഡ�(U��	��x����T*�A4V��n��I��������J�\�;�h�HK�[E^�����Ɲ���c��~���l��'��Ǎ��{�;�s��K�u���Uc&w���1��U����#�T F�(\VE�w�/l��q�VQ��z]u������L����~l�FD������,��wkGD�e:�~�;κף@��`�EC��Y���>�Ū ���
|4e�F�_���[������)��f�Kiy����ض��-G��nnMՍ}T,5V
�j\}w����	�K<��������b�ꠣY�����;��vtww�����Ii;���}��(���I�Le�
��DMz�u;����F�g�G��c�	wZ�����'X�G��u�"ْ�:1�A��Q���=��4��c��+��O�ϯ�X��[�r���SL�
������?��
�df�0�fLFjdr��'�X�s�(�b6,�q [/}��)�����X+h��t2/D��G�i/�#��o)��HMm&]T����d�Lȡ��g^Ԁ���f-��\"���I0rhj�8�)%�0�e}s�r#�~K���B��Ta�de&	�a�~�ح�����Ϩ���}����-�Pv	%�ъR)�u���ʈ�b��+f���G&t������K���0
��6�S��ύ��o�j��F�#���D'�>`�M�UVqS�]�����t3���s�����F�����X ?,��B|�זk��GvH���
+��|~��ޖZ�v~�zP�����ʞ��w�Fm��xz������{Ϭ:&|2��p@�f�S�~~�ѕ|dM U�,��8�y�bn���6�쨧e���k~��ʙ�}�T7�������~�tS��/�8��Y�h�E���x�g���0�JvU�W4�-&>Ina_ޣ ��j ��^���oNn�;���e[��f��zM�xih�8�����읹� ��I��{ξ��...]�yq��u@o �F[����bI  ��gw��K��̳28���FU��E�QmmH ��!��ke@������\u=�X�v���)|�����ǚ�=��U7������7�H6g�>��������.��B���2.�Yh���n>nh�����{��<�	pT��q�4�)��j�I���� �UpŘs�oB_cL��}�{q�?�i����9D���3l�g��(v�p"�׫(:�Ec��,޸��r\?Z�k��"��Vޡ:����
�q<5v7c��&ݟ�dQ[�r���@9���~��/N
ȟ��U�ꖙw��8�:L ���i�;�ܮF����s(���:��~[a%�&ӲS��&�_����AǻN��Yr�<Ff�7g�O5446.�:����,m�g30=�ι;�|�� 4*��Nv��AZh��{������O5z8�*��WEZi�./5V]�J`£�iAZ�7"�F��������.��U�ݱ��*jÂش2����k��=���C��
i��/7��Z�D�t=b�g3�^?�������ijI��h<�%�@z�k���g�"�~LQF��fxh��s�r��t�H�[/��ol�6e��"���2j��J����.��.��
幥��ʽa����+��C�Q"V-%���,K��^��/���dگ�i@Z����+�~�#��@̳�OC��k���3O�5��@�ݵ�Wdw�Q�,��������s
�!�[y��L�dw/���~;�Y�l/���'D�7��'���v���Ǥݮr6i��5ˮyI �0�m��1<�������;������ˀ8��؏��q5ңР뾓����E� a0��)��C��<�\M2!�r%��J`A�"���o�QY[LBGG�,j(�_k��߉*����`B�y7���jS�6��,�4^5[���ch��f:��?��uy9o_������c>�ei����D���㚴Ov�̜�PGN2cR��z��4�.�-$؋f���s��$��x�{�ޅ�����8�($%�k�����mU�&����m�	ue-ctF=�Z���@�x�,kI�ឿ�

Qٸ�p��H1F�̻�U�gbG��2wB�ZG92�Eri���^�F���݆��#K��@8[�+1��or�__�,mX>��g�g�a�^�w�z��>�z<1�A�@5s�y�V���&l/����]=A�Xx�\e�4�n�K�\��@3��$M�U���۱����ʺ�U����H �S�"\���P�����r��TO���q��ٕɼ������w�����{�n޵�.A�9fڃ��N�zÂ�����*W�V,	��E��9g)��EH<�ԗ�F��SG8r!B�d}�3�/ְ)���;1$+�g�CsA��(�>�Doϰ�4ub�HL|��q��n2[ߘ5�f�K�}�6���Wn4nID1������Dt��ްk��KL�Rt��
o��M6� ���~"���k��u��s��||�ݧ�L[�nf�Yas�A�Ki��kK����%�x���y��7 
-����ŉ����A�9~U���&՜�,�����1��_N�>y=d��_^��L%��F�q�A5��VP�%��.���߅M�N�	�򇮴ۜ$m�8��� �����F�?mpRh���<ᐵ�P�s%�Mf�4�L�,�$�<���,0�+�h�]�����,v^�ѳp�p\�D�������~Z�,�J�溝U�Y�e��8����v�Tt]���Omx�8�e��A��e��#R�g�u�m��;��Th��j�>�wx!���e��^�#~�� Q�75�t�7���`L䕚gF�Đ����s�@#�rÜ����И�e�}6oo�vl�|{����a����*�Zm�ƣ�K�ķ4
,���DE^AM���=�UOʪ�=+���7�;H 'E�sa�W��N8�]̀��@\���[�؉d���W�2\1{�j����8K_��^���ؾ����L,�������4tttj�2�S!����NY�7�Z��=է뚙����W{Yܻ��ۖv�^�WY�V>�N\)��\Hf�m{˷\�r����s&��� �x�3[P|�2�%۳�
�5�W�.�Do|���7�z��l9oH+}-��������K�B"u,8�!�B���҉�dJ5�i�8	7KS��\%)���m3�of������=_�=�"]�s�x�t�@�o�s��d��e����;V����(+�m꿁���F;���/��-��d`H9�,Q�J��ݦn�L��=�(#Ԭ������!I��pI7Mߵ~�WBO�K��K	T����:�- ��R3՞*�������|+y@m����+���,zob"���>���7�&?����J���m�G�0�W��v����v���C��I�>|l�)�p���a�j��1^��n��� ��t3o� (�L�}	lRnwoݜ���[�zE����1��("��Wc������Ӟ�&�/��s���Q>$ڇEXF���:��4�k5^��6x������I�Z��] ��	W.�w`���eҙ�k2��e���B@A���.�dB���h6�����s�7|�_v��5���.��!�3v�5��f�-·}�f"!���;�^�����X:- /����KӈgƂ��~�,�[�؀0����I >}����"��xΤ���V���t����}�����D��9ҹ�~���Qh�j��k���M����"�/�j��㽮�,sN��?@9B1��3U�o����o�'z>���i�&��cW$��F�;�!`�z��+���.:c�ON�ERP�[�	l
���1�W�ꪴ�a'Z�+А,�������.V��,H��L:�D���6���	��HƐ�*Nt���8�ah�e�|����K�]x��Ëf���?���d_�ǈCV<�4��Q_���U��b5;僪i��I7;�(�"�D����=�(ͨz�������`OK���9w�̏�L��)4�Y[����MXo�l�;�-�l�C���ή��a&K�}W�=�r>��z}Qi��70:I-��{��aN4(.�&�bn� e�2S��`��<�
���#�_s+���ܵ7�w6_�&��ggZ����Y�M�(�+�{���)mܜr6.x��ߐZț�Z�c=𕛏v7`u������5o}����!"�+"��?��z	p� �J�Cl;�I��Iz��R|��8��Sr![�#g��]�	��G��ωV<��$'��)�r�8ЇXA9��+��F����Ѕ����������l���:��YH\>��}}��B��+�7���+%-r	�Vv��Z�d�����(�a���F�1��9��=e9�L�LI�[���6�+�����=-�bl�wD��Ȋ����&>y��l�<b���T�-'rd��[�!IҼ���_�� ٫��a}��|�ʙ�}c=֮�"S���I�I>��ӈ/�ſb��H��r>U�(�8=/��!�0�j���e�w����oq���T��H���	ּ���*7`�)�H`%�<\|?���d��R]85���hV�I���\2nz���77v�����3��C�|n�b�
U��qx\7�_A��t��>�DV���\�&|Ua���K��Ri��l|xK�r��"@�p��H��)7��9*W�G���*�G)ZI����]���od��0գ�",��Z����y�P.��v���R���/�E��9�iir�fO=��,ME)�H�̿h���ΧM�P���*r��P2����^�#r�m�x�eX]@4��n޴}7�Ϊ���E������ZQ[��;���D�O�����I��7�/)�.�dW�$Ƨ��w�x��![YƔp\z�;h� �����t,���`��\�AX��8�܌�*cI�3��f��gg��r;�>�D�<�(U��Я�6�/W"�nU�M��3�l�v����g'�Z����h�g��r���^�x�Dy�.'K��Mg5Գ�c��g|	�S�?ʎ�tCT;���S�9[��^ɽ0QO��MY+������k����QPRF#  �"8��JI�M�Q�ъtMDBR@@��[jH����a���/�<��{����ڟ��}�u]�9׹g(��)��6w�!N��
��j:B�1�Eh$��v����e���V�F��wn��^a�Y�!�:���<`�Aj(�˫)y���x9l�TO;�@t���I~3]<i�!�����(�g�1�0�'4��<`�Tؗ.����K�{��˙�<>���I��p�_��ɡ	$놈=�{A�فE*�G����!gcE�U����ڴSSx*���Qd�A�9����۴D���m&\����a���:�+M�	��an�Rn��~5�n��1�=l6p�vu�t�W��n,�Օ��ɓf������`�]���~�a�ْ������^a�����W�Pѝ~�L�� ��Y-���=	�ƾO��3%�X�S��ckLj;	���C�j���j�.�X����1��eKs�I�[��L��r�e@��FZs�!����s�2�l�A:l�ӸYf�9ODݎ�xa����7ɗ@�::/���̚�٩/��V�7���������B��;0~�����=���J��f�2˨_�f�#��~8)w@]�f�+�G#���i�����:l��k�es�v6��Z�K�������᱉���A�Ў�`����I�p��:Ż�N�	·O"՜�7+��Sď��%����G��;�9=M�~���e�������E����Lîe�����Zlشi����IK�ִV9w#�5�q�:b�Ԓ���{�[��L����e��Q�[�|S���fg�/��,�������6�+h�=�k8��1�B����-���ٞ�Xk������p��fgN����5J�`��C`�e� �46�w;z��٪3�6{W0����p:Mth9+�Eܧ}���&,��±x*�b_�)�8�́�gc�٬�
�2��gEe.�q͟��%���&�����]�2ɍ��?��G�����:a�Ӷ'��"a���Q���wv:\>�9QC����y��5��٥<�)),$����VǮ��3�655M�k��y,�]�g_�_�B7o!�'O��|/9{܊��;�����]-�%<#��lߝOU��3��_Q��!�\@cw��t��Bf⧌�����I&��}��8��l��kr	�l�"V��f�~X��&9L�CX�V$:�W�{��X0��@���`��8+��б呫���N�MZ��� ��;��~�|YC�B@�}k�#�e��p�|:�0��g�'�`�� 5�ō��$Ǔ����x�X_��Z��Tx�D}�I�v������v@ۯ�ݪLc�Ќ�)��ˀS���ޜ���)�m�l���Ę�8�]'X�b~
�oc��rk>��<��S	���ދ�M��b֗�l�ڋ�>'����ӈ�-��┿�D�ُȯ���|��"��/��cہTI�����d=bV�kll����C�B�����oB�U�`�����͕s^�XE���T���� ��(- ����V|����C?��{� ��N")��Y����,��� �aO�]��}S�Ǎ��W,ޏ@�v%��L�).�^+[�_{.�m5��Bߙ��/���|#ߑђ�;i&�s<gV ,�Dޤ0<b�g#�)��lNO�M�Ma���*N[�=k^�{S��,�q�xxK���~��k#��3`�Ϣ�Ʉ����.�/���e��#r�����!�b����_��)��f����Q)�/���S�Un�mZ�S*	�\,Me�Gy���tv�����5R��if�j㡟5l��0�z�%m�3V�zu2=�OY>�j;�оo��8}��A��z��2$���,���������n����w�(E|g��݂ى��	F'�QM��&Rn��:a����s���0��E򧞯
�R��N���9�VbZ���}�\Y��[x�p-��_M_��x�r�ȋ?��R�D1+>��w������]I�XZLY%�Ʊ_�7(�I�a.����z&����}���p1�]��K9i��^�|��T�~3n�a��:oE��&��KR���&$���݂ ��X��b��u��X<�n�� �3���D�bmZ�Nu�����@p�;x��~P}�I��3ӫCw���՞���L%I��B.��,g/_��ٞ%jn$�mG�){�*x�L��Fy�Nc+/Q�eU	8&ެJ�·��b����w����z0.m�W�a���L���m��@����33��4P�*���o���;�2�c���]���7��!�2��Nb���(]�]yI�>��|ЙˬG��6��{S;�ù:���f��h�@hp���+�&)b�nZݽ	�8+�HCJI����Z�s�L�"��1HØ7B�`�6,��� ���p�:���{�H���,�
��U��=�d����~�)�|h�7�����@�3eP����l7/5*-�C�R
��[�d���Չ��fnHK����{7��6#F��N1�`z��"��0s��Z����@G(BU���$j�C��8ن40���K�X�{)+_zv�S͎N\�ve-�bWn�^��W��	aD���@��\�k���Ru�ڤ��\�怖��0�7�dޫRs��YY�5�[B����x<�v5}-�+\fj�
{�W+>����E��깯�T���Q����8ݸ��q��� =���]�F�����h��7�G�+����O�4�c��5�C��#�%� �;��d}z���wlsb��޳0����Zc��#yQ���4sB1���f�Ѻ�����$!^���_���q��%�,�`�H;�ڠ���EqK�����\<:]�@�����??Jz���[+!�QE3�2��ڸ�țY=�udn.�vힾ���I�|=�}|KE�@��^�{�p�g/Q�t�c�W�`��� ��ݝ�0@�
�۳��@j�c��͔�� �7$|%�^T�r~C?5�U*Ш�[����`D������ꋳ#li�|�w�b���5���5�+ߖ����y��"/�E��BM�Cr���D�2d=	ϫ��s�vpB�/ޑ��`-rt������|aL��@%�i�w���n���kА��)9c�L`s5���	��&�z���P�Y��ېz Ey���=���[��q��_w�S����Է*wV��e�y2a>�pjR��n$n ��[�.A�Х%��4o�tO��.�MAg4(Q����N��Ί���̌~�5�X����DJ����n��м?�D��.�ۧ*�+;����[iYT�k�@�VY�M�����g�"��TZ�>�Rʵ�9S��n�4p�\3ܼ��;�c��	:��^�A[��d���1s�yN����N�����Y��C�1��v��ua�ݙ��\��MC�^�������4oK�mc0*L�>��f�u�~c�zz�"�8=�=$����t�׭�9��MͽTɌ���q�qVK�:��g�J�r�;�$�(A_Ι������C��d�?ό@MS�D|K����"���'�nR�\�B��c)��������
.6I�tmj��2��a��1���������ìP/�T�'��u�:/�4�H�6PR�<�^�Ef�����ĩ xg�OY�u�E��ƽr�w�2�w|����4Vm��e������'�}EjX���5������Lu��7�L����x��0צAX�O����Kx�k��E�,���dћ�k�YI�x�3��+�<�My�|��"+�������^�� O���}�U�Pg�~�z��>떰IY����㫼�������t	y��O�Uv���'�ɀ��JI�c[��]$l�������$��#4ƞuY�x�e��ՋU:��k;��k�X}��B��>��{�~�. ��]Џ"���y�����SC:3�Iǳ���r�X��5
k����RcE2���\����=j�%i�X"�$�\��>��(�f�ff�;b%����j�v+�|�f�����!j?<,.>@g�Կ˼�Ҳo5q���Wov")��MB�]�0���|��~������CQ[���lD���D3����3R��jd�V��Wd�7�?bG0Us���G�]�U��~��WQܒ:��3�K<��)n;������u����b�q9mP�f�֮>GJ4�kg*�=�ˠ�z,*l�Jރ�0��)յt��u�ס})���u��3�XKs3#o��Pܙi[HG���M�]v�s�����p����G�X��7��;$IzYM���cw��c	1}�]�c��#]B����CPEc��i�����������i�}�.f��?C�k�;=�0yvU������-5W��@�+I�����N�g�ex;}q7󖛳�q.�,�����$�$�M��9�S:�W�kOO����y@l�L8�Ǚ-Z5N.Q��G�s{"l	%_ź��=ez�W�� [
�)0.-��`5�r?�oH��}E���E�k���h|�P�& y��tt��w�D`Y?�w�/�P1�w��=||*�2f��o���+��}���yvM�"C'o��d�V�j��)���J��N��#�#�7� ���K�4��9�<��ô�P�Wg,'dVh��n�կ���*�"8"� t�k�S�'d�����z�?u���-ݝ�M&�|�}sׇ3��7�ܝ-�M�M�\��Z7w�4�� ��W,v���?+��>�/���^���*'����J~�4|��y`�����bF""���.]�� N��=�gyt$*f��闶�k�-/8�B(^�vE�R�߅ː�C�I&q��+Ug�F���'�I�/8Hi��#�4�AM�<�n�ܬ9zpfi{����/�n	w�;��F�(^ng��-��O=�l��r�Hu�t�s�a��F�F@����N%�5J�ʰ���t�D���>7@���X���q��&7�Qq+�~�{y#*��E�U		t�~�R���???w|��yr^R>Vj��]��{�����/���ub�=���O���mv���Z_g�o&��Vw���F����@^ ��[���`G�F�A{��F�������ABV���2��V ��M�+�����N���@�Z�M��� ܄GA����h�k��"OGbH���A�d�s���F��K�=��_ɑ�,:��D�C�En9G��*Kd��M�����{ؤ������A�ՠ3��4�/v6�D�Ž|cV��&�}X��M�Ň������KO����If/�1���8�EB�Ӥ����򰢮�.�,sǉnwD�M�WV�[ļ��?J��]'>7��[� :��Nt�V����{<��T�Y�%�~J}T�
f�6w�\��b��Y�l���д�z��)쩙$^��**�G�uHm.����}�7����,ڏ��Z�C�\u�4Κ>��j��t�y�T��aV5GL���\+�5(w�p�JQ;9��<�跎mi���'Y�� `�j*|�UZ���M�-�us��V.i�]�RY*q������<`�����L��ݴl@G��u��e��Pcw��p�O
&0�9�yк$�Lt`8�����v�0��&��&Ή���i`��%,32*RFL��L��I�_��oxހ���� ��Ic�l$�v����(/��W��7 ^Ka�-�l�;����(A:��۫)Ş�5�Nab�h�^�$)��ɖ\�<>G�f?>��z���`v �F��۸"��o��bVn{�1~U��!.�ɢ��F��5o��fQa.��g�GlYu�"���eN'�j~����M�j�wͶ�n|�sO�Z�q[ى?�M�tM;(^~s'T3:տ�5�5�����d��ٯ�@�˷��η��w9wӷ���6�,?��1r��嘑^k�K�q���[�j"�`n��1.\k%@F��3�Y��^I/�xX�{�0�Qp�~V�QXFR�
����D�ggĹB?�'�MD�;W�w�J7���K�a묦R��=��q�}�ŉ���:Wd�%6��b��V����)©ͱc�ݺ�Swu�Qp��=�&H����m-*6�;��9l�`�����9��o����L��M�[�d���W������z����}
v󲡜��7�+�n�3f��Z����$��6�=��=����l<��*%�Ԣ�� 挰�N?<�b[�~{�}�����"�I��v�R�Tظt���C�q<��QͰ�g���3S3�8/t��o�k�؁˗ 1U���&�􁯬��NY��0�K��Q�����,0Ex���8 �_��^�_�_i0�:{�oқ~C�|����+�J�tV�P�7m��Vji�.uI�I.���{@�F�	�8q\�(v�,!���q�.�/��s��m��|>r�kӌ��dT6pԫp[�[*�I���[*�n6#�rƳ�+<�9�IՊ�n��6 7��NsW�ax���#�l��[��8��K�t�G.�@"�%�:�YJ�2O���|:L�'�UI1[��j�i�?
]K�\�}.��x�ot?���I2�VCM3���z8�s_̢��04ҹ:�m�ӷ����̀��p���9;�~'��K<Cs��{�m��/%9BS�`y?�!��㨳�ѝ��Po���a�$�N�+vc���ǲ��s��iw��A�^�����b�`��ݬ����F�\R�tɛ��-r�#*q�T�XA�U52j��S~Rv,-ZHc5D�Nn��Q��k�ÄE�t�Ge��B�g��/���o��=W����>yq����<�L���� �S��ի�5�c�/��~��^L�BA�4�lu��)ēF�-�u�ꖄ5��Z{)��m'��WA����pm�Dw<��,c��-;�[f�|��Z{kYz��H��u�}U�#����嘗�W0a�K�C�{�1���u4k>}]�ܯ�����5��I@|]�t�.��	z��z:�x�%��[ ��}��:U�Di6}���D�N$T�:3 ���m��M����Z����������mi<c��ڄ=�v�A�:R��m�#R��!�&a�����-���V�+�~�z]��m
�V���z��h۷L<����Yb�m�� ڒ���л�K�.Q��c�Vd���3"}x�{"Hɴ��L~"��'�r���'�+.�;�//r��Q�%:���� ���w:���&]NZv	7��ƨ�bV�# I��dBE�)£놽Bɷ!%��R2�_�W��'%��-%w�
��yC��n�oa侔�?�3����-�$|�1�#]���&��-S��� �]��5Q�@Z�γ���[��Ϸ ~��B�e��c�7�M�	� V
~X����Թ�k]f�Ҫ�������I��.��
�^]R���&��|'I�O>�T�5�1/��4V4$ �Ccڗ�n��;�Y�vV�Y
8�]հ��C�r�	)OBg���0E��K&��чl:(kO�����.$mX5I^���U_���.�X٥ؾT
tȶ?'^װ��>6t<vD�r��>C�Uz2���HD��t��~rx�����,u$��`�;��y���
G�L���[��m&���8�T�C���/F���>=�L�p���{�ِY��q���*aGE�̡�TX�^p�!��
:�b�wAU���&ݽ��?VR/�DNG����u�O��	=xގ�/����I����ݲ{5����۩��)D��Y\� �{�b�s�N�5N�pm��z���;w�ڮ.��Z�?jJ�LW���Ow�gw�.q�$3��kA	FI9"X/��f�	٣�$r'���v9ci����ܝ��V�k�w�)�6�Xt,� 4��f��呰�5=pK�b���(K[*Yb,� `���V�H���F�hQQ�#��i�9���;+-݂b$م�+����:���R���}�O$~�S�TN^>�b�h1}�b��1Q�ֿ�wV��ޖ�w�iQ�0��c�Y���a6�=e�}r�C+`-����𩋻V��Y�4׆�<ޯ�c,uf��J���g�F�el���k�h&��%g���j7�'��O�OG���Պ��<M�����R�#[�u���IA*��"�j#1X.MX;{*%zs�f�ϸsEM�o,��@����
��]�����W�&Z��!�rdSD�B^�'K?*�ư*�0�Y�xN�����Y�̘ ���e2o�r���R�I�~�\�lqYǧ��S��1�_;�|5��n�'%�.����V8�4��h�ˎL�n�Sɂ�6}Ug-mihEZ���{:�6�Tf�v
YQ�p�����;�u��t誨��BH*���=Z������`

iV������Ӟ�YYƫa$a�3�����萺�<�2�q?\8o�"@P��,맙dZD�1�S=Ul(�Yߘ��GTY�O�}y����'K-��0��l uWý8V {U�gX"�.�Wp������5����6aR3Xp+�g���/�Q/;oFa6��Q�%��!���C����"Z7-T�Ț��uk9��B0;�~-Ó�Y�r�@´�	e����􈄈�S�X�9*{~wq���b��+*0��?���IcL�<
��t�xK? �����#���	��v��4�����+cc'LD�wah�2U_�^��|����Nr�K�FD�˂�|��^�j)q�|��Z�K����Z������Ѝנ��*������p����3���	O���}�L����:�4�nTLKOA�8��ڻ�t(
��h��l�����vY2���Pq�;uJ���Q���H�U��X�������7�g����ӂ|��t�)��`��Q�iǩ�N��(:]���ض���+��o�<}-�����&@�4h%����P�s�����E�F �ʳ�+\����N��nx�[��q`��ֵ�&d%��UԑF~��Z�x�n��ycS{�4lD/��'q��F�4>�.�s��
@Vה��Ǫ՟d�SC�&'�t�����:�I߶��F�*�ӂi� �Ci��r���&1a�\j��	�	U�����Q�bV�!��U�?���{z``�̒=�^lga�d��`���j�Z���v��,8��� ��j����@�v��}$ޛǈ���j���)q���,��T�k~�F�W Bɞ�}��76se�}������j�љj�)���q��4*`c�.�Rcb��\z�.�Z�5pKgint����������J�&A�Y�@
�a�bۉ�N�f�2����rǲ�/Zs9'��uDn��pr��睭��F/UM *E-jOֲ{3'	WCH�B�B��i({��5S�\t�h�Q�G��R������s�V�I;��͵�����%��G�>�J�<Y����cr�����P����2`����%T��@�c�[�C�����U�UD�Q�"�&�Έ"�v��2��͠"�x����֍?-�^/�MBTw~�b6,W�*�P�/��Ha�
�q�Ɵʫa$'�<()�������O��N�3��	�fs�[���w���=)���X���=�L��s�.v[��D����QC�P��u+s�a���Ы'��+��L�H��W��W�mN� q�����3�XJ-��V�V�&|O������w�k�צȔ�-�U���������h��^������Qv���0����\��L�"[�;��,�[���S�kV~ع�:�|�l�?�����FFĺȰC �0�ɽ!���/p�1���Ǣ��~�q��eo�����̉�+�}!�d�;�v�Ͱ���{욿Hę�ړ���%�XY6��d�gUF������ʊDL�jr���`���Eۊ�����4W�����ך��a�r�Cm�*^��\}ڟQ&Gcw�����\]nP%�{����J%=3V��p٥�Qu;�?�H�pt�	B��Q�+_sN�ҳ7sP��!�oi�	"\����M���PC������s5��^Af��������}�B��_ѶI7d����r5�%��	�ӢwT�(���}8������6�.�?W�\�Ϸ}��>�%&��$�֬��;B�q�wÎ������ǧR&1���h��:�Ŕ�������&�e��c#���]b�����Qa��j�q�#�>��j{�Z��!Z�7���P��
\���ے���f����#���w���R�U��#y௃�䌊���S|�@J�L��GI�rZ��ړχ$�d:��/3�3-mI�}�4���\�R�I��-��-'*V�(�,A�C�L��Ůa�2g�r����=�a9��r���d��&���®3V��'��+��UBA��"� �qRP-���o���bI�:�|7+%6��f�0�;��8]�;�t�:��>k�!KJ�oK���]�%�n-�Iƿ���}\�8�p��j�d�:K��?I�p�����~C:���U�l�7f�?X�>=ݙ�?��ƕ]�zG��5��33��/B��B��	�lO������*�d]h�{R���ї�9ش�Y�X����n�hh�"�D�Tm�U���Ķ��d�c{)���s�cP�� fc5�A��d=FW~\�:��"�Uh.�3�l�
[���RG1��%�;<]�Y�_ÒgOV3z
M�՜�$>�F(���k�M�Aq�?+؆��M����� ���QlL��_;�WdAQ=Y���7Bh�j%SCi���;�$�b6gC�r��T��خ�mԛ�6�� �K�с);*�[g�����w<b�C�Tn�����̑!�%ق�G���1.��\]=7���N�d���Gfe���H-Φ��9=�>+��雲Ǯ=������H��X��T�����p��̌�`��{��F�wىi�b�Vf�:ba�����V�����#	����e�>�zh�2�!����X}�1�h}XP7�T�>翭i��-�ZM���D+��f�9͹�KJ����ُuNn��A�m��.��«�?_8Y� Ca�g�J�+�M� �u�\����A�k��nh@hSc����j�W a3�81����VA�*�I��?���deV�f�o�ZW��
�-߭���g��׻�#����%��#�gM���N�ָ9����{x��1��-�{~�Y 9b���Bi�.-=��_��0a��ԗ�rt�C�xJ1��;�V0E��G��ȶ��������.M�x�����׬�!>B�r�#	�}�����va�|VlP��Y}�ҵ00���)�׸u��&�IVZ�Q,i�:�M�-�-(���p�5q]���s��(su�|ja�;�+b�:UeOx��N�ڏË3��'��f^���-������g^�B���{��=��<�>&i�ɧ���H<�Gy��X��0����T��9w�����O�^�����0�F�?g���ٶ��wI������,��e*�!����c�� �Zl�B�ԭ)�nLa�����~� ���u�Y5�Q��G�(������d�$�������t�z[w���3V}�������zw�a�)0���$(�^^p����2	����b�ٶ�vƢ˪��=Î�=��^��;z;�B^��#�Y�k��CS�u�?+�����χ����kl�о����`ֈ���_:���z]i���G)|eL�>�I��ɉ�`��7�ب-eee�fe��R࿬(�$0�כ�������L�?��6n��5��A�-i�p�ZM%��8��j�����c;�	�����b O���g�wG�$kYm��kF\ �,����XH���x��Ó�()�!���̷o�鿬�}�:6�38�X�mll�68��Y�$���d�5�o��ŭ91� ��=�?:��e}�Ko/�j�>qH�۸m7��6.�,�$��\:�/7�G�g��s�,an�������o� �b�1��oL�"e��CL�����9~&|�j�o0��Gv���o�? m�*������"ڦ]�����
L�ЙҦ��F<(Wێ�`lp��f͡ޝ�f��3��q ��b���MeR �V>ɒ�1]/ԆRM�}�>J7��r�3�����y�r2��Ɗ4������D�f�+�N�KIJidm�>���N�5��/%���0q�Y_Qf�̴1�L� *���ʪB�؍�����^��^sf�{����`V��>�#��Ֆ����#F/��#L�716�[�~��&J��a�14Fv���p��甐�L�4ᩍ�ת�\������v�c�b~y� wԃ8���-�?��c�6�sZ����t�=t�(ء�i�"M>��	d���I�8k�e�jn��� ��;cv���CX~����=jYk��Ћ���{�������BV�<G�=��Ғ��2�m�"W$�ѫt��%AѴܼ�H�V��rN.�^�f����Jl��]�gH�C�a�c���a��%ݢ�w>��g��^FO>5�.U.����h��l߫��@劝��ě	1e�8�b�E�6�
���C@��;�G�lM+�t������~a0EOV`�i\ c������T'p`fU��	&�l����{P����;]QY�A+--��s>w ���
-��O�w ��Cr¥G&m��o
.5ϸE�(;G�ݾ��m"�}ɧ��vU1��Ș~�G'D�t��Õl��[BY�%'qoQ�weA�'��<~��j��%� g.��F�	��ePbb�����c�K	S��!�Z����k�k۹&Z"u4b�rS�$�����;<=���*\r񴋰O��)�{j!�鹬(ъ�0D�ɮ�N*���~1S�#z�h�����|b�iZ�[K��0��>MG�v��[��.\WX^#^�������v�|}�͍bǈ����1�8)��G����
8���%��q�����q�O�5���9�P�3钒'��=�qI

;k��[�a���x���&��͔f
�$B��� ����܆�n�i����=��6J������{_�NY��Ἰ�ٕGd��Z��H�A���>T)9Eɨ��� dT7�,���T/�A��)"����9����Y}��9`?��Ӱiʁr��&k��*ዤ�na =�瓩����8�&s����}�1���=���"O����G�C����]�R�t��¡����_d�~���b�W�@9�+�<d;�~"�U�}7�L�kz����בc��K"<Xq�R"�E?uJ�3U,�T�4<Ԝ��L�Z�MI��rnb�c�^A|�\�7�v�dA
H>��7 �d�}!�lp����9r��/�nFª���{�^`��71[s�"���/|N}�=�0r�+�Jʅ �Q8ө�}I��b+Z���,qO<gq	�3Q�γ��9�W�],t^>|(�3M��k��V��￤��0����*~{�7w�����Y8���AZq�Ζ*�����7������z���%{�3�1��a2�8O��; ���V���Ϳ�m;2�e���5+rβ��=SL�ĳ'ҁ�C��Y��=zI�J�c��eWDz�J�6�Y���xzFe�\���݋�Y*G� �Ճ�tdW��l]9jlz����?�f4K<��g�C]��t�÷�v C5�r��x-���:_�S�Wq���5�=[�Z9��[7_Kxl�T1�>nT�{lBӔ��<�'�!-T�����o�i.�����fq�e�T#��-��#���Y�[>����𗽻���[8�y]�,bJD��} �9G��5yゔ���)1Q����1�Lm�
�,��M´胲�5����h����T &����1}s85ZC[9����{˽�����z���������'��*�W����ܛj�䡾�ѤW7TR+��</�����0��K@ ��kp��K$Ө+Y����e�����5�ٻ��lg�����X�栺ڣ�9P�J���0�6-�M�s�FRƤ���[������b���⻖i�Ǟ=�;M�.J'��w0����[��>	�l�i��r��t��-�!�|� ���)�O���W��G������C�#�����k�s�mWA���B����LW�B�1���b��Ň44���z��be���7�H����su�˷��D�13�/%���iu&�(�<'\A�;Kt�jl��4�]u�)N��� �ee����*7����o���xU)C`Bt]y )d�����1��N��_��59�؄%e�=	:�<�(������{�8�r�l�ucv1��������(8�n��N%��q:}Wp�����F�F�8Cg8EG��c����VvɿC𛟽�j�6��":��d��o �]�X���}	).��y^�����,���ס�����@�m{����@��,����u��Ob�7��4�\���z��U� ��5��$-T�T�x;S��ʒӴ�؛TQ>��3�g�<���9\�M�0m��=bs�0�72V��l��\p�/���3M�m y�^�̈́G��0��t4F�C4�]����T��p���Ai;�>OT㧀0��[ �E��p;��E��|c@�B�X�9��*~��<w��P�MV$u�7�<�[d�80A�aF0�<mZ.����z9���`���[�2xsc�"k�fm�2�-w�;�a���t�����i=�]v��O��ޱ�"�������o-v�|\bʛs�{�����={9�.<�;��
ũ��uIN�Eމ��it���N��J�I�nH��?ܛ����]�{�>�L�oz�`�K�F�-ߓ���o5�ֺ��nii���%�sB�r�Ic�5?�,j�ߵ���m|v eD�?���ue3��|C%��w��|������?��ޏ��{�h?��զr|���-�ד�@�����wPwf咛o?�pt+�p+���:�sE�������K�0���(����[����[��c�9f��{��6t�"ܲGK"��D�	�C�� �ciDn�6� }b��S��^+����Ҭ��n�?���Ó�C�靕��,u��P�p)�>I�]7	�v�\m�CSٹ�?�9�SR����҆��؆�ie�\l�7�fÉ�p�S�:�fSre$��wS���y1�����c�F�o襶jT��+�-R�P������F�nyB���=ښ��ٞ��Ȅ�X��J6��gx��b�<����t��Q8𜀂ޱ$�߃�Ɋ�mM�XSႱ���;�=��.�7�V0D�-��1B._c{�;�v�����+��w"u?"{��!�!
��Q��g�3��<R�=b�>������L�5�,�i�}� � \;�p�Cc�ѵ�*����M+~
�qj-ge�~�?Îe?��Q� A�"�����3� r\�e	\1d)�N_Y����v�q��u����!�L���5��Ң��w���k��P7O�p�'��h$bJ�"�R��ʰ2k��WcG�Y,�]�oBd�N�*r��Է`OD��O�>'�,�1]:[�
z]Nx�,i����Ve&z{(��������:�ǫp�0��3Dz�~p2[��aF 0��x��_捦iʨ��'��%o�Ϊ������h0��҉ت��_����~]�N/9,3Bc�q�=~�'��eWi�t���-G,�^���󎘝��(��Q����[�\�%�����T�H�V��oL�g�z�����6�uޤ��mD �X��[�z|>Z%Oxw3����oT��,�
r��\C��q�:�-6�ED�ն�3��}%uO��y9}{y�^/�[9���� ���\92�Z�ƶ@�M�a����K�͹& �չn̸��^�I8��"i���ה���34�!�A@ �Ί�
��(���G/y����gX��5S�`����|�O�r�&�1	�t�Ni_�f���:쪋^iO�{V��_�����L⤶�-CO\��5ܠA�)�I]�4���ԻV��S��,"�^�C�s&�W����F�ii�t���|�[w���E����7EHq�}��n�蝄���Q�{�X�x߁	������G�����*�f3��sV���"6�2��~H������z���dq�
�c�f�����_#42Q*Q�� sw8r�jP�V�e�E���L=R�����2|�%�����y�c��LD�#�����1� ����f�����U���?qy�Y�2"֭�+%�Y
��ۗ[����t���M6����_K���Rs�	;���K?�
� �^�^���@0�'�:�S���7W~<� -��Xb�����Z籑�3�*r���o,E�^T_���NR3++J�>st����B��AD� ���'�tS��"&�����a������t�*���ɬ�rVq�����l�A�-qn:��=�O�}�p���X��'�o~�� ���j�"Dr��b?az<�Z7�|W�}? W9|s͹�BJ�˧tm�8w�[�u8@TA���z�w�#"�r�C=
�g��ArS����s�d~'(��{Kޛ�p���'11��gE�NO�Z�R��E���{�N���4tOQ�uY�+kZ̉��^���E2�����F��M\��鲼����"Q���`b峣:V�>������qI��i��ڰe�c���������n�/�o����Lv��xYN��������?CK�v@�_��b���"��$c9��ɚ�����[?4���� �]#!ݍRO@&�t� �RR�"9�F#H�������ޟ��v�s_�}]����7�����%�Jx���Ò�
|RJ�Eu�[���t�~/G���z��뎹�oo��>�x���F�4���`�<��~�)�2DA*7�:��bf�tR&��6�<\u���J���S���#�Hy�f`Jׂ(QM�o��r-���(����������y{A���#�Q�.b8�`�����Ax��$����(�����f� (݋z�.��`�-~עZ�m���o0���6���O)����ׄ�A'���##k_���|3�8bT4�t֟����{��1/�ӋYR�<���tp�����k��3�Dڵ�n���/��Gn���"�,��/�`M\W�$�>ce�:���;L��^��Wt��PY�s��?*q؃��ӷq)�=�U���ц��F���[��E��"7c>	�=�¡��O`��G��"S9��>����D���z�ݧL���-��[N��\S$��Ok":���̳�Ź�7"̍��D-~��t_A�������L�<���c�� ��gY^jv���so$#yз؄n��ޖL�����h� H�oL?`񽨵���8������ɥ��e�~eAZ7mR�JK~tZ�Vt�O�2L�yǯ��-J_�����o�>'�:v���[��nmU�V� xإ�W��r+i0��Y]D�u9ȣ�7N�P�{1�#�@��`���X\��e��s�'���/���:��IO��&�gX�7Ƣ�4�r��sT.���QF��z�y��iyKy�� =�������)�0����P�`��+l��֣d�A��nԘT
��[7)�-b#������)I]��|n��t".���-ذ8@��@���c���r��>��͉��"9�t3Xd���E2Z;���@�.���%��=���� �����3%�6�ҒV8&U�O�y���u�x���c&�~�W����M���]��L�X�nՊ�>�y���6����DZes�"����b
+�P(�w�k,I��ҥi��c���j�d"�X���m�XO����Є�D����y����U���KF�C�d2�{F�S�x�c�V���!;8����<��� ��9
g��D�Wl!�� ����k�kk���"џ�m��݇cQ̯�m� m9+sl�?�V���<Z�-�+1�_@��d�ݞ�^\����1��:��������|4>���!�s�Z�ۛ��E/�w�m�g=+�ᣞ���Q�t���E�G����U�l����o�8�o�ҷ��� �G����I���Q�-^���618[s�U����n�,	��I�~�9ȳ��{�	QW���
e��Gp�T_w>XGQ����"�"�fzGE<���y����ȭg���٢��M;CK���8�i1�v�qwǦbvTb����	�8#'�[��I���1�H�G8�8��-M��:��\�J��T���q:�.Z�F���Æ?Bȓ��L���@�7zޜ�t&�~���I�=��&�_,F�Du.���-@̀"��χ㯴�_���׽d�\>�$����M�W��S�w�a�P�����2!{�dIm���<�(��zZM����)]�73p�kú#/q���U�־!����0�@e��u��`�2O�'X�p��͂i�0ɽ�6!G�uo)�tֽ?]'���,�9yG������[��3�]��OYb �5b�X�E<zTi��-�@8-�]+6�Y�0��f����#�ڹ�ޛ�S۔3/T���� P���O�T����
�<�8�n����<�2�b*5����H'�x������
�n|��gγ/��_&Շ��t(]1��F� �X���o�v�
7�M_��c��7|(�ܟ:��	�b�}���C?u����0qJ:���{\?�{�z�q�ͫ�ÜK�E���C1P�ts��*ʈ��骾��Lx���ʁ=Y�������!����Wɫ�����~�q���"���������'�ﴻ:�ƯT&>^�����
��id��&������T*�����1��P�f���7�e�{�O�����7떴G�͙#�1Qjw�Y��e�y�l�'tn�6_M�gz��}�9�jV�i�V�~2��Y�$#���~-G$���@�|�a!�Y?�#6ϲ�r��;�t�D��E��^7�z��p�.gT�SP>���H�JvV�Gt�o���R���$�v)M�0�}�E�հ���!� 1�r����F�"/\�<:��0���@�jR�����C2�, .ð��������|=H�|7�z.�/�y�%��  E�z�ކ9j)�����덫6�.��giR��+��cU9�i=��.�p�S��祊=�	�y�R�;N���w}dv�y4�H�{�^y؁����Π�������e�k���	������e����2l��Z
R\�|�Pj�ן�$B����@K��� 	�s��X3�AQ���c�m ���ݭ��b*k��PY���t"�M�J+>��S˵1İ�SK��,'YϨ�
w�d���o�W�Xf-��{�J��+~�Q�;]��p֑��O�͇���=�GJ����u	#\o�?X\nMh�a�I�G�wrW��t�9k������H<^)�@�����=��O��	QqQzіյ"A�BY�pB�9��5������#���ɕK���aU���$.SXc�����ob.��&�e,t�O5E��E#,:/�W�(c���u�G�F0}��{c�XN����R?ǋn����2�?X�ca9�XU�PLB�Q�;�e?�1%�Rp3�^\Q,]D9�y��D��_�a�B�H�����-
F�=,��ӵy��t�q)�ޒ�1��u��B�ґg�#�=a)�rӻ���	F�Ԕ��"�k+UE�h��ǽk�{\E"-Kf�=���a#`n%����ք#��w57w�����/"DӼE���ɧ�G�KȂ��1t}�'H��(`�g;�_�xN����~^D��ۤm�Ks��~~3J���,����$y�A�y	�t�d*0�<��&j-�;�/����A9�����z7�1[�\y�Pfl�y�/�[�y���8OTʍc,ݢ��#�\O1�O���:�{} �{CΫٵ�.�iU�h��8�j�nEA�)�m4�h���R�<�yb���s�R���ZUC��a1J���\ oj`J�Y׍��2 �D|�4T6'��'�(��E[�-�_�E��Ţ�� #�"v����p䆈r=��� �K�X�x��;�H���ۇξ�D�?�mʕ\5S��Mmp1�}��S�����Q�8��&��:v���p0q�2!?�T 2x�#ʩ������H�(���"�npN�k%���Ņ��U��� K�Ry���n`qq�zI��+q�VQ��̹dg�~����/�p<R5������k�&�[՘��S�P����V:��e����r |b�F�ES��8P�0�+��:�\�=��!�Kb1V��� 2�u����Bh�	�q9�f��o<[ik�*H��<]�����'��.��)�cog���Nr&{�.�����|#����v�q�uTy}y��t?�=��wѿk�T9�\�|�а����:��������>��M�v��K��`Nlh��~1������G\Q��y���V�� �Ȯm�7�ߜU��{�&6N�2��aS٣Lj[GY��E)NS���,�lZP�N6�)xZ�1'(��[]� �BQ��h-��J<�q����>kh4<s���	��s�T8�ݳ*<&N��b��bA�l��EUQ<�#y[����=���m
.�i̥�,�۠n�*��vF�Qv��+�(���_YJ�iYi�}8���l1"L)q^)��}N���k�
?�=����qy��[۵+p���_-2;��|�G?մ���=��ʾ{�J/&��w��s��*?�0a|����ۺ�>�'��X�d��a�8���]�H��-7<�?mM�6 �*x��m���=Roʥ��~ ����_Vj�F��Vw)'�"�tUFz֣��4�'O/4�S/Ը��y�{��Qꞔ����4nh.s�H��?<���HH7�Q�k��s����Ndi�H{�(�vc��͑�a����*.���h����<�r�9�s�#�ܦ�8���x�\ k�B(,�J���'�UU���U��r�	[����2�p�{��.m���Jְu��t�Đ������h���ݏ��ݬ��
���ba�I�ڻ�6
�e��P8ò��1��E
ǘ������o�3������/H�[�S�Oy=������0H,�!ot����]ۡ#|�%��z����tIgT�8��˽r�����⫞�%�G_��򀓅�ۄZi�w��^ZD����~���G�t�)؅&�J��x!|�A��=�Й���5�q��>�5��.^:ڃ�Q�©���T^�К�7_0S��]*��M��Ni��[f\",��h�6�/�K���[�dI�P:/��(����&Nk {6��{���d�fm�霫Gp\�H����������~���[<˙=ӓ��{�6G�b�Iy��~uI�#�Y�V�f��e��/P��Z��'���W[$Y�UOqo9Z����X���X�G
������v��`70�k�:(�!~��9���I2�p�T��u�̣I�r[�uR�km<�|���-<��Zߛ�H\��'�Ů�C�%Z�z\Ip#=����+��Q���uJK�Q/H=�]z��ƢhA�r2��f&�#0���8�TI��t��F,�m�1���]FwN1_�s�h���S���.zz�gE�C0gG5'�MpV K�H�e{H���,8�Ԛ���7Fl
�ն����o.�'3��J(�˓�}��,���?]�m.�Ң0����7��H�0��c��}�n��G�]�3Yr�Յ���QK���ߑ&�d=Řъ�?�_��/�^���\6��*W�i?o5��R���x<���p{(�Hf�c�;��8�}�+{��S�?e�s�0)���
w�������Io�����,�ZƗ�KF�q9��5��z��t�sW��`y*X�$�&�՟�����|���7��u5���qp�:a��)n�'��+��O�'*�RN		>^�3╨��1uF.����b�?��UU kP6�R�����s2?�J�G/ 7=א
X�����.s��<�
����ˠnS�Y,��x���r�g����J��R�2��$�!�O?�U+��q5�^�������H;#m'*���#�m��1�0L��J�xV��r��Tz-�WS���ƂS�
.>�Q���d�5O���:�؟-�S�n}�OUkL�8�C���F��(<艭�ϒF�����fF�m�P�E�H)
́�Zu���(ۚV��Y%E��Y�1�;KĨGEz�8X���#ؔ�H@M�3�蝇[��lgV�u/U#�1�W�oHHԜNp8Š�y5����J�Ů%�����4@�f*���:;΁�c��ig�����}�
�����%�f��3��ٰ���Q�OM�:n�A����e�����Ӯ+!JB ���o�c�o�D�J��㎬�"����^{���Sz��͙UM���Wܶ��~X��\��$�f���ins-�d$\����m�Tu�wQA���~��sC[�P����OQ�7�b�%�M�h�@���ޫ�Үz[*�m������&���SKz� ��H���*<8Q�0>.K���h�H,f���K4N�M��7Bb�5�ڳv��W'�.�f�G��e�r��أ��ՏV8�S�������6�ϯ������!X���[-E&�R�����uDw~���?��ߠ�&��h�,]���an�"Ku6w����܃���ę&���T���)�s��˚��d��om_}߬��;?5(6�W��.?'�Q��X��6g�R��K�
�3#Xb�F�z�$��{+]7ԅGz
(D���cJkm�6eNw�Tu�ps�E��v�f�НFc����H����a�,���l;����$P|��"1�O7��!2/�ҋ3���>�D(7�MovI�^��N�d~(�-6�3�M:҈�hT�h�Ͻ��C�@O\�?�Mf|�n}�=����B�}C�)�M�L����e��?�w�)�y��G�^U/;��T�$�~�@���Vp�j^ 3�q(�Wх�kL��L��B�~3���wʀ�GN���ٴ4��"iFsh]���u���l`O_�mC�C��_X��Yy��׮�v�a(ɪ�vO]z-@��5���"���Ѝ�~�
�����HR�:�e�����Y�b�Y�tx��o�LH=�=��|�߱~-���pCq�`��?^����ٴ��nT=q�m���%OK8��{x��Z�=Dk�o���BKa���5����c�<��:#�5�vpr�hi?�lktw�ի�������!���2�ԝ�����£��U��9R� u���4*Qg�p���x�(HՑx�� ���3B'	ؼ�H���!��ݛӼ�6<��	ԯ��`��b	�?r\��b��vd�	���ˀ}�ՎT��ڃ�\�� �Y��s��fK�W��[h<�oV��ڱI����^�"����W!o�mu��!��]۱���DqxDp�£�ۅ�a��"�96�V&	¢iˑ�+
` W�I�[+*���<��Nh������h��(�f�?���H��Zj��C���<y�^šP��پ	�4㍪Ћ���x�Y_ը�p;ȊǡsҟKK�@���|�4��7uř�6*uBs�S/���1��{�}*�T���0�p���r�<�'��V%�?�_I>�sF�>��]�w�|3>����D�(��xw7�rW"W��]N��1ж�|އs��D=$p��ả�� �Oi.�Z�8�gN�"���ZQqi���M��ѝ��b_ŵ۩�nx��6Oxx~�d�@��~R���6��@ۻ_;�Rƙ�2�OB�i4׀�,��ޕ������XT؝���������mv�)v��hn6
�A����öA�[>�si��=���r�m�B�mi��<ٰ��^'��ɻ'��ӊY��G&�J�� ��B{�P巂�g}xGi���]u���Etz�E΃�@���������:�%��L���G��Z�I�|_�����j+x�3��7����5�~�2�
:X(��JS��\�<zt8''�wM�9�q��>�й<�ܢ�u2�z����Yo׳iԵ]��H��Ne�=,�G�Ȃs �߮�'�k�ww�j�6(�Ɋ��Wl���[ù_��k�M���J�&O����FM�"��JJv�j���� V�aj�gV(��Φ����0�y9�,���v���mÎ�q���Ef3�����"��Z���)x�`�3t�������5���R�%JT.p7^^`Q�������D�w����^�Ɉ�T|�� {h�j���� Ѷ
�Ԣx
p��#%��X,�u��6ha/h��E�cigb��/�0�,�8�O��ӎ�r8�!���OFT׃oE��d(�j��>=7��~��o��v/*_X	�Yy4����fL����؜?�ܰ�{�p6anJ\�g�����Wd��8y��}�%>?�!ֆ%�����1��V#�i^y�5b��q�� �S�q��b[%^�>gĔr.{�S��-�v4s_��q
c���<��X�}�J��5e~��Ef��� ��}�iv+��f:FG��u?��Nd9�	��lT�M����/��C�ޅͮq�ML�ڵ��Qe�1W����8���zԻBj��6�����7�P��ט4�3!� 'ʧ��aո��3f���	k!�Z�"1t.��+��O�����W<(Z��quI�ْ�4�zB�m�&#&\���@CU].��1���U���C�WI5��5�3�]�vo�aK�ÙOi����<��[�b\����U�х)����t[	���@������)����(��D(����?��Q���y/�J��i�=��r�6�Zt�'}�WtsUL�/Ӟ�^�q>.8ϥj�R��8:���B�R��cS�G�E�kl��;o�&o�IlX�t&T�#�7r�!�ưsNrttά%�#Gn%���H��|>f��Z��Y�&��o��.���R�����6P�d�A�� �����{{}L^�DT{Qrz��)�0�5s�w5u�����KL�E�G����-��F�+�l���Xk�ϰ��Os��N�K @��+~^����Cό��"l�@��	mkk�\&M�y~��r�x�Q �Z��8�U�>ǐ�bc	�����������r��4yP��h�1�!H��e`��$�l�>4�]j�n[�!B>�6�Q�8+;�PMX������W����Ie�`.U<��M�k+�ԃ,/H���s�P;�P#3���k���1���80��q���Ο:��z�o$�!�F�;�}}B_KJW<�S|�hK�����cj�:L��6�ٙ���A����Pz��^)�a��ŀ�ᣠ��� cZóڼsLV� ?`-�DT�K�xl�"x�ǿ֛�iB��7kycy:���.�lW�ʺ,����&z��0?V���/C[Z�n���F��r�xag�*��٨̶��Ú�H���N��]F���	G��k?�y�5�d������͍wY�Gh�ȏn/�Z�`��:4CnYK���*�jWg�hXabTR���vߎZ��瑐@��p�k���ux�s��Rw�v�� 0�P
�O�H�D��ƙ]�����x�����g��MI�3q�>޴��#!'Wyt<`����?D[�1���tě:ԝ��Ȭ7�=;��-�"ѩ$!��TOZ��]�>�m��@:#�{�^4�nƌ[�l�s%�ǃ&d>J�[�4.{��1�ΧK,+�>�Ud�9���1+@����-��ƾ/�xxy�nz�Oׂ	i4N�F�Н���B���h�����i��	���k�)��*S�{>w?j�H;�zU��������m�'�O	�<�s��X��%K1O
��ɴ��	�ݎ�����A�T�ې����@�'E�{��ɸ����Rm^��^/��M��J��j~w�/��F��P��N�����z�0Ƨh?AlJPW���I�S}����M���Գ�y~i4&�&��@Vر�l��z��n�R�
}^��b�2�iK��]
�( ��t��N�8h�g0��p�i5�NtV[ûeK��b� ����%~���b��I���8���c���vTЇ�0('j�ё��:8Q�T!��0g�u�k�|M[�=�i���~S?�U�\���x���8�*�.a�{�x)1�C׍��%�#����]0a��7�-��B��hֆӪ�0�ճu�q��vB��T��R�m��Ĵ%G��&�9�s:��Y�-s��i���!�,ٽ���x�F@I:��[Nݶ>!8&����P��C��1��=ص�+�r>N�����B��ky�]yQ�y��ɐم�t�چ��Y�_�^]/gvv�]�	�P�l�Լ�K:}���t���;1��������}lm�j *�|��s���e�*�����t��Yթ����u�lcT�y��&�Xhf��9�����"�uJ��HiaP����Z{�X�dT�^�vz
1��O�;5��D[\�_��V�I��cu��d������ⰻ���M�
utI\0N<aX�q��h
����hTs;�*j$��a�!�����wP���ʲ�Gw*���4��&�X�S�I�r����)������`0��� �6����G6�1�Ͷ�B-�W�BA���pM��$�ȋ�1!�/%�+�����\4<s˦�]��t��˖:6B�p7����u�^J��Jj/���<�����гҼ�ǭ�)"_�Vl��k�SW�Sx�p{nu
[T�^��/ú�_ڗU��r��ɿߖT�_�.�U�G��0�c��Ky߄�ٓ��ø ��4��b���ǐ�{8����
X��U��fq��AwFG�k��t�����gy�cWaFt��� ѨCj�.�5�FO��C{���G���SmQSMV]�X��$|��=�e	�Uh���=�47�X�(�P_�,��7����f�u���_�e&��5�y�F�<���Vk�q����VW��Y����Қ����b&�:��I?g�p�K=UU��B]��83��6�=�4(�8���/5!��h͸S�g�T0�L��Ea`�[Y���=rk����PQi�G$�W)3SSb+Q��Y)����ߨ�}h�W�Ȯ�^�D[JG�X��uK\v���Og��0H����)8r�-&�9�$�:����ǡ�~R$RrDBb
��ē�?���RV�{p
�}sF9M�0��HƘ8O�5��n��c����@��D�M�wQ�W��+�P�'kL@��?�UBKd�q�ůa����z�k߽�$� �ѧ@%3�ű�p���
��;�$Y(>sE�_�mӏ���}�s�I�Ѡ���L3��P��Y��ӷ�K�i����nl�&鞧�Q[M^^�(��v��L���S�]y!�����c*9��k��SOҸi����-3b8kףE�zʭ�#]��	䙁�w�l����k
����B�zp�$�|k�s�窡%3Hb�C�3ʌT���s����7ɭ��K
�jzyt��	1���y�m�"7(�:��Nڪ�0@�"�^|�pF"Ңl3�O�S�J�]ܧb!Pv��;)g4���4�=��{X���]���*.�����R%_�N�]�h�q:D���D�m���O.X�	��S���3�X���q��:�m;�k]f=Hd$�T�~�(�oT~���qX�D\�oA�B����O�$��6v�����F��֪����,�	AR?�û�ڴ�����T; �IB�O���Ŵ�jl�I' 4"�C,�{f{4�X�h#>�l��L��O�X��#ۼ8k?  �,LZ[H[���j�+���R��~<{�G��3p� Wr?�L$��M1�v_�UXE���`�O��흒����"5�y��l�P\�vo����y{���A&~6�^s����}�#I�OY��{�6�����m�h�i���3MY�����4M+�I�Ƹ��J�X�g����o;��������������hW�� 堞�B鈜	�?����j<��W�-��_��Q�������?���"�������eG`���|?���Esm����ˉ�հ�z����X��ްQ���8oY�PG� w�b@�	�C�>J�xFͥ�1�RQ����*_��9�/m>}���,���ƞC�
�!i��}�;�V5�\���M��Uŉ��VV7;���'���c�7|��(?����~O��w`�뉠i���f~�w�DO,o�>��v$�H�(|t����z�r�[�d��V�$:gb�Q��3��; �gN~�8�ږ�Fd��0�t�{�G?���[��n��z�^�ɒh��.䃱WM��Jt�nş�Yzˌ�nK��_f�M���AM��=���g}w~?��γ�]���ťF���ِ#L߽)��d��}��7�!��`=�}�!�)x���`�1����m��j��U�z�k��i̗s�_�պ#���6�N����(����o��%3���uȕʽ����4�9�G6��?���FI{Z�
4�����$ l�W��3!�'�$S<�(�2v��1[j���|
<bC?�yF_�ĳGc���=3@��a��(�iV�d�O�����n٘��(	�+S�h�u��`L�7�k�-�`�-U����8�D�>�P}-
�Ml�v��Alj�o�f�FJ_����U\��?1�c5�K�@K)�+�O���}l��
Y�[ޞsTb�aX1H����J+����,������f&������	Oc��&�߈�����H�j���v`�gU��r_��Y �Y銀4GM���RB����
@Pbr!Z���g��v�}�|XSN�}�
뫷0l1ˡ_5c���Y86�#.f������w�"f�?��-��Jd(��e�*V/�ဒ���O�Հ�R��o�˲^7w���NdSU�c�i���������uu��f����[{c�*�O^�R�t���s��V�!�*��B�<BP���f;�U��^J@�����^So�AR��ڣ����)ա�d4��z����� ��In7�㣻��Αɚ۰ʬ���w͹������	<����F�������~�{=a���#��l�C-R���>@�\;�ɶfE0����}��j�ڿD���we�{�Ӂ����u������B{9�ѣ����{��R����l���{�编z'���7�P��:�im�nE��=`~4rc)��ؤ"�����,�Z��+��~���/�i���"���KW4��<�B8�G��_��Hm�_�|'u��n��ڬ>xW�q�����s���0%�[��+>���*?�|�V q�Oԙe��:���Xn�Z� �?���x�VG����m��L���2�%����/���R�} �I��w�1�����Q�M|	g���ɅZ��^��ڙv��Q|$h��%|6��I=��9xx�U���(TB�`�R��7d��_���P����p��J1�/�`1�)�YK��즀:�}�7p����m�tB(��������܁d56��3+r�Ӻ�خ:�[f�c�E���=a�&-� �4�P|�`���<��?+��S��5���ûx/0�[�"���_��5(xz�SR�Yh�n��sJzE����޾'I�����Ǚb��2D֫r1�ua
��Wr�����R쯔��8�?��3y��,׋���%��֦��R!�o�����,co^�q�����q���EB9���ο��b/4R�ïl�z�yB��}n;�3,I+��Wy�-�'��ڝ%;��Ai%ؕ�Ջj*��%����fG5��0�O;�:���|Kߚ�-�a���ff:Ҥ�"�pCX�Y��A`�^p-At������p��z�������T9��@�#��L�����o��E�{Dd�X@�y������đ��asJdK^�����۾���i�I���aXN�S���8��|q<v>��PU� v��.]�C�qYO��E��(�D���n�㴖D2���d����]��^�����ţ��.�ح�T�OaFS�b����x�1�8�i���4UM`��m��H���?{�;vk!�kq�q�q���{ή�{IyP`��uȶΓj<�~aos��>�d7��[r��r�Y�?�a�s��rAjf��[� y�yo�]A�d{x8~�l3�ONE;2~HR���֘����K9��;��T��{=��B��Y�.�ؗ����!�\cc�.�o&�^���m=��o�rC�&	���Rj�a]�tD��Q~���\�,օ5M`����"���.W1$C�0m�E�V��ޗk��p��Vy���u3vx�"���p�y�g=a�g�1T'��2#�u�z9�vP���!7�ʤ�*B���X�F���9�$��6�=Yp����{:�#KEk3��y[���K��C"&�sm?��\�]F�!��~�m����JY��s6��m�+:o
�͑���ƃ�O뾩�:�8�0�>"��u �˨���QW�'����&��k��i~�EOv䐧%1�t������=���N�I6�*��=�cf��nN���k� ��9�~��Q!/}���Ï�]̑��z���rr}gHX�E�9�=հ�n���/3LK�Hd��^�{��}ז�)��I]ԾU�K��2VΖ����[��ܪ��Ԋ>n�s�j�tA�(�CD�0qS��B�U2ɜ�_!~U3�p��}=.&���`}���p���M��ঠx>������Q[F�>�FFv��/;ٚ�e�3�ʍ�y�H�볢��I��i�׮� ��ޯ��=�ۤ*���"-7�k˞eZ<ʶDyp&������?_;DI��u:J��o��l��Z�1H��NM��"Aw�؄�����w��:����D�*3(�?����T)�XOTƯ��2>p���-�R;����`��o1�z����i��;� ��[�w�_��"�X�'�}K23�v�eC�HE�ܷĶ	eG���|����Z��:���ќap&d��1���Լ��i�q�Dpp��W[�͚��5��yf�����[��~5O��(%v�Gv��EW���p*8o��s��
���fW�TI�~[J�\'Z��Ě��p�m���NN�|U@V��K�H��g�a7��')�o�A�궓�\6^9��.Ҟ�Ϲ�"�jD,�y$�H7��8.�e� �\AbA����Z@B�ۥzV$�*�� o���b����j�1{�u��J��g�_��}I'<�}�����V�̈́�6�?�gCQ���w�˰�i��%d�d+��|L�C��6c�3�?dy��x�x��:�����J?�qժLj�`ܭq/��������雂�m��5���8��f�C��@J�KG�sL��}|GV �ۧ�oD�x�U�^J~Oc�`e,Qʀ+(��q�������N�����ӎ�pO8˼��[��v]Wu��>
>V%Gʛ��\�h�/Q�n�L�˴���w��oC��z��DI+����\�~����v���*�;�ܝ4S�e.U;�|�m�Ta���y��x�ag~-&I/뛪.�W@	%�'��Ҏ��$�P=�j7�RQ۬KFۆ��i��_�Y�]�\�0)~����Ak�"���)��P~�ڞ�z�m ��Bp���|�9��s�D]�~����'�X~�U?zD$��� �+�b�&;���Z?�Ƚ���iG�Q{x&7���s����X,{���]CT�c��k�J� 2�V���ҋ�i�)��9%�s� ����S_%v��D?}��e4v!X�-��b�4���%�e������^w�}��V9[��[��Q�-~H�ۖɸ"�6U��K?���'�:��s��+/���O�yP�E;[�y��S@�f�ڧ��s�:�+��y�F��	G�X�����%i�Ŷ�ְ�\��?�$�[�d�L-�3��:���h�^`a�$B[�Dc�����z8
�8�,`����I�����^�Sl�g�F�u�������\�I3u��_��=
$�|�"g����U3!{��]qEZ�I�$�h�w~�u�=U�JQ@Əת1&�>O��<��Z>\��Mq��F�A���}O�͍��tܣRa�\��wdW�?p��4����ӯʦ9�LUGӮH�_����&��<���E ;�Z�����r�� SY;����ۅ��B��!Ő�t��UŖį-�[��8���>{������H���BO�XR �%m�&�%%��T$�՗����i<6�.5~���f��BG3֝�BM>���qk2@��d��{ �n���a�c��+����X踙_f����$�Fu�����I�Z%��#��anevo���l�������o�A�W2a�.`��Hzmؚ�5�7��ƎV�ֻ\���PO�Η�DC�����ń4�CT?ϫW��/��|p1���M=�g�"�Y���-���:����x���=ӗ����������!��7�UKLI�d�?,�$�n�E�]�������������D��c��y.Ȋc4u��E���l��˯Ro���9�r��-A���ηڭ��8}]�=�]8�����i� w|Մ��Q\=�e<��۫~��"��6�e��]8�(�薑z�%G_7�WR�PC�Lg�F�c%G����j��w9`~�0I!Kr���A����\���(s�B/��2���c((�0�C��؅�3���|L7�9�sf��P?$�޼A�2ٵ�E���x���5�k��E��
�V����&�����K�@�fB�����@7}7v���b�[���')��̞��r���Ҟ�� 4	D9��g��8D]��t{�&	YXUI|����XB��E�>�h�"IH�#�5��D�="O��tX��Y렶����C��Z���!g�#�Ǽ~49�Uj��"�q�X��'����+�5��/B�A�\��`��N)�a��}���Z��IG�����a��"2�}��)c�KMT�#v��fZ�x�X�T��o(j�B�J�ޥ�ױ\�*'��\�s���D�L"<�L%_��w4x���}�~(�R�弩L�W�-1�o��[�ϧ��^���1��,Jr��mV6�t�AE+D1J���7�LQ#���.�!)�*8���P(���z<a�M\Od�	���zƧ��·�˩����-����A���D��n�wf.��vӌ��9�h��2�}G�{vVs@u?�[����U)�Lac ���)�+0%���盟N}�]G<��` ��Au4�1)2~��� ��nJep�����KjG$�|��1�½��[f�� BcQ_�����m��I��M��}��*-scEӍ��[S�,tl(��� �t;����2������o3v�bo9���r�L3��u˚�o1��0������Z���%n���y��Ʃu�R<�~a�
� !��՘x>�#� �j���J"yw x�	��s�H�W��0/ؤE���|JԵ�����3�·p�0ݳ��^p�x&��Gf�ob=�s|��pp��1y%�!��(�@����f��ۤ�pa]�FS���8�ؓT�ޒ�?Ny����Ѯ~O�HM���O��B����#��~�9����������*e��MV��Qf"Bee�B���T�W(#+;�g���Ν���w��η>?� ���^��x�_��#�S�fZ��1�>'�9��I��[e����2�y�'�'��14��i����-�w i���٘!�/�HbƓ�2�h���Z��b��ǅ<� [�9��n[�}�fU��K}5������+9�4��dY+*[\�*�t9�Z���c��f����4��9����W8����2�@d|��k�1b7���.ȳN���γ;W�\���t�+�U�9]ϥ��Z5�.��~�oi��O��'[S��mD;r�;�{���(L�е/�4�%]�AWUXf�m��Z��]L՞��-�`�[��;���w�!o4��-��v�j.�D�k�:��W��Z��~�4�����bj��'���G���z��p�,��ţ<�Q��:�~�PF���s����c���˟��b��7�1�	PP���6�7qG_GO�Z���}.���[�OJ3!�DE˧��+�PM��.{=���6*�i©�s�mq���I+�?��C;�ǄU�.X�SR ��h�cm0��tPq�ؤ����sܶ������|hЭ�oȭ�H�����O�ņg|�0���̀|�����{����!��X��X"�.r�o�ʹtz��U�:��r�8F������Hw�iH�w��Aq+d�=���=����&fv]�'	��󄡹�&�V�DF!��d���5�w��[f�M��G��ܓj������}�����A�r��R�໦)Z0�Vg�5�c5#v~g>V�ck}k�rQ�5���B6�� A�6lq�	!�o�q�����\�I�,��ꁩ����@V6��k�u�a�������d6��I����8�5��z��==�d�Á}=����	Sv��MN�L�W��>ު�r�5ִ�3�~����\$&u&�<�\�*�Rv�?~y���}z���t~���;<d��iҼ	x�y�>0���\;IO�m�g��!��>���1,�h�x�<R�!ޑF/ϳ{\�ῧ�P)������gQ�N�`��ל���g�*�������bI�^��=���uװKҌ*��㍮˕�C�6�SV���q/����uv�z��x���Te,��b6���$��EB�j�K��d�"�'�n�{�����C���M�$Z���-�eA�cS^\�5ʏ���w٨�\Rw]%�O���럮�G{}����>�)����Fޞ3I�o��O��=2�s�\�zCS}�� �Y�@�m%���hM��J߀�$����^��i]�Ū�*�]p:[��-�e�y�H/��G	*��A���ݜ�y�ٿ8���X�?l&����6$#��(.��?�)����;B[}��{T ��xQ9�CD	�Qh6�=�zi��;�[!&6�1k�Og��Gӹ���P��U:��ob��hZ?��*��P�]��߲w�:��U������+��<\�7��5�ڝ;��{��r>�%��'T$,����ʊ��j�dp>�r�X�ڟJ��b�0o�y��WB�#�s0���,#%����b��S��"Z��
n�2����oL��a�93h�ʯ��ov��>���)�(��/J~�� ?3������yf
ꗠ?�T���-~0�9�y[����w�f�����p�
y�C��=xO��\�*޵�@��@��2u��-���D\����o\��Λ�]�H����D���,�p���_�^��H�°�kh�=|_��,��T��<�☰���pg�Elp	�
TY�`�h�}�毤��D%8��O����W��_��VZ��|C�.u�ޫ���os� ,j1q�-8g��
���"{u2����`u�Q]�=�QH�zE�5_Ry�|I�ِ.��-ّ$7n����Ю�v���!uBGdDY�ɹ����l��͝05�%
u@b�����SO2�Q�,�jJř>����c%��.�*@�5�����q��)IU�kРw�򕜍�O4���ݎ��.�֫v�A��-�=�}�e����N�Ų���(E�2�)%�}���PC�����<�۶fV���[i'7�E�4��]���X���ʬ[C�^=��*)��b��K}��o_H�q����Le����VvWT�v�J�%�
'��IG�Y6�L#�|���!�̓+�߲~�7�{�dI�fTz�P�X�_>��>z]��ԕ�S�5z����Ce������r�Zv�5��y�S��?�K�'�8�S^��I��o*��)��{xS $�J�H�A(;m�YL
���ZG9�h��\/J��s2^7�0�h!X�ƭ����m��fe9���G��vW����=k#c�kw�Q`�v���Y&��=V[xj�E�2�\�1_�|�s}D7�����zo0���]����C����=�F�-�zH�Ç����j������j��e��9�$����̖c|{��ڿ �*P��-�]������f����dɂP��3K�LX]o����p�ߖ9'fw8s�nJ�%����>�s�A��S{wn�y'������ �O'��2&!���e�0E�e��l�D�k%H�9��r�XBب2<� ��j�Voj��>*���]<j��;��Xљ�8x90�-�	-��@�U3�]Ky>	��q��#�:o���qS�� ����\x����Q��p��p�5���)`&���pE��a�n����;/M���U�E�.�O 钉��I�G���O˽��·���<�am��|���#M�%�P�q?��x�9"c&v�<�\0�O��y������-���S�gR%�1�J9\˺����H����VJ�� |���������kN��e��^X,��v�>�B�ր���Fƈ\6Jә�&��<���7�8j�����0��u�v�-�����{��"�؍}*�vK���n����3>�V�h�
V8��yI���7!+�"��Ѹ��4�7�Q�&^�g)�6Ƈs}�lR�7�qUr2�	����x&7����/�Y�����'ȇ�{�-g��\��=� 1}}Y�>������R��Zָ���ޥ+|�<]��nB4""��d�Tt��=jٸB5�����l�R eI2��^K17��$����CIDwޛ�R��J�����֭\4�����ޘ��"�7h��ㇷ����D_cy�t1��QO��%�_��3���+k]��uOs�9��Q���H�5ĕ��$�Q��-��ᡍj�?(��@s�X��UT��g���!]����x���Z}m�#��
�����4|��I�]�-�PN���qG��"P#d����]G����y+k�Ȭ���λj{��
���giC�W��nu�������hcEF�~�xx��@r���b��5�/X�-���~�T���`@�Ѝ���*��[?JB9����*���?F}*�����ܽ�Ƒ�\#4^a����d���W��K�X7#�ѱ��<������N�����f���u��U�tC�C�B���҉�`aggS�⌮�fQ���n����V�Eu|K5 e����Y����<��S�7a����`<([�Un�r�qu��~�vo�V����K�ݑ�
z ������?�ɡU?��|?�t�up�t[�)�ī��b�d*{<��T@����3��&u+9n������Ý����%��t`'�n֚�D�����i����\Q��CJ��^�Jo�m]�<P%*���1Ac�����ԨNHu�C�ztJ���a���p�����G
��"����x�Q TI��S��Jِ�������832�_� ��t��D^����ɧ�4O]�r�B��S1d\���/�D2�<ȳH:eeN���On��5���<���]XY�&Ł��/��Om��>�?�r��B�g�4��=�4�c���@�|�.��7��**+k��zT�pt�R.d��/�����C�A~������i)_3ƥ�I��5%j��T�ډ]�V~�u���ܟ��㙖�M*2u��-9�Y�M$��#y������������>p
�(�c�.��~���L�z�C�e߇���<0�Z�wEB�-<�͓�g<�ɖ#'��eE�&���J�1�Jh$o�[a�] [���l���\��eo}#'#�A:�4������7�p�)�Ѷ��8�NS�zHe�������k/lE�^�w=+��#�J}=��K-�^9�[MIP.���4��h�!Z�#V1")]��@�0��V��/��?�eS'�r�Da.(IX����)�:�hU!ll9���)��:��S%&�f��E���	��h�trm��"B����TѦ��������u���X�е�#��+W��G��.,n�*�`�浹.P�]CN�4iǖ��L����#�����X�ؕ:v�t�/�u-�.w����j�+W8ud�ܔW���4�❋������Ȭ-l�@Ԟ��`��8�ˀ4�L��,�� �ܽ���+P�-fPo�z/�x�L	L��??��_��m���``�):^����`:�nu[|7��rڣ�u;?i���ՠ�k��06��Gp���=�e8����r�[��\"����:II�Q�l��g�#�����)��23:�tꢀ��tQ�� ����u�`F?m�"g$�o��D��Q�.�zM�G���8�L7ezg�>�X��~5kN�߅4���u�j�|U�}���֊�b��u��V��U�\,�8s��s�E�zb���~�� ���ظ
%E�7%���$����]��)	�^�U�����s���w�x�R_���Q�����Nr�GX<^Z�7K]YV�5g��������qvI"X�$KdV<�\ϸ��E��\@��y�	=�ڈe��8mP��~E��M��7Q��2]��ӟ�1��ድɨ��c�&z����r�J�~+�.� �	�	y��)���$T�u�����޾�����7K�5��9�[��~�H��Ŷu��0�J[z�����{O�=L��?-��B{���)3Q�|)�[�m�=l�f2kF?�r�)����l���ؕ���Al��D�������1� ;������D?m:ղ��Np�U�<Z�>~7
	Z�8��;�\�2)�D�6���{B��}i7ϖ��.�í2�4�^���A嫉�٫)I�)��](n7�>�]XhC �?��>��	�֙~,r�əy������<]���$L�����rx�hqA^(�{f��2�6<�%�K>�9��kڟ^�IS�}&����<M,c�yg�@�{�>��뗮\J�K���s�:��Qn=�!��`W��Ze�a|)��u1��ԕ)���7�r��ͫ�r��Hz�����:�1e�#&���٘(F��yN[E��T�m#u���
&xs�9�tS(��(�	 3(9G�X2=M��j���r��V�K��W�3?\}�٧�uճ���>�/Eo+��?r1��4a����/0�cgt�/�~�$��^}��@W���D����D��Ѣ���1�`��ݶ���J`ػ^���T����:��t�SQ����:����ͤO�T������A� ��nTx������G�ki�_�����l�;|M�ߘa, 	7N�Հ���4P=b%l����|�큮�7���;6���[6����O��{���/R-8������Dy���jVb$; �-�P�\(��J�u��˶�Nڜ$�AB\��bn�uc��߻�o�61�T���<s�]q2Qkb�+g��T0K#P!^q�����H��GÃ�u��X+?���N{��{G|u����$=����ꉒ)���������C/ ���;џ�ߐ�n��.��,߰�/�fr������E��������نC)���#���i9�S-�3#̠�LX�Ю���{�����O�4������~�AQ��
�3�š��&F���[)�[�̆@2x�T�a�i�k=>�S��c+�H�6E"��}
����}���O�*q5!������O�)��x6�I���Q� �3P��|�kĮ.�@[j���3�x�����^����V���i4��Y?N�{��}X y�e"�R�1g����0�\�[/���SD�gE�!ޮ:N�ծ{�4�0��S��M8���2�����
��3�T�'y�����˺=�Y�}���]E�:�8�苛��U߇fb�K5���M�k��s�&� !�5�n`�%W����yu��;�`gyR�Ykr����o�!��Ms�ni���g���)��ׇ_Pi�I�m�yI������sp�Ύ=�TOe	��w���h��,�޵����BwЂ��IxG(g������>�>�Jj(�n�=޶!5���or��X���[����qI��R�^��W?��@h��"6m�/�ण7ܞ�W D�د�r��!ЩqY̃����+Jw0m�FQ�1�r4���T�V�U�����s"'�5��.�%Qy':��L�~b@z�1�m�_O���|�����E/~�}��I�	gZ���d^�<�F�٬��z��b���$�=k��V .r���P�L$A/K�X:m�蚜�.��&{�a��z�n�	��^��/w���� ����p�U��g��97�לw�:�ж���lG��ԕ�J�er�5�o<�2��$��.�>9����K=�f����
�Ι��'��K����y���η{QIw�-o����Of�ҫ0X0���Qc���z(Z'9�i�0�#��3l��.��?��&n9��**��Y`5h��C03=���EK2��q'�si>����� ����1!�栴�n�3�JU/?���W����W�Қ�����,}\��,��"L1�.p�l�K��q�VkO`]��F��*�M�~���ca.�a�563QZP+d��:������j���>�a'��#���FLlq\� >n����l�H��ǯe��@�۽}8�y�*x�1u��Y�"�M`�V�7����uk�֦�6��w"W�㹊�鳿��<��}J���5�a3z,6Y��m��{����n��Vd��d�p^%�U��lr��ʄ�`^��@oALR@�R	�y���u��P�����@Ù��Pͽo���Y���O8��]�h��$��7z�(��Pd��KT������{�L�ʉ����!1��~�B*1��n��ɡ���xF��[���1�8�Z���"U����اt��NI�EXђ������ݞ�8�"��j��g_:���y��&��͇w�w#�}58�L�S�.^�����p���A��^�j���L���������1�f9 L�?�Y1i�]�UyK���J���z��g��(V9άf����@���$�"tѺ���.�G�<i�P��>v�T��x��,���-r%_�bRܧ�bGi5�������N��%����/���v/�:qЃ=�7/��pr��!*�%2�18Į���w�_C�4.�(fĵ��紵�"z�]���Jj�\�w�R��of�|���F�ԨK�U9������9�c�c����>���f�0:a�4:m�;l5E�c1}B0��p����LbAŠ���7pT~`?x�_�7���+B��J)�,2w{5�nX��  �`<hܼ�ZO��@-�d�m�U-��Kew���=ci�Ot����X����,�/�C�{|X�_B�X��b��({��/��~�վ供���_w�K����:q���b�G���Q���!����B0�B���d���l�^���c »��/r���ޯU��/]�h`�K[���<"�����^#H?��A�~�ߣm%�1Y>p���lb�dX֯rU��ԊNÄ�ao!��c_L�7�d/�ib$�z�K	��l'bZ�lgG��~����V(����bw9q���Q����ϵ����}VZ�-��H.�>�.ЄKɷ̓��ji�B�E�_���P����?�L8��}zn0KS*���1��)�q7{�,7�)�n�[�1��g4T	����q]��lJhP!s@:v	41�y���0�C���}� AX���$�H���~
9�_�F�RD 6!�]h;�9�1���aƂ0IkJN���nQ����~�_�ھ��E�m�\�i *�Ze���S�!_���4��T�}���m.qP`č���e��`��ߦ�Y�� ֵ�%��\����B��PP��a?���������s�n����_<�"l���(a��!�|��2�S�� z�`h�����y�>CZԕ���v��ug-�����#J��C	m�9����w��ÙO]�=n�n��0.�ϝ������t�[p#�WV���.�<w�ͮ[c;3Αn����N:��C�����`�Mۏ�[�!��ĉX�����b��*%�e�S�NHޓ�.���������d�����S�!�N��Y��Q/�0[�q+�^L���d�z�W��x��_Q���c�l27��nY�Ͱ.�tV�g�J���:N�.��7Zu�e�>�f�4X(��넛(7PQћ<�:�s��r��ߠ�8	�lE�M ]��ŶI�ӰM�k=�������R^�@p�`��)� �&�	�"]�lM�'P-r�T�}�B.dzws�55/��K���$g �O'�'�{J/��J���gש���M#d]���7��-��>��;�H��p|�xT*��~OV���	�%;��#w�\(6`o�6H$�˙Ͳ����		/7�Ts�=�ұ��t[���Ca8�j>)q#�s�<��{��wS��S���/�}�į�&vb]�L��e`뺬?��g8��E�"y`��}�5�?���9�(Q�����{�/�����#vA.I�q1gy��c��f^(fx~��ꔣ�O7X����p�:����C�X ����n�#�4t�Ǥv�Sre�J��lqIT%
���Q��s����w������b�y{��.���)���zT�l�8���Z��et_�'Eg�h�+��������	��2ȿdµ�6�h��Mp<$��6��<�⁖?�3��HriBǺ��<��u�K�ͳ�~
ڹ���&6�;�fN�h�p�f����`�L�8�S)��^ߺ�P�O&z�۩�ue�����E0M���oPN^�Fs�U<n�&*�����g|]������˔�S~�2a_���i�9nwL�R�	�G)?�K���NN��]k<u�a/����a����d�[|��k�{}˺�V�}?�����'J�r�V4���� ����qL�����L��IE�!�8������> �.�����#N�D݀rn��Jgd�a�.�Y�����?����j�-w���.��{�VtK����C&HkQ�-�j��P��]N\�=:��:�ҥ�}��S��� o�RaOI����%�T @���>=!��\�E�{��f��w�ޯr�ʉ�$
���%��;�KB�9���%I��H�X��]���P�47��2�Y�C�R���b���k�j"1Y�(���#�� �g��9��A"��oJ�ѥ���a�f�Y;4�gx::{i�
�>��txQV�Ю+#���2K��Hbާ�X>�O�W��]��w�� �#q$!-`RR/R9,�H�u�.���1s����z�����!�W��l���.�׻�ܪ;�حv�ձ�社*���P"l�*"��U��aǦ� ���l���^.L���M��D|�����1��ğ*�Pݢqo�/��9�0��5�G�d<�c�������*���s�k\��R}6V9r:��1���QqO�^5N���?��'�s�r\\�n�-�-g˖�B@�n�n2u�S�D{���W��n�'���=�}�C���;0���H[�{̬(��)E��,�b��}ĉ�J���
�@f\����쯄	�s�;��w��~_1�S'I�?�J���֞Y���m�X7=/�ni*6E�B�8�" �ҝ��w_
���K�i�i�
"F>�N�qmȁ�� �&��ɸZl��+��\�t[��� ������Դ��c	�t{��1x5�"���~$Z��W�x���Z:ctM��>`�h*�ݒ��ۍ_���[�	�-M�k�˗�ð�	y�ƉV�3���uYg�4��:����ςu#�8��qb���thv(��dF;�r|��i<��,��t�Z�+s7��ؽ`�����+`����*����i66\Dns3F�*��X�]Onl5��>�YJ��X*��ꒆu��͓�]$a2Q��]�L�}o��笑����W�ifb��_gM�*��=)P1w[��~�,%��SIq]C��k��\��o��ɩ��#�8 \/�O5�|���%Q�p�d�;|�0
v�=)�8/�ֺ�<%���^;�k��V	��Fn�]A��x�9���Z��Nd����sR�'���k9Si?h.�d`�@��>��'�9����/�tc���uw���},k`-}�>�B6�؛���mrǷ5���ٰ�7Ea*�93�V�{��#w�T���=��c���K�]t��@?�rL�ol  ����5#~V��j��b��6��8aܭX�t��R��VJSh��f'��NO�G7%�� |HG�ɨb���$�~����+��X�z~ו��!#�	�f�h��i�9dK6������g�� ��+ى� C��x�f��)�i����Z��V5�G�4���5���[�rWΞ����S�.��Kk���F��1�ɫ�g����_�r��$b�a�U��$I)����n_L�h��IW�`-�s�*O��X�sW�d����o��wfj;M�	��k�05����xμ��\��u��[�p�U}�C;O�n<
�\]���6y9����,�R�o4��Az�f���P���;SB��c�x���W��*nrZ���Y�+�nW���򄂎���lU6-�'�r��d,2}b��5�/��a[Z����~�eۂ��i%�������QǬ�]� ��e_Ǒ��4�Q���G&7a<�1�io��(������+A���J��m���ɨ�=��B?�V@aS�d����=��;ו�T��na˯-v.UK<H�,E�Aܤ���H��L		�+l�R�8L:�}�AU� ^�I�q뼨�v�%G���A�b�-;庫% �r�P�j�����0c�_��d{��lбS����k��-鸬��e�������:矮���ۛ.$c�`
;:D7��zM}"��2��aR�{�P)[A�h�/��ҹ<�T�_Q�0���O�͉�&w��CnRl��$C;�M�H��(<y�Zu��|(+N߽"y-�Y�y�b�6��BY� �6?�T.W���8Z���}���y������J�ƙNӿ����7<����6�6��A%�6�M�;}��Y3���Yʺڮ��*[�4!Ao}����<k���馃�G�%��x&�O��E�>G��aF���j��c!�2Z��9���O-ʧ߀e�;�Pȯ��� Gf�{˫䷔��1{U��z��iw����.�b���=:��!',:��m-KN�:����&�v���g�^���I �A9n2`U�Q�l��&;,����S`a�6VA�a�	&Y����w��I�k�v�k�ހir^4�*Ϳ���z����n`?��� 3�!��ࠬA8᨜(�2`��lǖu�e�2�����A�5�g0ɾ��iɑb^e�*Z�#�E��� �4����?=���Q����X-�g2�=�ˍg�������4�\���o
�&|B���V������	=R���@$D(;?V�����iݰ	)kY]��;m�J������Nc-l�M�c4�������q<����O/
��$U��J
MGBT�i����.��Sb�"<o�3p;��v�~mɤ�D��{u?�*���~�/G�W�����H��L%����[?K{y�>�&��`���f`Z3�W�x`���x^6d��<N\u�YJ�`�:��㛚���G{��cѤ��[3v�3lE-�YHД�%?&���`q�`wh�&����#���_#�I��L�I��Q���M|���^?������$�� B��s�,8T��$�.�O����Y&]jɖ�<���:�Q�����eSt�lw���[pz���$�}��9��n�d��E{�Z�2�
E�/��,�ea
!�%	9������$��{ż��`��S^�����?��s�,���j�HT��k���z���N�!�vf�ˠō��3�K�'��F����>���rG���`��A�v@���Ό{�h��s6�Bĝ{��\�%��ƴ�r������Av3��y�s/-D\2�q?�J�s�F)��5�|���?����ć�-ܦQ;�� ʝ
:����Ua�ej������Е	.�y^ؿ���G)iy�I����~O X	ޣļ�'&��c�Z��<&#N��,o�ގz�x�~��1 �߽�K���ki�չje�B�t$r((9�!{�}%��P�����!����z*P}��o������᜷~��6��1���En-��DG�N������7��mu��*�r�0�'�d	<[KFwśR�xp��Y�.�-4.��'cW�L2NE�{��=���qi�e��&��[zm�d�ُ|��Q��eIGB��@�J(;jƩv6щv�#@GF/��u�~�xʎ��HR���_�u�����}�S�*��ز����=m�AXW�q��R����r���A�X���h�+3`�l!{/tf�y
y3t�[�3��Ey�A�ѭ���~S �`b���T�G4E���I+�)��kx|�qj��׻���9Vd����-�U��'��V���#0z�)ԍ���:'{�z�k�o���],7��H�s��Q�oڋ:�e �Φ؛��:
9��b�h"�r�:����\��GO�OvzJ&�`�?y��x9�y�
���DG��ᡱr�Ub�HK��w��C�ւq�������� �V�<�M�n>]#��s��Uf��vNE@L'�y��6���#�I��42���&�%�5~޶�yޭ�盼#���hϽ��?h�k��O�)i�GN�
}���M�����U��7��vs�����b��LQ����:\W�`+/�"�2Qw��_�E��W�!#q�G�@�B��,aG �$���~dv�ޚ2KD D�ͩ��������S�o\�b�%�3=��s��,�ďum�.Ǯ�b����"0��\C�Y�iM�?�_�)1u7�S����ʧ�����(;������l� 4�۱T6ɶ�<����U5��zAFiN� ��^���o�j��y{�댝֔d���NM������}��;�$l0����clεࡵwe�UX�
�?����Ѐ�5�&�@֪���q`�<�]��B�|6~i$3s+rnsOR�b$�λ��B	�A��Y�v�F����5�%pO+z���'Xy�J+t�T6FG��慿8��a鲱��^D�F�,N\�8��sŕ����M�97A�=�;���o7��%w]x�,�?�:�N�64���F�wM ��M}j<:{�p4���9�b"�����V�oH�#�WNK8��8�?ʁ����Y��3;��|B��u�ְ3t�v*�
��M��f�؇���Y2\�n�2�������9|��s:�OJ�D�CZ"]ܳ�#�]��Ϋ��_�N*`���sɊ��Aq�mO����*��H�҃�������E�T����H7�#�1t������D�V�&,����B�WZ�G������Ӛ�eW�ݪ��(�q�٬ϝ�7B��
8�SME�itB�t��̯�<'Y�Qn��ò�L�-�w'vFpY��~`�o�)/|f�`����u�5�5�-�~7!�F'L/05�)�C�� ��{7;C�E%;l������.;��(�V#��I=���:h��C�������t.��5��@�-+M@�x=�٧'���'%�d	�s�M�TЉw{}oF��,�s�*6R{�[m�Y=J�������A)G�D�zW覄>�f�1f��arL�l�F �ڥ��w��4WJ� �y�-�Fw���M�g9e�N�C77V���S�y�G�%�$���]2���.�m��F�&'���]��O�m�,ѐڹ�p\���5��:+g��s����&�*�=BvF��W�GE�_���i�;�mH� ����t$͗�k�W0��_.��t����^����=�v�ޜ5�>�d�Z�ʡ��?�ԹIR �>^���C�L��ߥ��FT��)���Z�x�ɽ�ӨF
�z�@�F7�wez��%���2qsWWv^�xb㭯���੗�i��V�V�B;��>=���H��N��{抋���D4����`�&��eqm�ᗖ~�%�쿘���NF$�h��5��QW׃7Kɯ���&�D��.����v��G5n�4}#��p /O�V�RX��$�XWc�us"�����Xw�^*����|[�&�:�%97��"���,6Ao	������H�և������6���=6��$���dӺ>��]צ`��ԝ���(�4�+=Z)�ԭ�R�9�������b>��p�~�6��ИN�����TK�e㠟���A
\��рY�-�e~ȾV��.�@���c��@�g���������Q�O��.]�.AAn)�G)D�l<0������.9'���C�Di�3O���	+��[��y�U��W��rU�}�XШ��-G�AڑN����M3+a�_����٥�Ba �6SO�N�)S�vMh+�I4��w1Tg-5�K`�m� ��iЂʂG?]�;��ť����C�d�Ҟ��$%e�~4h�'}�赉x�G��ٰ}�!<��	�=��[ڊ�Y!V_���?���@r�����Ҿ����1��f�t��/=�%a�H�[W\��*d(�6���M�]]Y;E����.�׼�_�f���7�F T�H6����4!Ҕ�y�0��:^|���ŘZ����%9��p���/����Ƌ���=q�go���=���-��zԖKY�Q$�8��;o��c)mO��׿�8���/z��MyH-��Qc&Ms�[eY�}Bj�L��}�-Ak�7��ݬ����G�L�X,)aGbF�W�Ċ��$��~�p�˥�h��!�r��������j8�Z��o�N��{�J�����:l!��U.����.xl&�W6^o�1�73^�?����v��$J2D6:i�9>+l��6���><1\��Ahv�,Dgx,�rD�R�3�=Њ��g3o<���5�)v�b �wʐ[۲A�I%��c��x�ur����b�{��V�N}���|>)|�U���ů���4$x$G/t�L����L�88n�ݿ�-
tduru����<��]'�\S�&�_����M7�z��%pZ�qaZ,�:_u�8�&{����\ߒY�[ș~�Sh`U��"�&G�'��#��.ޏ�N$g���\�w�r�l��A�z��f���%[����'}4~r�%���`�_bRTl(��	w���W�$0��� i7��� B���*������^�6���d�����Q[���މ�Qf�E1{�Y]#^�rN��ޏ�g5q�D-|��?;UjՂU�iB`��UT;K��V��J�����lS�5�j���A����PFg�X�m��!���AM��f�˴7�CQ%�i�v
'�h;2�G$�)�e�ԍ�R��M�J��c�du�{3|7L%�#�gmO5��~��ZC�f�T�Ւ�c%?���d����#թ�Ϻ���_6ʤi{��ξ���J�eX�Z}ng\H:���wL��� ��p*hk��t�.=�7-�1��.ERvß)?�+�s�MH�>VS8�N�9�L��d�[�)b�lᓓ����z7�h#,���+x��(�_�V��(��
�[	��N���pT<WuU�H;]��r����,Y���A��Q׾��]hrƻ��]d�sk��A4(� ���V[/����SNec�X�Ԁƽt�'p��	�Qsn1���.;���u����M���@fg;�}�k/|�53=O���ݪ�����,yn�y��2L&��]��B���\���df5.6	������� �ࢮxZ����������FZ7Ё?���=RH���x�9�C�����a������Έ��@'*(4�N�H4�Im�V17�ڪc����a���|�ah�؟k�R�Ώ��Nݜ�z��'t��P�-Er,��g]K�&fE|;��%���P�1!�m�G�p��O�R�J;m���
B�g��3���r����u)�>�n��������n��7����|M+�8�M5P��&��F�V}������}C9�Օ�?��`&����S|�(@����Ԩ���C���7�T->uM���!���������^w�L�����ͽ��]�^x
à�����ón��>�Z
p1G��vװt�U���ζp -����ޙ�V�H\�ݗx*�A/)�9k��	K�ې.�~���A5���aѿ�ףu��2����/�u��I+9�l7���g��E��Vo��c�������p}Uދ��F�mn�۪��5@w�#�mK��s���x���{��ji����Mk��gk����{ƦU�g�j�ĎR{�&{�X���=>|��y��z���z�a���>E�<�˹H�:,�%Q�@��fG=�3�tF�=�V��p`l�æF�C#AxmV����`&bl�(�������o���x���W֕�YCt,>zy����^]:wڿ����Uc��p��hh}�욧u��s�Շ���R���-
�@�2�3~r��dL��X��y�X�$��ƺ�2��S h��LZ(�<c�w�ޥ ōLW�9�����(oN<����4\T|�z����H���z��2@� ��u`{h9ڰ+�Gۺ	�������#�~�t�P�2k��M��(��E��gQK����z@*�Q�a�	��׈k���7o��L��'��F�fe @���%���U��v��k|�C͑OC��X:��$��o��g�uHU	V�uFN�i���X%��}/�eƾzOV�O7�y�Ԥ�
���W���?�Vac����m�/�t��-��.N#	�(4@JX�;�fI��"}��tu��o��˔�4�)��q�,蜜}����T߶
����(�L����M���҉��N����1������뮏���?4��4g1R�/�&�M����GB6����y�S���b���F�?����q?�k��[s��a�N�xŃ��H�=�V�Z��R���{�7�E!��]���^��$��dH�|_t�M8Ñ����3<��H�&!����q\m��'K�O+���i��B�B�ο�t�/J�`���ΫI��rh��8���ǌ^�ZyסPL7�hQ�n����Y�%�!j���ڄ����]�_W�T��E��I�i�� =}�C)�/���yd%e%�����9FI4R^�"�w�'O��\o�|9'Mvm��ox�A2홉�:>�V��~�*���-a��^.k��~Э�X>���v5�Ec���{1�v�گ$����B<3�KS�vv&�5f�Ͳʭ��~.���X�pC���� ��݆p��_�VחTt�|�l>ף�MzY�K����F=}�멘^ ��'%N]k�=��0�6�]�{�xeo���琈�Kg�:�-���lM~��l��0tA�4�4�w������"�eԳ{�ԉX��g�a��a�Kv�آ��"荒3���aS���b~�%t܊���*���7͢�b$t�TbOA�?�9���?��F��X<��q�l���h
V��	0�n�(;�#��J@0Ny��"�>�,���-J�m]����g��puRv�g�֤���H�S�s��GB��_�6�k�.���"�����Fh�GK���5ɇ2&�אz��O9~��αgQ~�L�#\pZ�����ԃ,��8��Yl�84j,l����/���m���i�v(�Kʰ4+�*�GyhlU$���7��CCc�b���m����?q��0��X����a%Pܟd����x��Y�ѿ�z!�RA9�U ҩγ ��.�'�.���]ɱf��OW��]�-��ೱ�L&?F}�{d�������ڣ߆�y�A5�3Z��>��lK�oW���$x��"7�a�����ZΜ5����J�z��y���f�せK�_�cB��ܛ���4���#ل��,����xڪ�z�m���d��B'��f�ˏŲad���[�[mQ=�MJW�w�f�K�����ڃ����7��B��fe'��Cf��ex34&K`|���P�:�{������8u�����|�^��x��H��_{��싈%-�bT���R�i�9�)n:+P�B�/=��g�:�Z��s�}����2>.!a��� y�-����\�Y�x�/q����,WKu�D�xڷz
ֿ��(�6��r��_౑^FN�V�뜯��g��3�Ia�\M�_�q�G��&C�{ߡr��-��'����7�S5$I�v&�u��r&��Q>{b���N�1�,�b�+I9�՝F+��g��P3��3UJ��[	;
}�v�S!q/�;�f�b��l��n����t� ��P��h\��|آV.���Lf���񮈟�(dﱗj�fsb�c�K~�E�g�0q=-�%�p�<ED�0����A��sЄK�v�n�"��3xm1Qf�X'�h�;�/@G�1F�qAQ�KFȎ�N�l���K�ʃğ�B��`��E�hh}0u5���fPVpz���W�T��aQ%�&1�+�\.V�*?�K_�ǋ`1�?��Uv�ds÷���C�I� K�b�!F�W��Ĕ�x<Xq�#t$��g܆���)8f�.聂���oAx<��M����\T"��ӂ�%�%wC0����I�>s׼����fK�m4����T��'��~����|�����U<��NY�@���s�(�;��Y�`�[�H ��&�F��5����t`�3�	�CP��v��=]a�r���s��YE7?z��L7'���@��c!�p)�5���q��w��d��y����g�q�H뽘�f1���o� -_0�+*��4�31�A9;�������˕���
QӪfz^Ιf����[�R�[*��"�elZ��<��#��W�܄�����
��؛/W_�s�`�\�/У�Hw��������o�@�ɗ�����z���~o����E�þe9x<�K˩���C�΍�j�-�;6!+�{攛���t1�>����A�w�j�0�q÷a,��@�����'��NV�\J���`�˝G�Q�(�u�,:Y'	�z_q���}y���g��KC(�0�Gx�BKHO�DN:$�RR���r��o�㚸ٚ���A���z;v��dY��v���j~aE&�����/��)��\hX4j_���Y�?��r���X�w�9g�[��kʂ#)4+�����ƫ����S����Pyo���E,<C�0��#�`z�M��eE�|��L�k�Bow��V8�3�x�*t"M�i�t���{�Wm�#����F�L~,�����)�mVt��b��?�o���64\��f>D��d��*h��$�S����C*���N�o���>L�d���O�4��KSxS_-��y
���L����ބ���/Q��R��>u�b����hr}�=�_��Z�V+U}Pj��u�x�I�i�Su��/b�bk[�[�Kf����5�<e�ӵ(������e�; ���{� x��S�@�A��r��e�!|-k(��?%/���:��$�<H�����%M?��U���ܷr��;�5��j�+<�Z�@���(����[ n�E�QYO��g~"���)�>$�?�eA�	1����ة���B+��}��Ln�dlv�"�2h,��B&�S�7� 2灃I*��4��s�q�����Z�P<�Z� ���[��ܙ'(V�6<Z��ѽ����ܽ�"1~��W�TS*��s~wňo��{QE�	�	�C����%�)����!X�G���%F�[4>�4���>ׂ�a��g��G�������M��|~�Z�͠S����dV����$_��~�S����g\���%�]
�� #!��6��n�G1!�&�{����h�;�������%�|B���!�N$���t�����/h�1$��������x �(�t�h���Â"�"�����˟�9� ���\��Y7j�[Xaޡ��@'�>�n�ד^*V;84j��<t�rJMV�^����_��� ���Ȗp����*�N<�b`U�H
3�k���D-vcX�=r�w`S���8?��V�[;�$�R���;���J<��~��1W1)��Q��Mr�v��&�dT����[����w~��N�.�U�����,u[�� �6aC�J8���q�)��1��8��1���O��:�;���t�E.��=;���4	���i�ގp��
�^�ˆX�ϸ���V�oq*�?D�T��h�\�;ӛ���x�t��,N�c��t5J�a��Z�Ț��wg .+ή���@�/6�W�+W%�����	N�X��X���ւa?���^rEO�.k�,�}U�-d_Ǚ�f�9/�&M�E���� ��}�������#��Dע��AӂέOM֐��%�.]O��"n8�S25��^�ּ�7?����>��x�ЧT�9�*��F~�I;�g�b���}�ӹڧ��B�M�LQ������0���C�.�(j��P��F�C�\�*�?�y�*���d�x�V��B�5�A���{�S{�ZO^�T��t�&�=DY�꯻�L�_yx Lv
9�ի�"=� ]%�cμA�b�t�����bӽ�zU~2����W��]���kx+��\���a3��1������!9)��e�[8&DH�5Ӹ�v�T��e巠����V��_���5L��������n|>c�D��n��N����r��	�_��U��\���F!�z|�s��}��e���|�~6)a!P��O��TTL�E�������j ���H���ĉv�@��h����g��u�
Ħ(쮰���N��OGǤQ��w��~%*�H���;�n�DQ���o,���jt(-�������^N
�$�I��)K_p����H4��Aô��0"$�6M\`"�Y�J�3����ҷ�D��[���k���g'���f|h�Ώ�!�yڕ������<��xS���+�-k�]�-���o�۽F�@k�7��^���(�dM�b@<�9$,�	��F�'��2VSg����o��P�����&?̯^�g�����sb�z:��}F���;���6��m���Ub��O?��^R�����h�Wslnny���|�;5�w��S�^��.����w��M���%��!aW}��lc���)2�2p1�%��Xc�KU�M��)o;k�:z�p���^��6F�g��si9�K�9]>��Sp��,,�1�r�;��p�>dy2jv6c��19s�4�2Gu��O�"�� (�� ���N�s�驉0���Ѱ�L݉9+;�����f��i {�1�y㝝�9x�	�3�����#�^�d6R�=���M��٩�ѡ����{8W�W�[��n��0@���0a�%z��U�uro_�Qu~�����ʘ��=��Y$��x���L�uu6pIu��R���1�HlG�Q��U��ÞW�ѐ3|�Y\L���ޗ�.��X�b����r��n��B��V��D[��X�u_j!a����x�i㾅P����Z�0ٵk�����HO yxO��w#�.�mVC�?��,�a��}[�g�*�w��0��5���\����_ ��_�Ҵ̠mWh;h�_>c��S������C͌���=��\�Xu���,�v�.�*X~]�j#���`{�ʊ�0���mbղe=�-i5���gt^}�-�G>�`Cӿ����Eb2���5g��*ƌ�p:-���n�~�)${���O���0��N���C��Yk�ނ����-�b;��U��`!�y�c��M�B�����B
b�����k0��Ҧo�|y]�P�eUm�l��d���bt�ë���B��k���[E5��e!�! jV��)�)@-���ǚ�<&r�����W�*��.|�������fFu_?��'G����}��<����Gi�����ȑ9S.c2a��N'U�G�#܉BX ��ݎ��5���f�vL���D�=������^�M��D��/ts���vv8L��P8.t�jwn��~���R�ȅS�&��Ic&��	{�R@�h:URG��f�Y�/�rt{v���<'.�����Ռ�{׆fZj�ߗ����(|th���'&G);N�br^�迃�Ȧ�qiV��\�j� m��᪩s4�u�7����Q�p��7�[�8���5�K3��#�l{���R9�Jǜ��3�������禢��	;���:�Ohc��'��Bh�BfcuQ�ő#�Ρ�5�����F_����Nz��1ve�;�H��Ԍ�a����HGI�24�$}A��7A3�M������psm�+���ߩ�Y��t�W�٬���{b�2'ɯ��j�bq�ї㘔e3�����~�n4.hxv�b��D{� ��_a�*���I
���ȸ�	 ʘ�J�6WP�{t��%%�J��o�7{>�'�0a�z��&��t�3�ik$*�:90X�\d�q��7)���:l�Q��0� n�,
c!�[��Aa�Ň��.�F�Α&5�S1�cW���O�c�ݎ_><�{vK��� ��k᪻�~���A��f(αV�7��N�1���N����؃���-X
	GS��~�w� �~�mP���ɑ��̍�j�n@>�5'亾�0�o�AfW�<��Мf��!�xߏ�;�PJ꾟F�dd��၏���I�-��j�O��v��(�=D3�"�%O��CUչ��CV�(���p�W�����%�}��P&�M�'�A�-��2?���W�gY��ՙ�)494��e��^��$Օ"�Z�V������h�w��|�2|���T	����,�]R�WE�S�N@�l��~��Q�#%x�ԧ���f��[��t�d��'=T�N���/�z�Z.z��H�uI��J��#g�
��z���{}�sC�f��E��_��mg������j*͆����TNE���"��pe�Wvz�kj�&�p��js���/7�	��xf�԰u8h�掴�C��|J<��]�nw#:&�̓�f���9����}�X�9�ߜ6����������r����mt��"L�䳊�[V@�Ƒwٱ�d��:�{sS.3���%����Q�p7��;X�?R:b �H�\=I#��;�i5z��h����}yXY�:��E��]��@z4���O�Ԭ��K����+��9�/�X�9�l�����e�Ʉ��U�A��g.�3p�ZЊK����E}۽O@���B6��GS�J;��J�e��^`ZOG��^ �a�P`s�w�Ǧ?������S�m����X�Ԝ֘}���,a�o�e�F�ny�!۟���n�Hl�K7�-�΀���t�5V{:� UZr���L����0�u�Z[�2c"��9a�(�ƥ穢^�p���@);�Ge�`�e��2�g�����7(E��Z��k�8OdhwL}�CΑj.�e�h)EXRHFL\Fe�*�m�lA���zCl�.l�/ĸx�H߻�'����R/z/=��Qﱳ,���31u��v��	�6��=$��cs���%ʁ	/�q������t@�>�k��`���F>�΃9���o�]QSBoŮA� `�E���LP��(��>����i�ַ�������MF�f��nj�y�o�s�G�FI{ꛞ���F���_6q�'���L���N�{�h���7�/�[����m�\1�5?#���Z�,rޛ"$��-ސ��_�-^햁�V�-��[���`I���(\C���8oL��D�}�5���ߨ�a��	+o�Q�=�`��Igj�/��1��	ƌ�$~T���7�l�(��23�J��_�+�p?c�[�>=���&{[2B�Z3~���rބ��1�\畹L�UtW�=����^�&�U���@Z��GK`����E%hQߗC�G�Lኹ,���Zm�7$�7��ՒK��u�H��z�?�_
��-�%(������UJ�
����y�xߚ���W�dN�/��C-��J�զ�!2�$�wBe9gRe�s2XU�%� �Jg3��MOzm�)A��J���C�	�`Ԝ�4�E��96g�o��K^���9�94�������v��<~~1�}ǣ�s�����k.��:<�vxut~�[oy�,���a�5�w��X�N��/����G�Y�pa	ώN�A��l,��2.���C��'$x�%G���S�zn�5�
�	�YI�:,�����mv��"Zl�g�V�(v��s6��n�����o�E�uѻ��k,N��L�l(ƽM��.�xI��~�MtzvE��*�Y�7{�w�Kc�r�
���7�	֜M	(����q1[I�qu��ߛ�$�pU��@s�B(�\��#������V�oB���m�,���yvK�<�b*��^��{-mA���V䀾bβ�5��f�W�<�8j�������1	�e��s�4=��&l���w�pt8P�!�7��r��s`n�^ sI�d�x�B�)��:4i��/��|�����S�� ->_����?�����J#��u�x���tJ2l	�Is�Kb:�IU��hܱ�c�+أ 
���&������ cW��zm�
cnz�+Y�Km�=Ң���4����(g[\�:),T�3M�b@V���l�y��O����>~`o~�;Vek,s�I�'tk�C�v��9��q��DFSy�y觵zxG!�������|��N	v+>�Y�j�������`K��O�ZQ>�à9�Ӫg9@��^�,q����$�'�]�A�� ��ئ<ǨE�ש�u%�;B_�u��p�׸;&�+šA4�4�3G]�H�>9(P'�ف �e(?HP��^K��^P��0-�����F&�֔��k�,�(о�=��Ky���s}oA����.}dO��+�[�*s�ޟѐ:�3���Zs�V��ռ����%���k<R��+�Hwsso �p�����Oǉ����H���۞y"�P�XA��Q�	�������o�(�V�����Ѷ��߱���O����~E��b�s[�2�;�~'���Xc���N�� ��ȴ�qc�i��|�7����g�x>��;�_��x�Ϥ�w�69�ᴐ�6��>�vz�눾�`�˫"O$�����D!��ʹO��}�d���\f˥�1�C �bJGag]G��isy��ʬDY�_��w��J�������*���|$]��N�oN}�M1.��O� ���7㹭���s��Lf�l2�b�-i�FC>��ʘU�/��Ɩ��1�U JO*H�B�B����u���E���q�4DZ��I\T4Uy���([��?�1�NL$�x����k}����gCK��5�]�ݞ���f�I�l�p�Xz'��tS򡸖,_��g�l�i !�ߏ���8}�ub#�\�oo��0����Љ��rҊTk�S�b���b_`'���-�|juZ���_���ږ�"梛����a��to!u�mV����5�/�q��t�7�.+D/4/�z}i�S_$̘.ʙ�j|�?��7�s6Q�Sb�ϬgM]�u�=��V�\l����p�H�ة!�/��ߧY�˘*����p�)���zĉ�t���Ǭ`����V��r4�$�=V�9bx'8�&����/�/��<l�U�"�Qw}��5� C����t(!��`�߆oo�0��%�}J������3��x5,:Vnw�+�T���y{ϼ׈+��?�()}�Dw8�KT�?�~E.���^�wk���a�c<�pH#k����.�4�*W��Z:��4a�Kі��B�jyY���c�([]�6�h%$�o3!h��6����WR�<��U���/�XX^��^�oZs<���[Y=���E�)����B���?���kWK.d8���"�0^���O/��ɺ`bJ��*����,V������B:�D�G��a�o-��G.��{ǯ�k�M�[�H�i5X�@�	�f}�A>	�_!����\��/Y�׏-1%�G��u�pߛ`�ZO���޻�B�NVb��X�8!��|���Z~<����h��@u⬄���;��C_��d�w�����'֪�j�;��-�a+r3D����1��A�oO{�ԛˠ�9��X� TwV�`6�O'�>����M�) =7Ξ;��@:������g��x1q����鮼��ې��3о��3A{���x���T��|���
�xl�jx
|g��3E�|΃�J�=�;�Hv@��Yg����!Q�k�������چ}�i���bi�˴�ŵ�`ۼ��s|_�}��Og^1��S��W�۠���Ң����-�_)�k���7c����6VTV�9؈���d�iN+^���X�̝"��g��A:J���	����0�pWt�7|~�~9~~�q#.�������|����t����S��N`%�g%��m1A���n�(�?/��nA��>ܤ�GO�nrC���e��F�7k�`z?����dz�9�/��d��E+���\��1�Ġa�Zs��Syw�PY�H� ��ҩ��ޯ���0Ǫ���]�m�%󃩸��Z>>�\���p^S�'Y�
JlA-�RO�&���p�|:��2>����c�	c(�1JN�LL�*_�}�q�Bh�)�f�i����ڷ4�9� Q��L#93�@xRʻ<��o0�f�ڪ?�S�Xtc{�b��7�A��H�^+h�'�}m  .�b�ꓝ�z�ܿ;=�����k����P�CX�4�V��`8���]\���]��Ir��g%-��-�7t+�*� a�
�Ꟊ[@mՌ��bllt�UOf[u7r0p.�N񍟅��G2)3u�pS6k�T���5&&��XIUH��E>���y�����9��}�Vة�w��L6o��GQ:�ξ��A��	�&Fx��Z��Z�����=;�����W�+�
{gc�ϔ�sEC>%��o&u�,P�W1�N]�Q�j⽇�@�椓_�A=�5C3G>*��R.����dy��3�y[�sm�[Rs\폥rZ�3m�O�w)�C2���f�/���(l�"�@��Q)�dyI��������cDs�*���7Ă�[4-f�5å�%���Ju{��ס��Q����	#�w�?.!]Ne�4���Ԫ�˅��$��%�!ܝ!���o#��&��\��� �g�c:S�y��n3�-W�ה�����*�-�܉�3��U�����h�i�8��$Z�ǋrl3�[4*�s���6.y���	<�c����C���7��S���a�L>�N�9�K3O�� Q�:�&��{�T�w��v���v��[ �n B�Q��^�|{��ؓ���׏�{#todm�1�����6���[�u�n3wOA��ɀ�H��O,�\NۗC�`�Ef*&��?��ŵ��j8ژ�P��Y���+\�#RKԠpOD.r���FM��ctdGS�����+k_�Q݈�oG ��8�1�����b`I�0lL�b����ߓ�R\�ui���F���H��E:��a,b�~h�z�%$_�L�b�Ǌ�4ᢉ ϔ>�A��߿?�j�̼�t��3K�� )
��?7��nW;ܟ#}�%W�\2� R��E�1Y�ڢ�2	��..��G�F��q�Y�2��r���e�����j{a�a�Y�zŤ͠�������_u;�]���J&z�K�O�Y�AÅzuP���8��ͦ$l��at��efl�آJ�R�Җ\}���;����������JT^M:z���HVw��ÀjCD��.W���	�d����Y�|�s����|��-ead�Üy�	��e��6���=��S^ݙ����n���?-�	,\ߝ�L�k�Y/�s:��b�FcD��s@��B�ɑ�yɑJ��Z��e�&��>��u���Y~�7Q��Iļ��.S�<��_�վ`��}��E��zI1��3)��3:ߐ�	��t�f���z���jxiZ�W6w>�	�;�B�/�Z%z�0�E���V���ZoB��	�9��GG�E=���
twj'�����2�ˇ]B�bbi�	2?i�ƪ��@尀!�o:�V��qs �8M��r��Z�n���_Pap�Ǔ��	T�.4��4����w<=z��D��%���$l��º�I�����{�L<.0w*��0��`��&�i�Vf�j��_��8L0r98��X9�=܎̈́;�����S�E�~5��\˴��%E� �e�
 ~$_����[^�����>�o�k��
7�W5(���/d������Q9�pQ���{Y�H�HaVO�dN�H#h��xY�?a�I�^�^�����ΫE�	~F3�������$(�w�a��������f������Ĉ�c��������\�Z��.b^��-�׻eIǍ��_ �{p��gx�S�1�d��HDGO�pk��#��"�y�"�V�����B\<C�4������$��0Fmrl�.E�R��e�pgeaY��+m��]�W��[�h�
w~<�6�8~(��;��������>}V^��T����)�(g�����YA������}�g)���QW�~���h�4E��׀�%F7�Ow�t�)�aʽ!���a~����I�m�Mװ�l��y6�4S�L��Ί��l�6���/�
6�[С~��@:��Q�uY3ύ?�<ˁ�:��:�p&eN�)~�F��%���'�g4Gw{��.&�b��*ź�@��{_H��4?��Td�@O���gT�玐l>��
��m�E�@nm���1�p����f��\�e��]l��z��yr�K
تE�ʳP�<YK��M���P�\cc#-,)������ݝ�~9m{�&j~����B_O�d��ku��!:1b���Ѭ�/4R��w!�r�׼B��Z��-O�ZM81����1�_ζu+F0ם��;����[3ֶ,�O�f��vn��YV]3g��;ϒ��/6��e=��/n�k�����ƪ�@X�%]��!t�]��xEm�mX,�,l��܊p��G��þL�4��g�k8 �_����E
;N����]��= h��&���Ղ�{2%A��)2G�b��C��o	�������ɇnC��چ
)����w=u@Z=��Y��b�4mA�4�3i���i$��Uz���%�q���	��1��&�w�H��O&GNa�D�v�g+ōZ��h/�u�O��옓���H�W�О�Df�$b���z4´%w�0�/d��D�����z��k!1ᮟ$�N���m+藟���ؖ:���:	�+W�ԣ���1�k�?̌�k��X��P0��� jޏ���#
%h%6������������#5{���Z6ه�Re��76�7lQ�@]��j�$�r����}�f
����7O�%���뒪�,c6��V�t�����6w�7�zOE����AC�pT�s����=��%�� �7�-A˾)�9F1~�rTDd��ߧ�?��[�C'��r��L�d�#��[
�Δ̘r|�AŨo+�[����q�];CSv�.�w��@��o�I����J�Jf� �)�"}V�񫙚�t��!"�=��p޻R���39w*����o�:�lJN!J�X=�z]��:?"͐�N��O��T���3r_)�����1��{+Y����*�P�2d>����6l� ޞ<�qRE��[(��)����@�P $��<��&2@�
*\ޒ���X-��g��*׶� ĩ�UN����~㥬<��t�%ʥ׿17�K}���颂���M96������p*ܹ���F/���,���	Ck���*U��]@��!�L����A£�����k�HO&u�9T?��x�&��M�ƃ�FQq�0J$
5�Ճ�;r�zt0M���`s�@��ia��iX]ѣ�߱��g���� j��U���Y4|�`1�e�J�M!o4���E�J�_|�d 摔�H(���v�k�\��2?�x�Bi�^�9h�w=��Ǵ�nF�'͎rBD�S��s��)�8�9�C���RI���RW{�1EC����և8O�ddnԧ���;�S�SE��| i�}Y�;v��|�Vޘ���B��Yv2{�m�U_ĭ·V�C�]�=v��z�Kϟp��Z�Ӟ֨'�4����n¼���fϿ���1�aa�p�9�w�(��l�b�vdR��LMe�ԅ�v-6�/7����x�޳�[���4!���T7�� K��V	��|������M�݌��s�nJ�>̟��O-cR�ժ�*�a�ݩk��C�Ɲ��)82-�i p����ӭ����ؕ|�b��!�u�q��le����H��7��,��ф���
�E�H�DF�j_R1�5�B֭�[&mI�~��V�y}�� y���vUR�y��Yq�G��pz_c3���YIs�pG�P �%8�>w�����tn뢥�_�6�����/R�9��Vpp[h��-%�[?ƺ�=�Tg�RKy^g'_�jԾ�	[�2��F���ަ�&C�j#��(���;ʬXޤ�?.�����}|��	��)ΙNG�b�����%~��Z�Ѽ-����5��2O���[S=�Ԁڷo߹%���K5�(i�g�d�3@��Ш�Q��9�b��~�?��rD�a���K��D7o��r�=�����S_�w>ݰV�^-� q.<i���5�V��Y�cr�j�?����UN2,� Jѽ0r�2�_�5��F�`��T��,� 3sg�kp���Xꚓ[��j��'rBۡ/&���m��$n�R��3�X�kt�����z&�Q$e����_�^>q�L�7��G\���	�/6}.�����wԧ��Z��T�i���L���qD�y{z=	�"z��WL#�^�/�0��0,�D8�%���Q(�6ؾ��"�6LX����~1���*�)��_�|Q�q�l���`Mq�g��d*L��0��;Fv�g�
���g:�O:�v\� ��}��}�<t��l�4\�g%�M���nG��ڤ�_ퟟτ�3�x��<z�$�i��B�p�w���p1��)�8�8|Vᢳ2"yZ�w���IZ�����9���M͟��..A��6�Q�xD��F��2�v<ƽ��tIِ�݉������k���CR�4�%��[/� �K[6�W) ҝ����W*�׾�pq����G�Ng�B���8t(��^��.�6�����v��"������o�TX���rԲKMݕ�
�+����P�p,Մ��I�����&\� ���^��M.^���a�4D��
������r�߀ji�?S�u~]B]� /�v?Lx!���;����/�?�f��t$���Z��_�[�O���Ц^�Њծ�)��ۏ7�����c�½���Z�WCP����{�v�[=:)SW���ڴ�5PMq6�S���Ɇ�	\]�t�x����¬ ��dA���ۢ�cM��^�-��OY���|�����ITԎ�,|�Hѣ����������3=���em��M���\���qc,��:�= Q��-S�x5k���#I�v2�|Yj�@>F8��~%_��P�zJR=ކ�^[��v�����~X��	��0�¸�8�0=o��+6��:)�:�[K7���9c"���3f��
��H��ם`S;�������g\�p��ȓF&����)�`>M̱Z��q���u�f�P��t�TC[d�%����!��c]eq�Ƙ�����-B��,2Ћ	0l�b��W�sēh����TN�n����2�qj��g���C�6�h�3�H79���"��d�!z�9���5�v�twh��f��O�5~��n+�",F�_ۉ
�
��Dv_O�e����^;=��m�s�.���K`��3Cf�ͣ�Mu1;]�S?�D?���N����	yr�����!.����qR���%e�Ф�>p7���l4�&��l��Q��$�/��%�%����^��_ �|��������a�{���5W(�Uh|�El_��vV��x�DN��	ze2I����݄�1���6�B�CL��l���9w;�l�+��iȀ$1�s�Vw�ɫ,�����k�?;D�\��7�w*�9�?���C����6��8�X�V�i�qa��$���7��Y�������E���z&z�[흿�C �=�(j��q$<�<�Q�mX�����A˴"�7�q�����>����W^�+�9��M ʜ�B�o������~8����b�F��(�OF���	j��Q�=���ֆ���!Dͣ�kZg�����0�h�]���f`|�������uř�����#ۭ�]�[L7U0��~$�8�,T��ze����D�'C�F���E�udH��CG�6��k4V�7��w�dZ���NZU];�&�j�f]T��y�������'s?�0W�UF-���g%��`*:T�eY�Ӧ���؃��۳�ŉfm�4hy�����;�G��7���(���	���'��ŷ����n\����
s����I�7�7X{�\n�<fp�/�J6�s<�����YU�_�1�������v	�bo��	D�C�R�+�S�(P,�Ǭ��?H�qBk��Wk&&��Gi����"�5|����J�T3�]�k>���DQ��4�Gv��IK0�&-)s��|�!�T�wxxAݘh-�9>�;n��/y��;[�6a�vMg����������^�c���P�pt��e�~���d�{�gAx�c�^�������Z�{���rO�6��r�h��Kˍ�L#�3�{�#Յ���,��:��iP��"#�p�Ʌ�_z� @�e���0��BC�]����'J��h���'8�D ?&6�j�+g�Sw��e��*~�27��r9	��M�τ@ڞ�	UHd~Q�d�L�Q
���詋m~�?#.vZ���^�s�3�2�e�{�d�:Ǌ�n�5: �堼��YEu�� Jl��
���iI����ռ܇8�n�>�5�y���Nf�n�B���k�/f����S������o��RTծ�-����ڊګv�Q3H[j��+(j��"�T��ֈ��#� ~����~��s��u^��<�3ށ8{/,��N�ǦN�>#�/ҥ,���I�
��kZ�6�8�9s�������K0̾��?�rM����	���p�fڰm9R����O�Q��������l�����	�&�v���`H�q�D"�_�2�R*�xL��+�P��|p@1 ����+�r���&W���7Fc�#T�l��u���sC�G�pB[m���x�R���er|Ϩ�j�z�������U�Ţ!��2P_c�G��j�߂�������Yy��9�Z�q_[��/!Z'�#i4��c5V���m�'�%�;�9:�8��G5:s����� $���}szzJ���b?�ڊ���5s�(��[(�4P{탢�P��G�~H������%���d_������pd��j�ܼ�(g�T�G1��x[�-�@��a����'��,�@ʖ�����E�.����0��j$u��KD�&(�$��Md��7���{���שS0Ur��ɿ� �7�!�eD�C[���O7ëø9��F�l��т��u��.n��˞V�"�[5uNq8�f^Ď��������*X^d�ŭ؞RX�e`Z�I �;)q��r2��{{P�ZK�z^&ZjL�nB����L��ς�lF�I9�9j���L���%[/�B��@���Q����t23�(�s�r�
w���dj��?'>I	�?���G!�1u6[�9���9��GJ����J����#e��s��VN�͋���-�3�Ҝ	�z��u�0c�� �C�;�a��Y��<��g��m�������ԗ6x�!�rL���~��^>�0�׏��M.������������g$3Y2ol4�cl#h�	�L��g�iR��S���yV�?]��qi��G�0�<�T��tN�UnQ�> �鐈��B<w��^��p�l�ֶF��^���B
�6�3��֒'C	����!�\.��w��
�'[�ue�H���\�5�����2$3,�=徊5��퟈6?�V����<M�7[	���khߊx�e;L���@�x�Ī�X�L�C�ao_�N7��y��%?;����Yi��غ�� ��Iʽ�D��������y\�M�.,.H��Eu��{k(C��`��R����t��P��H��}S$kj�ţ$��w�R�'�%�V�L���t���L��w��W�c�l9�w��g�^����<���? �+��󴥢"QyIH_J��vi=�:W��묱9�TUۂ��Yl�kߛ��N�lh �u�1&�M��)J����k�騿-�ky���&����.�R�g長4��b
����A�����G�	��r2�e�ѫjq&-����A~�3HLd�#Ԁ��g��/2��w(9�.S��a�?��ۼ�3}N�15�6iS|���������p���cM=��Vc�|NB+��(C��ۂ�~���[�jp���`Ͷ3S=
)�mVÈQ�}FZV���qO��k�/��By���S�2-u%>�9d�˹SY��v	g�ǰ�$��ϸӕf=�ĉ<�i��j9���,��Y#N��{�˪
�>"����P�l�l�K����>���)���h�.Q֔/��� &�ޤ�Ԏ~c���c�j=f���� Le�/�!���n���O�6^�S�zs���Ag������s7��A;�7��
�	��R�L���e��.t���d��,'�)qM�X��ˡ��3�O�3u�����Y�/�?t/'q�!E�[ Ŵz�L|)��&�2�_y�P�e�Q��v_��A~�nҮ�%�ӏN��� �/gY?�ڟ��u(�q}ti��񦲲pI�r�NQ,*�HrM�~%a����ND$5��C���a�i��ryԱ�v^ix�i%��a �E����)<.�Վ2�B��HJ��h�d�Ϝa~0���X��9/�����[��%l�Rµ(�4�{L���_}����K�"��Jq%�;�S6���F������$V��	��a��*v�ǁnh�/�;ы�K�eP��Z�[���)���(_s����l?�2�gA��6�=�bC�M�4=�w%��(qK>B�%����\!�}<6�B~��8�r$�*��oE���[*����ݐQ?lH*�D6�J�)��o�ͭ��}#j�G��yXG�赹�g&{ Ɨ���������Y3���^�8������3�η~J��[�fz���+�I��W��Ȯ���q����ǁ�V���'#K��}1�h�ަ�/������ƞ�_�I�{�Y�k��ƚ��jWk��bʆ�W sa�]j�]�6�Hzs 	�'�0����+w]���8[��.���Ɲ̤�g��O���}�6r�X>�K�`�wt������mC�'L;N��GGG71%OR�a�ON�b�^�fd�ss�5���!�HQ�EZ6l�j{�[�f�� ���3`^n�Od|&�%�*x��O*S�*��z��h<Z,Z��33B�Io<�#����]�M��T��clw~�#�X�#T.)Gjؾ���m;ku���U��^O��fM;�*��$�CC<��<<�ʃ(��}� ����\��'�����'+Ҿ%���)�t&�E�� �X`�ђʁ�:�ӑ��Gc66���oG	Z� �%��D$����c�=��0�Ȑ J��F`ل#��d*V�F�OJ�L�o
�f��7έQ�L���� Yf��z����s���l��!�o��KIO�I�F�;Tg���	�,��\M}je���hL����RVG�\�J��b���w������͑�=v����)��>�	R��!��~$�2�F��|3��������+�3����nr�R���U|�<ut^�Ƶhtʯ�0֨�^M�|@��
���p�6kyb��{�u�0�Iɷ�V~�#O�Y���[">�1BU�7�O�ps����J�������t��wN7��q�����q�3ʨ�LN�{�jѮ�_}����߸���EL�v�:��1ڒ�Ǐ��Ӗ;T�l\t�zM�\th�OK�J�<U�{�,7 g@G���!���"]@����{��ė�7B���!9�?#�vys��k�n�a?�.�ߑ�Xr-�p���0ͿC��|����C��iaj�����
�c��uH������l��"�J g��ꉀ�O
���Wnl�e����I���T��m�ļ�-2�'{�7}��<��������;��{I\����1�܁��;M]޼����A�9�����/�?T0Z�򛟎d8^{�ykǌ��p��E0�wģ�ސ��v�M���!Z�
l9��v���p�����E�]��K+9P(	���-�p°Ȣ6����o�=]�]�����k�����]�}5e�G��TRy��0L��$ii��a��f��Vq�v�)����=7jn����oG7 Ȁ\�з�\��i[�d}��O�	ݱp��+#�Κ��Ȱ}�.�y�m�g 0�*6�r^T~����N��dB��lH��|���鏗��,g�c�Uϫ��K-��i7Rㅭ�}��t9+��tsS�~���<7]�:���I W���N� �a~�	�[��5��R�(�6r�΃�1Eh�gd5ݹ�|"�Y������*�3¢�{�kC�.0����3L��scof~��^j���d7'�����)��s���b��QDM��<����q����&$��8��75�P(�݅sTƿhr�^�Ҧ��������%����d䓱�Y�����b�w$}K��"�`��>0����g�X\���lW�0bC.��C'�h�Z������xs�4�ө|��w �R�b5��h�=Pώ��ȴ%P�W?/Qj���[1�4`�ـ���D�~WR-�7��W�x������D.g��Ŷ�R�{I-�ɦJ�L�)�/�,=[x[��`�Rz�e�?�y��X�;�NӬ��a2����4���y�[y�.��Nț�:~��lW �%WV7�-+���<��DD�edZ����GA����}8��Ee4qyy��E�:azx���p�똹=�=�!4��ɴ�#��Tl>-q��y�h��m�Zն\	�!�L�^T�]i�}�x^��2�3M���#j�����Tq��I�m:�@7t���H�U��m=�'�"S�WSx�D(�<!����8�W��̧[S��1$h�ц�8�H<�nGpi��x{�S�ձ���`׃���TGH��?���^����S
�1�.$�;PP�0�LY��/_����L�XD ��&[�-�۵����a���[v�J�.��?�ĹlBʑ��y�r���KAO�s�[}{ȮO�2]� L4�>����� �6�����_�양��d���lJ�G�m������=���.I��0� ��K�w��^�`��--�,��GD,�*�6�4���k�T/��
!nT���r@ϡ�D��(%�eJ�N�40�2���B��*7��C�#_	o��П�m�5㚨�R*�WG�>�T��a� q5���AT9�w��AM�v��@@Scb��p�}ǾV|b�a!i��zw��:�97�����Y�%�g�,��6���g_�������m>c؍�����gg�S䏕�%�3�=lV�<~��ՠ������ܢ�}�,y��t�W�L�WG]ӭ�j<�g���2밻u�6�4?^z�zZ��`T���e=Y�\��n�%��F�v���7� �^��Y�K�M�|���f��t�v����`�Տ�a��R@�bKΗ�%�?�:=�}�V��+;�&B����L�w> �h��#�������%(
�;z1	{��K�k��������}Ͻh\feb�{"�]�t���W�U!h	7��;C��U���7&��R�!Yá'�^bz+<�#P��y��C-�"l�����=�a�<��<����~�H��Ձ�.��tSR��PN��[�}m+��g�ʍrN�z�z"�z�9��ۇ0�a#���f��/���p(m���d�ꭁ����N��}��t?UH�:t�ZXQ\;�np�3�;� O�;O��K9,�W+�	VFq��C�>���'mѧ��8����f�66�޻U����s����2��:=u1}:�	U�S������}#�Ҋ���i�c�8s�8��ɦ�.e؊��ۄ��B�L�`s8N��;���u�\��G�4�p�����UO<�y��ஶ��&�(�ɩ_p(�����x��_�O}枌Ԣ�N*�ͭ@��� bܨ��.�\�	;}�rBoX1G#h�q3��F�^���h�V�������5��s�vǕ��Gmʁ:��Ԩ��Oo:��]��Q?���w�k$3G[{{1�N2O���vTu����8�q��)���Cu?<hA�n�,�o�"���=���
�]�z�f��5��z�.�=����Z��Z;���oW
���t��a�&�D��*J�ɟ�
#K��$�H���&��Y��.�P�O
Ul�b�KZ\C����g���U��̿���J�Z
ͮ�H&�H�%�D�*�c�*�������^[��U���B�%n��p$BB�6.+�:!��01?|kι}��R��J�s����&'���8j.JBF2�6rY���<�}�Q5�gf2o�5ڥ��Sl֔�ץX��r"~���P�PPH�b�*#L�90�����pu�����������ԓJ�QX`�ɏ9��L��,X3��f>�0��W�F�å�ϓ��1Vב�k�u�[>�8K+�)����!mo[�r�o�%c��?�E��!������4��)0�#-��$0&E4���]�=�:�����m�����>V�K��;��� ��+_��\]��U
[f���aʁ%��.�Ưz�ή�����/n!���X����w��Q؃�E�6оO�}e�E+�l N�Z�0+Mߛ2`�u
"Ŧ��@��Ol2^�|���x��bі��v�N�����$MrC4z@���Z(-f�ǀ~ykO?A\��)7Yc��Q=�<�6�4�kޙ5{�ٟ�x�t���|��~��`������[�P҄0�"��VӢ���Ô��,eB�NmS�^8+|�G����k�!�}�M;�K�����z���_lo�,�h7n�F��jİ�1z3�/�sv<�#�Z˾�iV""�c�vk�<㥰CY܌V˪�n`.M�Y�/0<\����hV�v��oV��_��m*?Hzm�E2���M���:r9�12>ax�_��>�Qi�XR�=�QV�Z�7����11�ϻ��#���9�l���}]����j�|k���7U~��c�X�r��1���_;��^q�z�T�
_5`�E8K�P]�C����	u�t"@�Ͼ̴(���T�څ�9y�h���X5>���52�ye�:|�B���Q�����{��,q��k@��X���`�Y.w-�G���7�_08@#�\F��:���P�n0������U2��b3u#���Av|<��G�@-!wz����))�1�8�2	���r �fr�|��~���O��M��"<��׎Ez�Ľ�������zUx�����W����igW^Z9��J��N�dz�_�u1pkp_W��c/��%%�W��6��9} Q��L�V�)�OQ>K,�B�Y?��gf;�Y��O?Y��uי��"&`Y�~.���g����)��>o�S��s:���B՘��MdH�js�d��mX3B_yp��២մ��$rO�c�f�Wu-^r�z������|�����U�^���I��|�Ѿ���ldh_��q4v���Q֫5�H�pK���C*�s���w�1vg��r!�'�֫�a�:)�T�	iJ���r�9��؝�3�01Tm
p�{`���ddde��q��bWV"�C�=@
+�* �u0�xj
S�7�X��8|��j��q��	#�.�߰>.�t���]?<����`���JYk�iف����>8�VM.�xv�"gp��L�ع�@_��@��U�w&ȁS�د����Ͽ͹��+�D�P�}�7�5�����/�0�A���;U�e~�7��˼�\S�4��� =���jO9'�e�\����m8�4=�^���QS�̱����v�+UZO�p�U���/5`��~���1uL�P�j�R���Q�OQ�96}��9����������,_��X�[ئ���8xir���&��ƃC2~�s���t 7o�T�������Ħ��9T�se�yZc�F��u��.��r�yEC�X<�����;��!,9"\x��U��H[��B4?�/.^}+u��������Ƈ��'n���DK\mŪ�-j�`���{9������, �j��4B�a��g&36��p�j�'��y�}��[�m�>������0�����YoJfa.-�RW|���~��|s��^��?�����f��G���(�]>>�	IX^.�TSAO��ڜ^/�B�Ib��)�y �U�?�J�A���^�O�] �p�?e6쓓�Y���$?~.:1�I�Q��xA�������������{�W#����ȓ�1����-��Y�avG�9@������P׶;!vq=�&	߷N��Vu�}��~���d�n���p�w&�{+�A�[ ���dV�U����K��v^����C	���AǍb߄�}�,-Y?R\�Kڄ���:�Er��1OE��O����,7q�:y� a<��?:O>�+Z������6�{�h�|d���-���|�W|$%���GۭT{�w.�@mU�2����=�����������W���� }����J�u�hq���<�W�]3}Hjq#���5�K��>�S�?�+�o�D��� ����o��Ŷa���1�����S-��L����.j����ATa��j� ~�Vd�,SP~��0��&�I�O��i#�I��4��,q�;Ń��P��k������>�����
�Z�'����M�����n~�d��k��#������s������Z�=x�d�S��ܞ؎���m�nw���(���҉��zɁ}�'�;�,�"ubx���Gkl�6�UϨ�j͢�W�ӥ����ac��7���G{.��r�1�s��CC?�ճL���g1�'�5~Y���ldvLgjB^�L2��E��^�i~��,_�w�"���SjC�������K�p*٪%]=]'ׅ�U�����<� =e���8�"{���J�n*V��Uu��-A_g��3���e_,�}r~�����Jߨ�S-]����U,�B��'�ZjQ����+#+y g�/	 ,6)3ݯ��Y@�Q��ym�ݸ�B!����Jݦ���ô6
{)�ЗpYUn&�p�T��
�0m[p;���)|x�wD�os!����wS���+����[��V����316	�!�~�,�픝�?-V�nE�\|J_�[} @)�!���;���ՅP�咑B��P�u�H�<�����{*�v-�� �oUݴ� *Q��L�X���jI��g�����UjuR�M��iz5��$
R������T��Y�M� �,�.^��m����[��S�1�R"�0q1�#��j@*��MȨ����J�Y�J7�yO��ï5g�]ea��%�kkc{]�`��J�A���<Y �؇8n�*܃a�Q.�߽���\3Kͼ�����㡥۪`{~��b��;���/iA<�)���b	�1@2�5���x)���3�T���_g#'9M7�[j�Qv�����hM4�[�V��k��Wy�K� k����zA-��>�2'�w���������^�q�n��s9�O�+�i��5�(������*����氌���J�DJ��0�4ɚ���Y��(�O�Qϓ)��/�{q��p�Z-h��J3�p��Yiӛ����
n]mn�2����M��K�������X�efC
B��`q��U����VG�O��М�רO)F�)����T�@��N���؎.��\�X
��9�����{a���n�;��-�+�G	�:�r9s����V,��M�~��rK1s�i��܄��XSI��gѴw���/8��ͻ=!!���N�n�v�H��Q�Q���M��&�i,n����I¤+%h��n�����ٷ�0��W_jW�}�4��b�\d�rHz�1wMcKv�1i�\�� I�'�I��<i�Hy�Gٿ���HO�z��0����������S��҃�n ����6���+JE��#�� o?����0������ӻ�4�ݫ����d��{��_������"�f�L{��6b��1<�0b�����o�{Ի^��s6qp՞7RI[�X�Y����KA�u���ﾄ%4��L���O��m��mYu�lt��0�MY�����w������.l�t �E��.wҖ!�����{ZӰ�v�0i1�-��f��[���7[�	����$y�b֍��뢞g��E����n�����O���u2"Y>�y`��1�IGkR��GZm�� �e�o�d�T�F�����.��G��%��!���*>�B~8{bͽbR���$��5;���*|�AF���b��)���]L��,[��.)*��o{�D�k��{n���?���T'q��\��נM�d삱^��0L4��{�j��̓�˘fc���o��v��wq���KמΜܝ�ʚ�� �ڔ�?������2���4rD�������n�����^�ģ��$q��8kt{t�}-�j�W��u_Toٟ��y�@��z�1�tL����xz+{O^N*y���$�h�H��৫�@��/�;L-KH`a�a��5�P�d���׫f��Y'�������8�r��R[�K�n/���oh��L6�'($�p�/Y���#/zR2sb, +�B7�I��_�1���yh�(P%�b���+�G�����#����n/ERt�F�qe�di
. ��Zd�N�l���tNv��qq�/�?�k?�]_���E�w�[����?C�sJ���V�[wc���гJ��x���&ǯ��pK�����;�\׷��x�Ϟ��`�u�䴝IVj�Μ�1K~s8�\��̦K�(�%�5� � 9;7GV�x'Q&�m��Y.[c�ix��"�k����vr��::ȉ:_��	.�������5���qc_��YZ��&Y�w3�I��z��r���<��珣<_L�g��bH�/KU,���԰��6����SRn7i_ŦrM$[���x�r3}���&��l����,�ۜr��"���2�d���ҍ&};v�:�"��m>�qN|�k�*�3�|蓟�X����(.>v��$��O!䫔��OCDg�Cʹ���Ho�E$|^!d3��H4������ٻ �ddi>e�	�Ʈ�4?�EΔ�ǮL��0�w��/����q�ݼl�)�&wL|]3��"H�m;@���⃁ Qۦ���r��UBMN /���'x{���.��LI�Uz�i��%'.�tl�4m�N,����Jx�{��ꖘ��(���Js������i2�u�+7G���贿�Ik<��.��n	"^��K�IKK׷ @�a�ɘr)����xB���!�]4�`�o�����da/���W���A(�wt,,��c51��@��jtF��}��> �Dy������$-����Q༼.�Ʒy���E�*���Ua�Q�R�yRW>��1@T@}=C��"��Gb(h����=/��WJڣʷR��Ey�$a�T�տ]��I5�2��)��컁�؊L&�Qp�h�f��xP�dU���VGdq�F��E��Z��}FIG����C�>��*���wu���ڊKܘ\�@�M���;O�S��G��6/�j��9�����|����`ϸ�e�Kͦ��z�<|]0{�mTbb�6�&Y6u�?���n�Sߨ&>d���a��ڸ���N���R?�����u�Aa����bW�t�C�B��WhF!��*��d���>xJ9��z��T|#�LOOC@�����34�\��{�x�c�C������2�6�K���5zas���CRq�M�i�2�	U�a|�`.�V,%�rl��Ҟ:�K�OPH\^���nZ^	"���� 5$�*b7[��;͜P	���R-�8���AK�(��$��%��lP�c����`܎�]Un��񪨌뿣j���Y{Q�/yt)�˝fV���BV�Z�;If2�)#�\n[�Ӳ͈wI��ݾ����~�Gn�S��*d��i���8}�KS��jJ������(����(����}�w-�yS5L?'�#v{�Q]d����nѯ׍�z,�wa�Q�l�\�T糏S���{��u�.��}�eK�a�����7��+���E 9��>�o
,j݉� <?�v�kK���~z��Շ�!�r�^����m���������%��ck�:&w*e���S+�$�����G^[mY�W��y��<D�����'2O�s�e�f0�x+����E���	�0	��I�c�GY���Uk��t4��-M�3L�FQb
��)�z��UX��z�H,��m��h����k�,Ù���G�Ux��'���~�3�-=�,gwW�xD��n��g�� a���cEVᦛfW��c�������g�=
���{i��fQ�2�<F�1u��o�_����P��rA!nfT��U��ƭm���!,����$��
L��Ju��:Vk5$����a�W��a户�r
_(�-HB�=��o��/�i�e�Z	���v�w2� ��2eI�#���'<���+��;F�ݹ����%�c��\a���� �C�m������eu���o'�*���Q}ht���˴ԋ%Cß������~ߠ��~�e],��~�U��r���c��E:ȿ�ƞПBr���r��!�j�������5JB7�T���¢��9��Br_�y/,TH�4��侌~���jpOT�?����F�0��������!_�G?i��!!Γ��/t���n����E����ӡY�;o3����"�<0���ܦ^�ս�5�m�>����\�����4�'�e����S��~�i���I�Y(�)`�L�����B�94���g����=&��~��l��W���2�vv�4g����?	�%F���VZ�Ƶ��t��{_�wvN:�ȋs�Ҝ^W��uh�N<�ToP�*B�������QZ�,�����[�H 4il���͵*ƃ��3��� �0mm�A��5��x��P���9#b�x?�m�[�_s�?�\���4����D�0$��I�����id�?�?(�+&������U�Q�/�����]�o�d�x������+dͼ�����0�2
�����m�Y�uVL�gf#�4���$\��ީ���I'xKrvq��S-� �1Y�v��2HV��ٲQ�ñ�]�6�W'��� )R]Z��̵�G9
Z��J�Ff�9�MF��x6������*߷Si�ul����iX��Z�3��O�le�����r�Ί�����'� ���}�h�G_cأ�N��?����C�����-�MYIC|_�c�<�
�2���*�A��<3��W_�8�e�P�WM$/���|���69bu��O�4��h4����(��D7��;�=<��w$���[��G6U!�ښs�_O �����l�fJ鶍�𪏤���*Vc����\���ݕ��C����!�T)�|���Ӯ���� �#�� IO�kϭ�lVլZ�lޠl�T[�7���̦�wO��c"N���^��l�|�7V��uY扌���l��L�G9��H;?'j�1��6���ϸ�-�[zh�В���>��E���vw�YV������g`cdTC��dy��hO?Y��W[/[����Kd[���/g��[�k�[V�b��y�+k� ���
K�-�Դ�&2_�5Mb��(�<���62t���p�����ɓ	l�sO�w˦2�}�-��A�BD�i��l56w�D�`����]������X��ERo��@�ϛ =�+��p��h���jI��-�����K�� CG��QOq���+��O�E[�/��r�[��-�is;�܌��m�b#�m����ں(Xg;5�PRD1�G�k��������0{M�mW���G�=��w��_��h��9T9�Bݛ��8��EL7k䂫�R;�揓�b�r��V�}Ǻ�ظh���[��3��5�@�Ϯ8M��_��;��ˋR�W��,d��L�]2�B����|�y�O�#��/HSg�����Va��a{��I���ć�ɚ��t���9I�sM���Ltt�˓�Xض�����mR���w�����_A��L���t�(E�eлZ��X�]�H1�,�=m����k98V���
���^��3+�F���G����G�ظ,�qC��i(�!����IO��nz�2��ꏱ�쫗�R
���w,���Ď??����7RMz¡�KtA�ڏL�E(�k��I A���]����a������1 [��d2�MC:��X0a��U�eTc���Cw�e�9K��?L��;J_���S�5��>w�k�F ��������S^���>+�J� ׼->�ݷ�Z�������,:�޲�X���e�B��ꌣĕ��w��O�����&�>W������͑�ġ!)w1��4���ȧ�%ͽM���E��x�7+K�D7%����[�D�����o��6.����}��g�)���m��AL����hG��z��1>�����gZZ��>9�]tP:���(��|[GQ��K�x5�d��:8���,߹	f�n\%����ϝ��ft���:��U�G	����:�7���? �I�x�|�U_�`_n�'��Z"��Q� �8R8IG�0c��2v�|x���<��݈`���I��X�������[�2���Y̻���epkb?Zl0CZ�&i�I�E��=��%A���v����Ҽ�@��/���P��>���U[Z�i����}�m\[2kB�\�+��[���mӻI����i�7M��L����xSdE{%%���\���Zn5=��SxJ�ٹ�`�
�y�ߛ6C�_a���yR���0�CC���6^ ���`���LdP�^�^���y����\P�-î~�������8
���kkٖ��v�noƩ�l2L��O��E����wȸ*�-Y����X�㙻x�T���3au�W{��9��U`��|LYeV��t"����z�Ox4{�y�*!"'1���r�}9W ���(&&�@cg���O-�5��S.���r���@.�_�{�5g�L�M,e����Fkou��J�ӎr�!��j� >�F ��(�%�MO��r����K������0H���E�H�����"5��"Y�/j��4 ��Կn�w)�P��%V�9/v�ۓ9��Z7y�%@�� \̋iʶ� �^�Y����%۪^�??l�1/Ϲ�;���v�����ΏNJ>����#+����_�<�9�IE-���f��ny�Hi���U�Ry���%�7���a��d�[�-��w��:>n�D��q�~֟�������������}�]�lx���v�C�PO�bɭcO7��ۏ]����>���:*QT@�c�W�4�S�׏P(�^�7�������2���R����f�)�����#�D8���׍��هI~u\�l����|A#'���/Hs��<f[E��>x_L(�@6�;���wu�`�g���;ޑ%�5��<�Eu��� Ҋ���@B��P �H��3�P�����$�F����2��%t݌yk�ܝ�7�,`�^̍�`�����f�uo��#�R�^܏qk��������\*@���G]�]�=?ƿ�6w�o����dd�UZ���KzJ�H����'�O��}�{��'����QQ/d�������e�> �H{�S9�/?�u���1kt��P?���t��#������)�W&�l��#O��>}���D�GVZ�]D�o����K
{�9m��5��������ё��M�?u�ۙ�U����e�t&:�D���4Lk���x�DC!���ߔ�?�����B���I�c_&T��c*g�r�d�K��)��qB������
{N�����2��ĕ^A�2��4����C�lT�R���%�=�5�`?ړ�-��u�H?�h2UV���z?���_We�om�V�6�Q�ɶ����E�4!K�,����PV�Z8�͓�
W�"��Wᜣ����t�oT��A$���Z:(���O�;̧����X9E2Uڄ���/�K�A�U]��,��r&��8�굎�t;�럼*r�^���yz84>���	!9�����w,�'�\�3>�o~�(��ϝR5�uww?�+�{�d4i��Z"�:�'�YJ���W���hN��?���E�JV'}�a��^�5����x\G��?X0_��W����tB����J�/a���:��l���Q1žH�">�މ�ϐʨ��J��`8dq�IIp�ve��?gU�B���V�d�8��O��敖��_'/N(��?4ex���/V�W�v�zN-���$�>;6�-[�Ǌ^7z|-��΂Y��p0����˒����?�e�%�)N\�,�58C�ihOg,�!��G�d�׺8#��e�vA�ɹ��<S��$N���ֲ~Ir-6d����^i�W�e�'XJ�����Oc�1�#���k�O����< i�3�?'9��'
���Bs>Ӭ�RVIs�)�R�9_ǣaCT���gU�7[�C�����z)k��8��Fۿe(������[k,����ʵ����;}f�����711���P�=�u�W��ޘ|ƔA]���CKE���D�b�\����[՞�1c�˛Y��˖��oY��V�Q�*G�(f����JA�bd�w��;���C6
��@�������s�1q��� �M!��M-�V]|1h�W�q������F�}q�X$��6M�sD�F�3w�XO�����\��rH3ء�#4`R�o��f�t��$b��@��t�_9Q�6����A�G���ҳ�ayCH���f��� ן��$�°���y��Tx���uBR���5�ȫ>Oz���V��m��瑪�*פ&~�.���}�A����;��C��/�fw8�B�_A�^,���dK�������ɕT
�챺����K�̐m�.T��Y�M�$��Z���I�ʷ�.�����4U�f>�cS��`������X�ƒ'�{L������r(��^�A%����"[;���5N� �cp���:�=b�PZ��d�k�-JJ"�}�Yi��\>�z?�G�y��|,uʂ鮕i��� ��x�66��2I�@�?2 1�&�%���_N���eJ���g�G���L�ƆS��-;l��3��/��3�W<Xʾʦݵz�.�+.W�#v:�`^��X4��0d}�gdR��{D[xP�*'Cp����@Kvj�7K���Mz��M�vG����d*��r��E�W��B���ַE�s��n�F�N5�S3�d��K�Ǩ��G�:e����?��:����ۄ"""% H(!R�Jwww����t��tIF����0JJjHlF���^�}��s��{�����s��;�\"W��y0�����<e����{-+ �{�+$�cOP�lY�Z�v�N�G����y�OXA���<x�7;��Dt<&�]>"|��J�׊d��e��)�|�;{�$)yx�T�EhnT=�5��1�$|��0�N i]rXc܄]�t��9%��bp�z�e��xz�AWyz�=��=+1��=X���Ru��_�҂vV�BB�7$�R�����z:�@���J]��`l�EWX8��T��ђ#A���BFB}|2DQM�1������b�#hɑ��5b������sA�e���m�k���y��j-��D������Aѱ^I�A�Sb�dK����e+���4����g�1Z���nΩb��z�?ީ�cX��P���6g�-潟�Ә��fZ#@4eu��{/C���tT�/앓�%��)+iM7�.o����c���O֝?�I=Vw�����|��y^i1�c�n6m�+��3��L8n��K�4��Y����`w�L��S���J��w�`����M�hЖ�������<�)��SX����~C�������3H��LS#�f>fu���
q:YE����B"��v�Q����C����%w�>:�h~�؉�ig�E��P�+�8��o�+��$�jN�0�I���P�v`�g����,��v�y����f7�Ύn'�Z�������Q��E�g5�R���2u-��N$<��d-��z�*�8g�B"�>�O*SaFE��b8+x�b��`Y�"s0���,4��*�Y��t��]7� ˺:I؜�<~*-j���e{i�{35��K=?���h��$�h�i
�w���h��qX�{k�^')Wp���{w���?�B�IJ�����׎N1�7$�m�z��dU�cHڟ��.o�-���+t��!Q$�4tD#M� A>M>R�5�E$b���.s�ćrwv�}c�pi��QH횇5��3�ʫ"{9zN�S?j�f62��㙺
��9
�<+*�7c`4ɉ8�5��k�aT�<z�o $ 8Rs
zY���g(�`S�*��c���� n�FӒoLޝ�^E���R�xt��ϫ"�Dj�����޴��������N �k$�,4����`��O '?�2��pؘ��{_�,��e}��.��.|�x/��&2\X�qG;%���n=��m�h^j:��!����R��P4����f���6J���4�Xu�rk�+n�y��m�q�ln����\��?%�8(����'��kh�uQ?�R5��eא�%%oQ꠵��z]��$�$�ǘ� ��ݏ�������N`��7mZ��b*g�d^��]�i?�i�J'�/x�,��)+w!�N��1�{>�=!ɥ'����qu=eF�"mm;w��'Ø�ߞԃ(�b������}�-}��'�z_�̗d���b_��i�{ٯe����c����dop�Rе7��6| ����4�����O�W�l�ЯFV��A�)Κ��©�����i�rw����!�.�N��)��K"bnw��EUSE��/�6�)�����V���f��,{���;L����� ��@�]�R���Ǘtj��2!l�Ǥ�l�)��������7>�{ʡA�R�7��L��O�V3��o�Ē��9�n��P$����|��0��5W��o|���z� �TE���?�E���Z /7UxoX���Ӥ�3��봏����վ[9��wC�i�%�ה�~����n��pKa���i�h��1� |u?�� ��;�\�GK�#��Ȱ�pc��+��erd��vjH�'fEUA��� 邏�Iy��ب�;�ׁQ?ˑT���isBq�8GϑCթxŚ��	ܸǟ|V&B2��U���_,�6X~%76�/V5�˴�+/�����t����~�<��rPej'�a���S�_��)�C!׾���P5̩{P�~uNi}���i�<q��~�5�׼�ɼ�A��؂��������w,M��^�|q����.�v��,���KU���*�ùM'��#��u�F��^ۨN������J�-l�ui!N�����-԰zG�6;՛�Э�����Q�G��4�n$,�|g{�Z�!� y��ߎ\_�?И?��8JF9���v�)�H=./<��-u�����c�oJC�]|��4��N)�sE-	G�����я�~��Kr��2��~y��!�����D�@�@�Ӯ�uwb52��NWO&~ ���$<#&���ɸP�DS9��46��Rז��6�k�E��3�M~��^�>ld#A�$~#d(Ì�U�=�#?�m�c�;��}���?�J��nOw��,侺l"��Z���,�y|�s�'��^F�^)iLr�� �͎�)�^0E�洀>|�������'�S��<ŋ���M+�L�^����V ���	c����$�������TCo�>p���k�ӕ�_���s|Y��
W�e�@�%��ĀQпn���P��ݷ45���z�e�>��Ws���L��49��e�{>�ٟ���;19fE�YW��ym<�Fkk&�)?�y��m�Zy��wA]|e�+C�=3�?J�����eX[�2�9r[>��Ƿ�����W5;�ᦋ�v	�R����' 2���x!E����^
�$�K����ɞ�دG��٦Po5���h��BfX�V�	����\�xH��+����III� �ʱ)d�����yj��K�W��F߮�T7�^��[(�ߗ�� �3���CU��N��t�,��;�jmB�qi!1I(/� �~�%%����Q�<�wYau��9W��-�8ǿM��|w9uZ��L,�ذ�� ��p��yARoj�f�*�k�a�{������hZ���v#��ɯJX9C���Oe�(��k�{_�EK����Yi�t,��&�"��g}��87j
���~>ˑ�%�Έi�ac�&�V���\�����&��Xo��IV��vO���3�sI�).�(*K%���9�ջE���-aN:l[${���m�����ʨ�3@��D?�M����{_�7ê��?�?�ڮ�.����K���Ur�T���<�R�l�Ө}Y�`c��B{DЦ	m"a��Qqk���v�D�-f���yS���&��?��D�|cZ�5��^���x��w��G�|n�FNܦ��HB���@'�����愁]�[G�Vp�K8�N�<��5���U�'5I��?)dۘ�_U�Uʉ<#����+�?��Q#A|���c"�ӲE��R�c��&�R
�7�b�M�P7�ڮe��כ[�_�Z��y�w�}H�z��N	����Rj����=��c��e�
��B7���N�M�D�����c�î��z�6��c(���r_'�S��|\��uZYX$ �����pt<Ք'�����?9����֑��Z�r���>K�vH��`k���1� ��lpr�B�z�#gy����f�����S*=}��:e��3
�8D'I��F��'$'�B��0\;�����h��s^?����ңk�W�<3�n���nnj7����]X�����X���+�������:�`��eg�w�P.�ͤ��Wp����x�rW6
�g�DF֔=��I���^{��^����!��U�&�d�(�/� �l)�i!��02�E�ݷ@'}�$4�̄��+��T�ɯ���1o<�[FZ?x[IB����9�������؎$���P��;۩"s��n-{S�;���CA���/��(��
��%��>ao%D�8m�&�)0ޗ����'C>����l!���&�?^��诘u�!��m���v7��>Dz�j�fs�98f��p*=�K�N���3��PȴZ��/v�Ө�26�<%͛�OH�0ow������e�%
u�V�$E2����Pd0�?}�͹����-z���Q.�~�ĈUqv^���gI}��`�����;����2jJi�붒�p�ΌU��M�x����w�ͩu��w�����j+(�����f��ք��}}���j�}"�˙���v�F2fYnT��_����3��?H��C`:�*�*�w��Q�~5��4(��q ��es*b^�f>�� ����uN�e6�j�n�!�);�\b��[�ƾ����I�DaS㭧��_�7��Z[~I������8��v��H��E��pz�b)�!���OyIM!�[�x�ᆏ6�Mqp����N�ԇ3PL�
 W���'��(��G�5�L@�AJ��L�1������o!*BU#�T���'Tm�'n���j g^B&Z>o������䰜w�=]̺���w�?Gz�؏v��<��>�Y!d�v2�2�R�H-&MSy�*9`>Ah�ۑ�.������w�@��O�e��=Z`\����h�dؖcR�خ!���;�s��hڊ)������m��z�=�p����IM����H������5��h|+���>������{*����J�0�bҐ�X��F��7JR���KF �X���lr@��4�Xj�[J�Z�x9*3��hC�d�ʞv�NktEH^�F����$�� 6�[s�1�g�k���cQ㾌1�Q����Q�V�� �x�vNΡ���P<3��2mƻ2S�5](�V׆c%h��^"�Z۬���P]�_���qUݍ�
��)P�q�)�I��Z�����[oX�Vs!����p-g��A��>�s9�ҜQ\D[�So�k?�P�-ꆄ�d�<�-yM��������L1�+�Ӕ:q�p�* ĕ�F�sͰ%̱��R��V��"�R�6�G?��T�w�^�[���[���tMoM[4k`^� _�$Fث�Ɔ���$�P�A'�C �qJ����/�َe����]D��Jl�n�.ĩxj�0��cw��H�>�aP��A��
��Nf�j��'�sܿǅ��P�A��#
WC�؈�>S�vB�L'��g�e��r��j���Ck�&׸��ȅ�^;n?�/��0�������_%�h�PR��j�!�{�R s�����G��\��^�G����SkA�8��(+wRL�Ң˦�(������ck�]-�?ig����i؊Q	k��˘o��B�/|Ԥ�&[�x��M�C�V���to�o���z�Jz	璄���͓d#~VZ��,�H���9
�Gڦ �
Z���43R2�GX0s��QG2������ښRe��sZ�4ݿ)_ub#�<�l��[�bnzhmS���P/��R"y���:b�-��QCAYѽ�A*w0�h�d�������V����a�_|�)�5�7�;d�PM�$;NAjd@�.�6aZ��;^��5gc�)��ɂ`��~Ķ���A�[5��N�����-�F����(�F��ʇT���T���;�q��'�PU���u8�Է�@��f���]?9�z��k�F��dx�?5﷥�7�sKp(e�V���P`F�7�W7Y���Ǹ�߾���(T4Y��Q��?��B�"W���]8[�M�
p����qY=��%y�ɉ�v��&r<撷���	�yj���2{N���|�]&�9��;���^꟣���ᆬ����J뵤$�\S2QÙ���=��8���E ���v��D3=Hp��F;�bU�� ȾWn��	�$Uá�I��tI����۫����8|���I�G�˭����	��X��A����=���:�u�M}�3}jm��v�z��G�+��=�daE��ݨ�Y��{�4��4|�Rɒ҅9�l��{�yR<���\ ��r�<�b)I�����0���M�z�(�28�'�U�Md ��|5#�95�������D�Ny۩�٬�c��y��Q��S[S\��;�6g__��+��Wś;����.2�K�����ލ�1�#�	��濋�)��2%��9�q`m`����=�y<�3,��e���o,@�v�j�U��l��Ivg����E�5���9Uk���{RǍpo�8O�\��>|��¥��=k��g�]f��ߟ�t��ʩ?�+�Ul�W���Ld�c�*[��B����c���q
��݀�A�-j��)�/=#��n� ��"�*"���LG���I��g���w��7�����Y��A:���M��q���8���P�A��ӗ�)�7#� �]U`Y꧃t.���_j(�3%��r��"
A��Ԋ���cM(�P����f���v��zx3�p��w�hF����r�\G/=W�m�
�F܏��+U�y OT`����P�ҷX:�>O��<�`Fg�����NE;�j���Ô �N#���A�X`-\Ni�ɈP�P+i��fc�jz�iTg3��BQ#gI��U,햯��l�=�i2I��;�����Ӗxخ���8vӇ�F_�*��$�c��.zjP�V��3����gzd#Iؚ��MJ�������Kr_A�	ϣ��OU�^ ���l�4�������V�^*I�=��3�� ��ҀʯG��1xsb��5,̗y�7��^u��h
.��Ȯ�2;��/XN}a�9A���>�oY��k%!5��uK��._�^d�pt�> ��Io��/���J�/f[7�ָ�?��p[�D�	[����&�I2�L;cJ�	�b(�J��F_Wǋ��*/Vs2�i�-��o�0���i�n^��َ ��mcQܫ�g%Rf��6b#H������_��MUض�Ԓ$�%Ok,�n��S��y���%ny���j���_�A����/vʝ�H�5��` �$�}�i �|���-V��4&���q-��YZc�k��4[/�`�8`�a\���:s3����Y�\4dgQ��J�'���#��k:N�����j�]��!-����#O�`��%6US|������6.[�lb�t��^�tՙp�5M��T|��[Z��t�6x�+�tuJ�O�Fm���cE���$U�x�Rp��9}�j3E�*4F����Rؐ-���3�d�-����HP��٢t����kT�5+��Ktz߃Gm6�!i��T�ݣ"iI�[a�>�?�kJ"��'�T���ԗ�K���?������z�;S~Y�Y��%k.�5-�f��oah��G�щ�jj�u���f������ƪ�3��<��
n�[k̷���6{��p/ʃ����̤�-��MW/[r9qE`��k�y�s9�a�i	�Ri՜A9������4��`�E�P���i�}+��W��K�{AS��Y&쀬��������ӷ����{�<���}�J��Sd�{+x6��{Lr�$�U]�$��'/������:��!���P��W�'Z��O�e��1��k8Y���<��hvME7-��س툉�)Kx���KC�.���8dϝ%#=�:���-`4J�g�\�~�fr�X���`�#l=q4Ҿ������U [7�O�v:n4U4 ��_��H�1<r�d̈m�<Y����� ��Of'
�ia��YA����<��������L����1���f�R���0�mdOVMt	��)�>k*�hu/p�{���#���B:
5��Y$A2x���<������xTtn~k�+�jZb�2A8˷�̭i��6��N��\�H��SI!��f z駫W$���	���FcG�~6�4r�F���u.������]���\W�<���i*�\-�^iԋ��9[S}m�d#�}��Fq��N�����Ff56ɻ��yw�i����z����������Hs�t�/K��KJt�����$P��*9��
�A�����Sg�|ꭼ�/[�SV6ڀ�'���x}����ɖQZ�m��1;�9��	v���+��Fd��4 ,t������.�����;m�,F�w�jB��1�- ��5f�r24XN�|�_ּ�)s5q�`r$��c�f℗$Zz��Ȉ
Ľ��Rߑ'������}
7����ӧeM�������i�%�O��Ԛ�O�9�7m��S�^�.�=o���X�R��$lLQ��rZ�/H�]� zyN�?�z�����~U}��@�;�8�;�S��X
 : M5_c(X��"#l����Ny��Ue��Q)�{�@���!�rw�ݧ\D�舣�����7l��A�������-������欔�����d�E�$��<s5z0-�<oq�G�������	�Z�Z��R���9l�����2�����w݂�H�䪃aP�tWp��c�˄�����I�1�\B�FA��9>��:�o:�B�@S#x[��F]�_�J�.���������  ���'T�$J�>�I�[���X#��b�G��o=i�aٷ`��)������)���?#���xK5�݆ۇ��_�������%Z�d�s�D�_"ޫ���r��U�Q���u�i�4�	�)��Z�l��C/L�L���
��m�pWG�1�V�!�X�k�֗�{�z4�Cx�Q('���4��k,{��^�4/x���"mU\��-���\`d��s?��b�d-ץv���.��R���c�4~�j��Z��M�}(7�3�֥S�O�|xS�.�9�ҳE��udr�@��7��ۗIT�s�����>���lJs��ﳢO��2�s ��L�x�<��}?h�%��к�,�$���B��C�>3��2«s�F�D̈����a$��=D<���8���}ei)p���:	�"'�fň�j"!��Y.�͍X"����c�[���~l�����ȶ��ۗ=��-�H9�rL'4�MH\�R�����C�*���IZW)&8E�$Т��ݨ�m���sģM��q��:�>]kK�s��r��;j7d�3*>���ܤ�F�7'�{��4��7����sϞ���l��1))X��wX���_�$|:N�2�L���g. mؓ_I2��%������޼WXb�|�S��o����%���b"?��f�RR���9&;��G~�:�FO�Kك������.���Փ�#5?䰃����{&0+�y��jyPl��y�Tk���n�(f\uy��ʭ�v��.�愇s/���rj����7.�\_43BFQ�9��� ��m��H����z�4���A�(c�TDJy�)�,,�ٟV�>��c�k�ħ�"\�m�7fjz�.{ӿg�y`#ic�I#�����^.K2�?%cOU�fc�����)���B-'���0�4����2#d����H�Q4g���P�%L���c�?�U>*Ucl���fԐ�UO՗���(�*���
�^�d�;����T��J�HM�˓�I�X��8�hq�W�ލQ���$���8��C�n��Qm'��1�^���,f,���U�E#'�@�Ȝ��,��U���cGH��G�I���Y�����?�<�l��a��Z
,pQ��4X�LK���r��w��\��bЉU6��|A*U�y�����z�#�%c�������4B�w�ktX��^Zs!���,��3b3�յ�T p��C:�ܛ1�^���?W�ycw�
�g��3�:!�92�@�����F�,�*5Ph��DƮ�E�8�Z,��m� �.nj0e���G���@��hr�����ͱs�^K��wp�D?�E�Koo� �&d��v	gI=���2���������+E�Z��I��Y��*Dl�crY�o&A����>C| w��H����N�BI��ڊ�h�T>9�1��5���G:��ιɦ�H�����3�%fzG�܃WY�	�J�b����2�?lP�UQͽ�O{�'\�� 9ѭK.��;�X�n��s�6f=�f�3u����J�A�vbIf�j��B��4�Ϟy:s���7*E�de"�H8���69��疶���ڤ~zq87s�/��y]iܮd�<�ч��?�+2U�J��@�F�IсҌgI��U��7u��R*����W �m}��F����n)f��#='1��$�m���^ϒ=f?� �l{���ʒ�hB��%"�Z_���[�	�J"�ĮQ��CY��+��t�����
��\S~��ɮ�`�>�=*�tYxM����i�ʴ�! L�h�s�~��*0�g�S�&oG�6R�漠��������d�dD�j|Y^v�t�ύՕK[����|�:���r|����1�+O�)�޸A礲8��È�X&�E��P�.�~R�`�s4�,�}�_.xքj��ļ��Y,�{��)��a���M����}�㚲���-��Y���� <�6.ܯ
�nwM~��F��"�l	~�8��y�|����6{t ["�9��{C FA�+���9]��d'n�]�$O��2���U� [o
@�b� ��OER	ʞ�T͉x�y7��8]��>o�r��5��k~j�eO�S��z�>fP�}q���Ze������Z�k�b��#����;�E���4���|5�E)����F���wH�Q_��/ȳm��@��&�L��L�m����Gó��G�k�蠪���]��k�"�����L�W���![�`�����Zl&�p�E�|�/��tB(+�|�z�U��>P|u�@=�����䨝��\�҈��ù�Lv�K:��=^�l� q�s�����<4�%#�&����-��.E^����������4��8H�P֪�O0���WB7����*�Le���)pf@u�M;��$*҅w���j�5���T���=_�6P|i�4	2���*��ҁ���^�<Q�R��;H���ϳ��Cj
=>bn�A���.9pᛏ������'�Z���Y�і�JL�l���R��)u�o0X��p��w�Yl��40W�\���Pr��<������5����������G�}��N
#����Ǖk��y%�g��?����/���pӬu�}zM;U�fp3`������$c�z���.���s�8%#��C�;~�{�㕑y����Q��w�~�� |���,C�*鴸ڔhI��v��<%�G��.A��(��jx���*n�h�Ƴ����*�ʰ�ɘ��]7�+;��̫�~�}A�Sv�tM�K�C�S2ش1?�M�m?�<�����ɳ"�w�X�=Bڲ軜�)�~d�������JhC�cp��ʾ�΍�W���w�r�Y�*w�e�H�J���T��/�+5n�ܻp��N�+<�5݈[&��;נ<M��!�Q�%F^����������,q������.��m���ם]ҫT3�ϰ�*�4�X�����(4�z��]j�Ii>�T3 ��mdNW�����P�����.��=�8�S�N_�\�d2���O���ٚ�D��7a\�L����s`���K���o�P�As�+��ǭ��Z��k�}�~`e��ޅ�u%�$]ҸD�k?0�Ѹ�K[��������9%1������-P��b�G�`�w���8�$'p��2ޛ����%���1�Bz)��}�kX,:�pM�ͦ�L���m�,��t��Lc�jfBb'���ſ:e�����������w����L	(k���O6M^W�kdks㵴G���������
'��Wq���mpy�c�-��=�����pqE�W�g 2�>�=}�����,f�i�_n��*'h�m�HH���r{7|�2��,��xN�
uB۶��4ż�5�1�
b�f��U���yx6����;^�4�#$�՞�C�'rYT$�k�_��c�S�����DN*�k���gm��{��8un��m�q��Df��s#A�'=+���>���;3X�.֚��]&�W�7�5"2{���i��C�;b<�Qv��q�'*;3c��`�⶗���~�L�|�N��Cܕ���I�\�/y0��W#�̠�
�}=��R؜��E1Mi�L~��"��T]4h��;��f�4}E֬<j�x3L����_M�;,�˓�ʛx���~�yw��֦l-��V��6����R̿O����P�;�K��Z�1?��5Gk�ύT"sۊ}��
0e�H,��Uoq�
�K;�di��'x>�Ii8
eA�P�x��J�2��â���Õj���Q`#�Q�~��h��nG�b�=�z�0Gֽ �C�+$�ɀ�W;��1�#w�S�q�eT�e��x�����6Fe�47B�0���-L��T���������<�k�+Ҩ��f^����!�-��J)���u�تϾ�ݬr L�o�ϰ��[��@��D�m"�㘢����?���S�Y�r��$nvTs9�h_��B�F��m�d������1J@;9��2�{>���

��k�$#m������6��.o�W�`��uj:�\G�O�l^؟OgK��9�)��r���ʨ�~5��u�z�oxG}���� �� �>&�������F6y��ͯwxa�����ʞ����^n�{��ϊ�'	4���d,��ZmF9?�v� ���ʚ7�C,����X�\�T/6�w��Q��U��p�����1�I	��`%��xF9F-Q�̂�ɍ}�W�b�8ԤC��^.��m�������#�x͂j���xjܚ�����
���/v\��i9���-P���fw=�c>_y|�ƈ$���7GY���IN�g����3ƣ^NK��P����L��n9���wV� 4Ȩ#��r�j7���4<�e�g�N�BP�W�B�@�o��c�� ~p�}�3�J�6O�������z�l�7=�/����6������Fv��KF�mI?���|J~j�+Cy�2�x	���3�i0��+�$�e�CL�C���^Z���Zhw��p[#�j�Ĳ��e>m� q��N*�8�q�4�����(�qE^���y�r�>s#�e�)���9Z�T��W�%��&ı���g����Q�~+�����ݐ�׻�Քy���ʈ�hn �J+��J2~n��B� {IҔ��Ȉy��CWЋhW�Yz��	���2CT�EPm6.%��.#s��yK��^��A�#X�ҕ��5k�(��-����#1wQk:4�ݣ���� `IlyZX�{����}�3ƏT@(I�q����W��1�I��>L��捱u냔0��d�x-�
0���'+��O�W��2�غ�'S��`�s� �Y�!NT�&^S��<���kJ���nB=�@�$&��#6����U��lj��aq�0����!�F;y;��5�BI'r����F�z��9S�+�ʑ!CU��ߘ��~�A�K'��W��3��F+~ ��ޙ� �(At��� G33&�}�S���'c'Y�,�9Mu�a�������G.6J������r�|G�z�mc�������3@������D�?O�!'{����~��9��kQS2�����e[:n*4I!�5#n3#t,���u�p���d��\�iw��䏞Y�����]���H�w����o�O��ѵ|GL߄����W��w~H�O}0�=o�6��W�=b�%���J��������ZG>�pz6�M��G
`A�)�R�����)35f��ZI��������� z>��l��D�*����򟠳0.���Wj�[R7��q�] ����FF{xnP "��bm�=�p��<ZS(�z�f�kR�A�5�3���CK퀬;=
H�Og$J���1��4jv�{Nd��	�=�ee�0�*y�xO��	-Ŕ�urd6�K;�v�_E#0�j0�dB�&qJ�Wf�^4��2Z�k�1f��ߍn6��x6�Q��*�ʸ��9���V��8��3 ?qT>���}��N�7\ɪ9���M>�.$���D�����w ƃ�ׁ;����l��l���,܁Z���t�Z�Yl��;ea�bv�#�YX�I~��.*3��o�;��8T��w�;G5�7��
Zո5��Nn+�S�~=AC�Ov=ߌ܁ݽӴ���ְi���=Y�i.������f|�l#5�`8�}q��Rx`I�j���KpLj)Z�ߧZ @�u
�P.�k*q{ّ��V�]�����WV�_,�g�͇���[M/���I��+~�d�Ù��5밸p}��a���A	��v#�Jמx�ve7�7��`�,z��u�#d)�ˌ:�w%Q�o�̉�f���{Y)k9��lG�D�t���.�R���0]�q���7fh�G;��b<�Z<
+��k1dYP5qK�)}��,��)�y������O���g#~��q{�E��}ŎU>v��������l��	�>g��sͧ9 ����R�}C+*�F]%��Qc���z��-`Xg$��t̄�'%v�9�"� �"��%�
��|<��"�G,1Q�ӈ�xu��(�׿&ܲ!��W�����g�!��yh��hox���mG�)�N[�B�� ���6��o}ri��V��r�@��j�Xߙ�]��Fʩ�|�IwC�\9K(s�[�	4����v�x%�;�1��6��8\5�cx�"dNP��!Ϟ\��W|��?,D��ؤL�ѹ�G�5/K��Ȑ�&�n��Z�1�i��9Q���!d�\���î��&�7o��R#�4��#+������X|6�C�YO*�L`ln��`/�T"C���4"��c�L&��Xˠ�z���e�âq\1�ȧCsJ�����n�������N�&]�ZN�*G���BJX����T,ѧc�{g���J/P��li�=t�ыgb���
j,�[���=s�7�"'��:gm=����;�m n:�%�?����56?��2e@	v���<�W�� x��|\#gx�jn.�R�� ��:�U�0;=6kZPɢ��������4Lr���딬,E�T��%���(럻F7넜,��@�E�)�'���4^w�^�z��h�x���^�00C���A�Đ�^�� ܇3����k��E��M��l�|���H��O/������~xcG 54���g�jl�ļ$�SGy�ƚl���槕w�
������Ք��=�ے~�F�X�ݢ�}2��7� (4@�qq��>�jJj����d�;���N,aճ�iN�!}%�$�f�;����w�I���N"�h�s��}qp�Tu"ը��04|�Mh3���o���@�}PԦ>XXe)�:���즻q��$7 �CI��n32�+:��s�_�e$�k8::�!�j���ky�y�*of8S�!w����s�?m���ز/ ��r�z׃h$Kgf�mB���( ݿn��Ej�cQ��x��߰1� �]�@�~o�r�;~�A]���`A�sL$���s���BͶU)׮��o��G�Qf�Q:��âZc��L�i]gNQk�\�p�ӱ��䶂�`�,:HM�_�uK�ȝ����t)�(������%Х�
q�y���N�tʵ����z7�*ܑ���~�V����5�Y��|��>ҍ�3�na�������M[m<KɆHݼ�U�RGp��)I/X��,��x@"�c���$�ޘ�ʇ�e�o#Pe�V��Ў+�~������]h�%�f����Qk`i��(j��"��H%��3{`I��/���ԟ���*����½�5%b�ۧ�jxR,���lK�zh�}��7��JZ�^�%�'�Y� �"^��A�Lm�ΊU���,��ՔM��wY�w
U�nD�X�v��V�WE�pw��|̷��-?��O��1;7�꺝
+�S��^��XE:>�yeC��Լ�����c��[�)W�pwfr1�6����*���.��-���-8��U%�!�뤺���{�R9��>��#A�Wu���������E��O��2��J��g����M#%{�I�}�f4����y��rE d;�����5���R��t���]/J��[�|L�pr��2�B����Z�m\�LH]�j��~��b&��๐�A�G˅�$�\��c�G�����?���͡h�F��ǌ����t��W�G^��#��$�,-|�m�� t��ņ\L�y�[O�G��%����ѭ� ��ܛA]��J\Q�?])ܲ͆_���O��t���9���1��qlxjY���y=!�i��~h�$#�x�M���9�tyJ:�������c�B��7B���<y����Ț3�͠»�wmi���m�ɻ��>�^�U�2�%z���v� Z7s[��,�b�7��-��(��� ��
��,�o�J<�s%򆧊�.ѺAr>�포���(�E�T#-��ooL)���I�k��R쨬���R���DkrdZ]��j�>`��/�;6&��U�xh�Ы��`� ���cY�>��Yk��Ŷ�'흞���^`���t�=��z��¾`�����i�b�� �Y���~�97��>b5�������c�s��9l|�����4}����j�N���	�F��p�b9�ަ��ν=���Ɨ�c�&>la{q
�q����o�i;�t�i���Gӑ��ik��7��ϰͣ���ɿ�Hs�mD짩GL���JH|�3/�W��ʐ�̪���Ǌ!7g��fgrɚ��4>}�Vèr�9˪���$���))��05�ʳl�W:J���n�Mv]z���J>�g���]�\�:�G����<�����%��h0�2�b��j�FJ'GjV��V^~�������P�be��-Lb�e�}�nSs�w��h|Q���bӵ��f��s[N�eͧ��	$Qr����=����u��^����V�NC�������C��س-#J����T��Z�{=JSj���!�մ�B�bLV� �Ƹ1����ˁB>Cơ���q%�h����}���<�.�n�Q�qM�1�a(�TY���T�kV3J0�xԏd��+�{Ķc^�O��!��d8=8�X0�1֤C/ra������6zaH�	�:Rc��<��nK�}�wB��P
��YL����Ī��=\�����dcgZ�{������.�V���+r�Ie��=��oW��Qa4�M�~�7�7Ydz��6���s�S���+d���D�HrE�\��\�RR�}��ܷaX��r$w2]���嘈af�#�6�ff�[?|���>���y=�����ߡ��ؔw��|��=G���Ash)�����{A�H�V^�����+	�{��}��(�G&7":<u(q��&~��zp#��o�"]m�&g}u�5��/C�q���~�U��y�s��3^R�Q��c�_��胙�<���༙_�y��f)�+�U�X���0M�ڿػ7ΛO\.�%:V �)2������۵�
�F���T�9��c�:�x[� 鶌��D�uϴ���>b����j���㯯�g@�]�yj��"#��%���|zHz��V���f/	�Q|����x�d�+)6�ɲ1�  $)a�-��Ź�<�̹��5�h�@�ٗͥ�@t���)�#Y�;���:��kd�n��}�����;��pJ�5��Ό���]�g4t�yЭ:���"��Wt��U���f�u㍧k�������%�(����T~TV2f9S�'�'�&����/����4H p�*�G�L�uBܯ���ħ��������Ԝ
����?u�1����@���Å���L9��-��ȈG\�>_> ��:p��E���٧��	��`1�� �nj��H��L�s0�1(�Yr�MHx�@�㥉	WE��P���І��
�ӛ�h8-������=?�3+���)Z�Zu�%����ڋQ����G��_�7��@���u������\X�%[)eu(�Y���٧������Z�zO>�|'>�D�'-qC�Q[�R6�O��l<7v�z���రw^U�1�Z������c0/G�hsr�c���>V1,�@-l&��ڡjR����L��-��D��͝�9uo���
C��J�� �F���0�b��m��z�1f&��"y�u���ӗS�k�,з��R�sj�h8��(D�a�����4Yӻ�Of�a��AA��4����o�5����5�ԯ�-�s�_C��T��1�ƦVT��En���ȶ��?e��A��ǃa����2��N�U������n���z�eCp�6��q��cr����/W�.~g�x��`^+�ܹ]Jѕ�9��Lw�ٮ0�Jy-�?��R��D�2�&N"���OC+�*��Xg�����hx��[��[�?r���!�+�.�vÕ�@���(��.�8��E�8r9ƻ���5/-�4�8�WIl�Y\�<Tr���So�q2��������R+(e\��PS��mB�_��\��'�_��8�?2�O��4;�U[�˹Z9?0X�iҟ�����F,�v1U��O�C�=:}�5��l�L|)e ��g�B~Ii��C��=����d��/�ϱ����Ft��>%�!�
2�;}��-"�v����Kw?ݵ�lm�\P�$tbi�̿�Ay��������r��Jb�^P�AD��?��[t[��f�6Q�a���OO� ����1(���<�N�sba9g%2&�8��JEm��&S��0�CU�aJ����G���:����g�rI�	��������\���F�[���s�굦�k[������
�s�Z�/��cvq,���Tx�$��c/��S��@���~��o�K�}u�<�+/ӧ�F`�ެ|*�sT���)��Ϭu�T���
-�cx��pק��O� ��{yS�fm�z��d�n�OT���/��ݷz|����I�A��k@<#�b�>i��/���1#���/~�?�޿���jb\�-~֥E�-�\�=�J"����%���,�eT��b�xe8���/�A��>�3�/�aF�Q
:��z2k�D�b>Ӻ�Y�T-�ue�'�n͹�lY ����S$�������(��N%_���A�C�N���r�������`����¼E4�l�_q��EM:f��؆��@����3�9���c�T��5���<+lYx}2��3� .⋗�I\��`$ 9d����'��#OSJ5_�%���;?�I[_�r��[ʇ�r��������e�I�\Dh����c���t%I��_��j&��T�f�T�St���wZ�gܧT24�u�����}���j:�N��j�W`Rr�ܞ�G˱@D��:7o9���hi���|Y��C�d�ˍ�~�o�����X�'��t���k�����5��@@�����S��D��OL��W�羨̓�:�i��ξ�Z��p�/��GA�X�u�̊'�%��=�l��}���g
�}�:d�Dg�����,��dN�s��M\�
H����O�����km?_����`��#/��mZ,�����3�N#�Q,�i��$
���I$�wq�
�t� ����r��6�k��fQ�� y�*f� ���4Y�_F'V�DhB�\v����Dn�5O���6n��W�csX#ޝ6c�i�ymFO�/�(��羲nc�&���;���wGs�[v�^��&�;
ڢ�]�p���CK[˗\H��z����~%�������9���8s.m3)mF�I�t�����c�ND3�(Sz���is��j��5��u����B��F�%ˎ�Bk����{:�Ԩ̿�4�UM{�FWa/��bO]���q�`z*.�(��8����%��G9M,�ة�����y�!�T�2���h��3�aΦl�`^'���
���oam5N������f(�w�d���
�{徔:��VR�f�@�'����S1����T -�R�����S�"��_�+s<����Р����]1��s�U�o��s�;|W�ΕG�](�Ww	R��{��%Z�U8���-�8ر�*��v���^�Gb�Um]���9��\4EG���}��=-��k��6����G��+wͤft�[��C�`�S�ȩ��gx��>n��a�{s]�rǺ9;l�����)�O���.��!7��8���C�v�����Z��-ry�Ledd$�jE�8���9^����cZ�~�/+`���������K�������[�(�,����c>�������/E�N9:v�0����Y����A�$��bg&��3f��%���#[�ˣW�$E��wB��Z��R�%�Ͼ�ls����g>V��M;x��'��K��cӨ����a��_�$�����@��`�.�oW�*쨉?j[��A�f�)�c���U����Fr|k�z7c�~&|�����U��C�B��� ۧ��u���`��H��N���.�ѷAy��%m�DoȬ�^ȸk�u�w(`Ulg�r�y���I�z;�/����{C6Շ)��$/D>Xg�n��Mx�v���G�����G)r���y `f{�����w}B�l�������61��q��,���;�yﱼ���㵜y�Y��#�ֵ�f��R����|�ޗe�R��>���O	4		;�_I���1@�q!@=��gq�$�����
����}+��鐎!��
�};�sެ�������o�J�7+3��� �_<��������8ǜGq ��}��Lmz`�`t�|T�́Ul��Hm� �Е"�$����Ϻ��q�kC���,^1ɇN�D��2�7m��m݌,+Y'笟!���b����[�"�z���w^�![V�.�4l �yC����+����[o�o5Ӌ挥4��x h���������>_�	P������A��Ϟ�ѽS��� ��������{C
�%,����_���%$*��k�	v�]~Ӂ�����?�3���H��L�=F!f���;�������ã�y�x��K�O��g�Z�8U��x_o(W5�����&U�����SV�@��Ւmz�+m� �Ǌ\�l{�~X�����ݐ�!p�'�៎b	�2�g��1�4	���IT�A�{�dЍ�ŷ�n��Ӯ��Q�&|�5�!{?����ܗ�9b�7�~����Y�*I�#4�W?�Wc*8�]�$������s�.��s^�ŕs����%1uv��������W��ǆ7��]_!��">����G9h&4��b5�DPs������� Lդ�l������ݼ���|�gz���.h��l��}B0�w���<
RKc��Ŷ/�{�����!m%*vX�rg_�K�Br�q��k��p�#|��\� ����{�Ӟ�v�H����L�Z&9cpH{7U_�E�3�W������#붆d�/������hf�k��[����!�����L����v�]d��x"b���W�q|,��X��GJ�Z��U��%5�ҫ(��������*����-c�|-������*�J�X	��}�5�l0�G]���Ϧc�d����Q�?���w�����c�5�Y�?���w�ꛟ�̓�����Лqa?酱�V���_mp�1��@����� ʆī�
v;�:�3�е����!N�ٶlJ��
�x�$���Y*���ӄ������ב�um�a=oɠ����~���n�V�t"e���}/ھ4y�x�Z���#�w$j�Q��:j:�
ũa���_�mO
��a�GHW�W{�Ȱ�YbS���R�|U�����֕�JQH~Rggm�7����9	!��C�(V������A0G�3T�r;yy5p����g3�"�D��Жv�~��B՘���B����h�����]K���z- BoBI-�L��[tI:�9�i���p��8����^�/j�d�����������LŤ)�j},���N	o�ψߟ��h�k|NBP���f��i��C Ȇ^���Pvܸ[��#ځ�竰j�T�+�9d���=�3p�d��	i�ހ�s�etѣ���+箮�;Upa�
"P��������{;�<vt�_f��$=�i�l�4� �Ç��k=ܛ��(vb�(u8�)9�VZ�9���f=���ߐ
�ux��r�"����0��;e0�	x�|cx�\�릟YW��ܗ/�6�����7U�R���ח�}�N׌�'od,�v�a�eyx�\��r�F]�~��\]B��ދ&:h���� �����o���I�"��O��8\pł6�	D���y�/�Fe����tI3�{qa�<ETQ�[��������Cn��r�{���q�ȕ�r�q�)"oC^��}g�Pd�Ɋ�2���K�ОqW����ū�֩�
N���W"�rU�Ab��$���X��iDb�^Rń㶟E��NwSU���u����7kȽk�jr�RJE�)}�9^�N�&��?x���v2�/��!��H����p#;7;���f�*��b��c��
��F�G�<?�tU�:ω�gxF
������~ r�^�N^� B�H�CHE�g@��op��-�C�U�gd�ЖXƟ �_�, ���!�h]ٟo�Z�(��v �G���`������_u������4u�d�`�����@�Ixk��9��őrZ�e�n^��_��T���f[4����eY��h�_���PF�S��u?��S��k�;����j���ܮ�������+,(M8��W�f��i+N<�m�4�o�|!Y��]�PzWvt��d�N�q���r��3�e�֮H`�f�Eʉ��9ޫ����=�6��SN�_<$��;i
�v�}��k�r�k���m����Z�O��I��;���C ��*l�58���^F�H&����}z��GyY9LUq�%:���r��v#�d�FjQ��/�x*�G��b��Nv�ߗ�?���ӣ�!/��[��܏�;l�������2a������+j<nyr�5t?���o{�;W3�ы�1�Nwt�l;�ĝ����- ��BR���`Z���ؘs���^�գ��i�B��Ȼ{CW�Xd�+�d�������|(m�]l���	]#��j�|��(Hŧ�/�8ZND���~��^���s�m`>��7�h��:��z��R^we��{��{��*^�'���2�yW���f䇔s����U�uxE�(uzp�h��wZ���1�w�7���;���M{Hծ��^�o�r��Da]����1��(,������y~���3�?��~��Fi�̵���6�-^�4�';�<��Cwā��5������ a��}��f����d�f�lU�4T-�8��~�̵D4,�9���^���7�f��%�x�VZꖅ�e�2����%0~�]�5���p�~;-[Τ&^�F�SIAw$�j�N6�+ϭ�S�_.�O�vifWT1}�0��?]�avG�,��r���g����8�v�w}WlZ����i��h����k�í�iɤ��Ƣ a$j���׉g����A���?5���}��A䇗ɖq�!�H���m�eb4oF����8�ba���������Z���bSSn��Ru�4z
em8��ۦ�Z9������/��S�V�~΋Ȩ �ڬ����L#}��"U�$�X�]���D7�¡�� �+����嘯x�g��.5L��NLY��X�%��;���6|d!X�.��Y��#��M�r��!�J{M/���`�u���� �����'�.�����4�Js���2�C&O��	�e:�Y��_k�/X��@�9�"Pd�f{��V�s��6��@;T����4Ax�U~�$C����xno"����JA����n�R��*�ϥyI�}x�Y�mIj�{b�^��	Z�
���`x\�/�X����,�Սv��/|���wjc���#���Y�ġ�<!�M�����c@��n�F��q�իp��1�����iP$ߔ-* �w�Y����PqH��Le��x��5�����k*�L|��Ђ�q+^6��U?��%*�+����F�q}�Լ�ݮY�^����X�<Q>$����]ZNr�,^�9��a������`���^�=|?D�Lsm\�����./۟�@�|�j��,��@wd�'�CǴw?X�����A���1�3�l{ �`!��4�XX~R�pӆ�z��9�)n]�o~᚝�JQa�_�I_ʸ��mXZU*���^WK�]'�#k.u@���f�>cv��=݀��)��vC�t�s�3+�ӯ:y��*��B����k�����̨�[u�g��Y\8ydf��( =��"��h�oq�F5���x#�5������ a|M����K�#)M�v���1��̣���]a:��%m��3C�ԕ��9Dzx�R�.{gl�1s{��q*zh���lz�\���Ί?�����-&�<���쀷�Xt ʗ(�Q�[n�����l�Z�Rݑ˦δ����Ί��Z*N��L̮_>���vFs������j�
���U	��#�!e:�`I��g��S�Ӂ�[�o~���fC��x	����$�)�5�+�#W�ƥ�x�}�����r��E����i���#'�ģ�TW���Z���o1f���t�3�5�|����E9[��Ga1ؗ��Nm��}�G�>$-q(mK�t�1�l,�e�i1�í;u���~��^M��g�����)�8���������i���%0	��>��u���[�!֟�� B�ռ4v4S����|��>��Gx�$��H��m����8�#T��D7����4��"WC~�m���Ә��8���b"W�>�RW�[��A�BK�UZ�_�Δ)�:��P�cc�.�^�{���$Ԙ�,|�E��>�3M�ݠ\�}��Ӳ�ϡJRs�P�^s�O���?�� �ċIbekm��:֤�_����$��4��OmK�t�t:m{)	�#��X{���Μ�s�ƾ:n���Prh���J"+��+��j��z�zT`f��=0�5�y�|�[���n��0(�L�V��+Y%�O9?3�qi2TI��ͨ`�ӄF�7�'
�`ͼ���"9��🡾��ǣm��8|��(��˗��o�v�Ț�>�𩩹pXL �q�x�۞\R+�zi3��,Y:�f�#j3�8���L���/���+^]����.G������}3��ٱ���E}Ǐ|�F�3|/�{�9j�S�'ު!6j���քJWpY�-V����a����׋1�<T�?�հ�Uԉ����J�����`�XI��`���b�P�|m��,���p��CO_�@�!KA��<��'���h_����̭�����nj�����P%�릮��?v�x+�iI���v9^Gݹ������Ƭ��(:��cݶE0��{�ҕ���X����j؇�Y!��%F����E�:��d+�ݘ�(T�{>G0t�n������?���&�տ���������y��;�5g�N�RR�j��g�@��O�������4��C�h�U5�����m8\�\V��y'k�����.נ儞�2����)��W���$t#�0| �7�CT���[��kk���n�l�{�$F�i��ʰ
NU@?��H�T*O��>��v��.2[��I���ؐj�w�B/~��"�]�������~���8����}�c���/û��Ǐ�`F]�P��=��~��3�a���8����j��j�Q�o^��7�%c�,�b���͟�'?ܮ��Dq �B[�:	�c�[�k�u65c����F�<;7vV@f���uN+-d�3��)ķ�ʜ6a;���] ޥU���$�$�+��ws<��9�q,4���~�W��G�W:p���1H����{m��T�fr<�[��|��ϱ[C^�@�>s~U�F�v�E4�Ϲ�L�y�.Z`}7���?�<B�v�ڰU׀Y5�1�����a�	�uG��I�&��/��w!�c_��q[H �0��w�=�\�u�|=�����c�r�w,����	D#&��j>�(Tr|\Z�g�	�� G/Gm�[��,y�dL��a�A�����ջ�G����B_"f�6���P�Na���Nc��i�̭Jg~[7��{�J|��X���dQE���Q� �ό�nv��c���&��#��a^y_9�|�;l���:�>s7�{�1a j������hn<�S2���5������(�t��	��?��s^�D���SA�nQ H��}����+�l��Fm�� 縰@�(�<�	��E>���1D�h�ڑ��x��K�ѕQ�P%���̭��4��y/��[&�C����[�ږe5��t�$/�ѯ��{m���?p{���M;��	��d�Dtt��r�"sZ���#[j��x�h��s��%j��eyF���w�����ֵ|4�d2sƽB�ͧ����v��W˩x���X�p�K��ƅ��P2ie9A/��?�Go��!y��/��&'�����d��ڿ!u�4�����{M�L���o���(>7��/b_���Wďc����~���i��N�[�zu|�1�W(�]�Q�Qӫ�D�魍'�}��3V�,���d#J|�mU$��|��uh�Iy܎{��^��G==���sB��m��"Շ�b�C-H�՗��`�K������=��!����Dww�Xǿ6s>� �<:���Ǚ
��!T+H�1�z����Z(Д�U����U�Jɶg��,��]=�9p�$;�;WÈɝ�WVv/rמ[�V ��j�w�y����'�
9����!�fZ�ֻ�7�N*�M����H�7:���/��cM�R_�cg�/j��r���6�#�z
-K#x�u�~�L��1rBV��H��S?��3Ԝ~�@.��qk��NMa����l��"�:�n
OR�d��s���-I��Ӝ1!�þ�{����|��i�[e�����d��F?n3����a��
���Ɇ)���.���:�N�����$�H!Fv^5;������9�����:�1t���FP��;�sY;[��N.�I�'��ޟ�t�Xԯ�Yu��j��]����у}��TG������X{/��+qbCdN�/�>L���k�{��'a�� V�L��t����R���ӀjN�2Xߑ�^�����M��F�_�:���R���.(�'&/,!��]F�|4����0�c}�淙Rce��yK�Ly��FT	(=z�2�u��R�T���~#�U�F�7L���ΗG�UFXx����6��	��G��~�'%�?d�Oxș��j���?Zx������N
^��}:��p|�Ch��`�h��;�%>�7����ݍ���A�q���3�Ѧlb��~` 
�h�(�r��^�c��	�P�,$����u9|���h��������E�^�3�A����K��#���ٻ���S��F_���^}��,)npkh���7f�X@��0.0�A�y[��l��1��UC��2��^���eT�b�5�0����'H�(��X�Z#!?����嗢F��ѣ�{#Q�k����^��X�J�xJ� ��Q��*�=�vP�`�I��)�E'-��/K�Ӑr-A�H���� �������Xx����
~�Ёb�u��B�A��{'q���Yn]w[� �Pp��s��n��pp�{j�yTH�w�����0��[�6fJ|�c%E�����>�f%�����60Ɖ�����k;�-8ަ9e�gi�Z���	;׬������V�I��SC�s�䏚�������|R�{�B�K*
��C'6ڞ�#����ns���P�����V�
�\�^�F�Q�t6
�iO�<����Z�6{�mo�gT���}���?��\U�����X���W���{�$��RL�35�V=�����1�(��apnYx)�Gmp���^��X[<�{��2�v�����M����u�����~��2x��O��U�?���st�*�%.v�����݆'�c��:(�M�)�^�A~����ݧ왛�>�V\`�����)w{���"m�pg��v��(4�����~�,���=4Q�o�ĩ�Ю�|�1��i�Y;|u���IJCyW������`�g�-�$z !F=��/�ٗ��V�0;���kkt�K�}j��܉r���<n��:�����Rj�ٟ_�#K?����r��gG�c&��l#v��[��-����>�oN�s��a��+V?Q�,������Uq4�=�6��l-<ߕ��`�~���Ã�lA��8�}�ECu6!�{�����<�_.w[�$_�,Ԧ�MA �o�66�ax�{���8�乢r����!���6~�H��6���\c�!�\���Fe.� ���G��Q5�+眿e���~�n���|

���P�C��S��e��3c�<�k���>�K���ʿ�Ւ�,s�?[��43�Y�O~(�&nL�|������Cmf��t�Cm���7k}�T�>=�z���Q|M3�38E)��>G5o�rܐ��ɇ��O�x,��de9e���Aae�X�-��M�k*#�����Y�3���Vo㒫�ǚ*�?�sl�k��"�J�� �J�X�MSrr��G!|K|-�wA�<�c�]P~�O���Յ�{�M���|�oޏ�VL�4T�}ʽs��5��/��8l��.l9�o�-\=��.o���_��)���SV�H�&{tS��q���[&��w���@,F~m|�A�'�F��&���R���S�M:BF���\�W���٭�v�ꕥ�л|����J�k�FR����&6,.aJ];~(�Pͮ{G]�D+'܏|=ұv7��n���Fҳ�c"?!�Ή�����Xw}I��(,��j�%w��$�|��l�O4\΍�!�ғ��RFj
����lQ�ۼ1�`�?7��@1>�A)v�&2?�F�s��o�����`�9OX� �+f/� ��6i�ę��wJ|�.�b�/JYp��� S���󦃶���=�$�ޒ������s��x!_^�:gj��H+cy'�Ec�g�b�w�*���'�j��st{KH����Un���{��T�� �\eG����*B�+L��mo�\m���і$�#�OvEl�x��a���>b�ȁ��4#�='��0���h;�'��_Jx�Vc�Gۢ(E��<n�qq�P�m����F��N�H��̱)�0N�J
k�mO^�:��o��>�G�2� �2,�ac�5�8Պ��g��x�T߽�M��*
�&���+Z�uӗ�T:):=��7̻eA�t����Olt�ρe��~ֿKS��,w4{�`��/�KGH;�<#O����v��t�v��KW��;\�TӹHz3�ְ��0A�
��ðr��@��o([�\�����M��/^��VW	)��Ν�k�H4	�Mʋ��"�������h�Ǫӿ��-kwDB�'b���o�CUA�&7�w0@�L�>x�,����V�P���<�̌���@a�����H�f*I��c(���.�����Y'��t�V�U:�m����n�ɏ���;��*���q�;W&I���|
�!9OQM~\��b�2���x�����oq"u�Xp�HV�e$�g36&��0���T��#L�(ŃU"o�zr;��bC�_��b�ģ��`��Dk����J��H�;��"~� ɢQ,��ܵ�MU�o}Ժ��iWծ�y�69��z��qm=��,���+��1��9\�5�@)ډV���*�)��fx��FE��k��N�ڃ4�Y�v��k����Y�b�����؟�t�N�h���(sւSe���x�o��-V��d�ϰ���=��W[%�^.���ӓ�^p��`�V���`��0H�����~����P֌ +'��Wr
�E��&�8Q�*����q������è@(`Vv�	Yկ{�5�6�<:��B����ҿR�j���o���Y�s���������a�O������И�����Hx�	S���5�/�S�(��᜿����U��`i򲅔�s������s���l!p����!7��[D���b-'��9��6�W �r����..Q�haƈЭ:��)q�;ż��E�G^��
�����󙂴��FL���9�	��qp�\j�_@�N�n��鏜�e��'��z�EpIHĸ�V�aB(��ql\��r~	sZrn��H}'�?Q�@��m��E{]�5��k������e����5����5��MN��������M���;eM�7~���zΕL�=H�l��a+9����U1hV���Wf�����?tT�n�jR;}������xo����֞���F���WYa>��炟p�G���n'z�t-@���>�ZeMÈp'+�Ə�1�>��[8=4��5+7�� ��Z��! ՜.�#śB:���?��c��e�O����ߺ�V��P�R&t�꼬���N<�{�$�0p໏e�B��e[������Oͽ��%�����6.
�&��d"�4R�ũ�a��lK@����)�J�m�Ů�h}��=�Q3���V#\\�]g�v��!�[K�F��������n+zG@�9Dd��I�Y�c0��5���0�I� Rg���S��KV��G����M6�H\�#��@���L�{��xH9'0���s��h_����DߋflG����8xh, �aNGкg���?^D8N�@�1�q����p�޴eݱh�9�r����F�|���l�Թn�;�L���J>ʯ��#��u�+*t�DGx���.c�ۓ��ʫâ"q�d��g�~��N�)p^�WP�)��C�
�!S��x
�W͠&I��df1��>vH��ZNx�3`�3TI�3�m�D!vMp��_Y>1pBOާ3:J�SNo�B�7��zp!�{l=q-�ԟ���ѳ��(x�4�U�9��]N���S	�(�l%ƣԖ�(��ņ
��=�y�EG�a.���>djM�=��҇��(��N�x�2m� �N���N�O%�_�)�۷q(����ob|(������~"����y��+.��2;�E[쇰-�V���Zp����rs�Ew�2��z�?"���ct��O���4�N�BJwh�H"���-��Rï�A.�F�Gl�t5�Y��Ѓ�)Z�����s�U*NYI�����Tug��M{�N;L�^��m�	tzz�1�/ʘ���B$kAQ�ˮ5���2�Up[�s��{��8�P��]�T=_ƹ	Ax���Lq�\��X<x��3�DBZ
�}�y]����`c���ˣ!����m��������+n��ey!Vz�)�U����ȷ^�Df���E�5u؊�£\�p�G�Yb�Ϲ��e���{�����B�/�^��"	����]M^^����0�ZP��8�X���0�.#��a��!�՞����b�ã�1�:7�BS:�,bj?j��W9��:��M ���Re�z^A=��>Ԛv>��B}k��n�����Y���Y4O;�U�tq�J��ŵ	Q<}qQ�X�d�a�2�O��p7�(-eo�~��	Oɛ�s(�D�L�ꏶ�HΞy��8S�m	�{d0����C��V����zS��g�RI���?�~��7��kʐ��J���:i�W1�#)jH.�lh/�Nk^��`Y�Z�����n��Z,$أ#z�f��AkC��w����J��l�k��¿سB�����s�>���ܜ���*5T'�}��ǡ�+׀������Wz���U?G1�W�u�,/�p���p��F���w������Q:��	"���ܫ0f(�oڒ����p��%�0U����6A�-�>j�$ʾ0�xp}�Ƕ΃~�ˡJ�[��ho��=�{v?����'*�� >�I���k��S�c�u��3���s����Ct����K�ݾ��/}���y\Sv���R�g�f6h�sQ�w�9�М�r���2j���i�do���ϛЬS򆁪D�剾�ƅHaĂ��G	��R{1������:N/_ky4�6B���e"ZY�����nE_4`���y�W2QNc�{�a�*m��O�	z琅C��=�!c��^��7��-�I�ļ#�����}��|�Q�����Y^��K��i!|6����]�C�����7�����.�"�Z1����qh�r˽0ԬqS�����d�SO�E��d2�ԏC����+22?1�3�r�ݡ��Ymgܓ�9��<uBaP� 
Z6��w�K�5�!�7��-�o�?��'���y�Wh����o݃�V���(�}�k^���7�/����7��O/n(%��3/@������=$�d
rE�^D4����wS��5S�����2��C$�F(������ =�+T��r\�1Oр0���f��ZW�BGqdSC���d��W���f�xP�]�b�4�A>�+��އ�)�:\�s�+�.�aᖒ��a�`���_Q��:�x���h2�X	���R�R?����W�>��s~~	3�h��P&��V(�8��ش}�	�,��k�Z��}\���Jn��]N�e{}B�s��>*Z=2q��Z�$�O��af�An��o�k�ٗ�q�B��[6Őp�B���AB�:��d+/P���<�va���y���E�O*��we�M)����G)��(��u�C�oi;ʒ�t���d{�ԁ�W�N�/���c�[ş�� <�@���S��(W�;ZKj^�d��y��7�X�"�H�Y�aI�dW�	#.���b���z���0��V=���@�U=����V�UPou{��i��Z/��	�EE!���l�U�������w��O����&Y���ng׌�fp�X�� w�+���J~��x�:s	�Ɠ�"��,�w�~͓!D�ж��kڦ�8j/�Z���t7����v>�c1J�8ߑ7�wUr��i��۞&K��0`n�E\�������t>��`��Ey;��u��-�\o>�	ւP߼wOۯ-պ2�vj;iņ�D#-�3��G��󅵍@
������B����}�?Tyz, ���>�PQ���(��ʊ��h�+5��u��A����C7.5a����&��̎g)��<X���Fީ�������4v�K��ߡ9�����Xd���L<��WlZ���z#I��=�8�����4�;\��$]t��!q��	��$u����gZ��_',a�jNa�M�򣵪#Z5�u �Q����+6�T�����M��)�!����^�]���Ѳ��^��RaZV�H]�5]\�CL����:K�d����ᙜ��9���.*3z���>&^�лnQ_�s�oƋ�i{���.c���M(��^e��^�¥f#�>;D�������>�l2#g��F�*�����I�#~��[�|��2����uj���uھz��y�^�j���>��`'�%4�-@O�^�Ae��5��I�/m��i��+�NZ����a�ie�'$��<Xv)_f�����J>	��W����G��@�����.� �b�n����+1Oj
�d���^6c�ɫ�F>*���w�ېBUq�5��dm5��F0~����]:�~�Y����I�L�U=���כ���A��C�z�i�#:ږ����,�*�:�5�*˻�Lk���%9����V�6 ���k���ϼ��S�Sd=�	�,L�h�N��5�Д��j��cí� ���n�a�a��S���nX�r�FĚ�(M���%����%:bX$-m�m�Y��E��k��8����'�v�$����"Z�|��[������b�fg7�����K��Z���	�_�q�J}`�%8a���yhbOZ��=W�+8x��Om03�|�V��&3���^�r���A��.m)��+L�fQ����~�Ḫ�G�3&È�I��7�i��-p��<�I���L����l]��������QX��u��������GP��qc�|q��q�EPtB����U{�+�)�.���=
g�������yކ˹�=-�݌�T�x{��J��ʇ��t8x٣��|_���h�UA���s������r"�w���{!:��?7���+*3�m���h e�|���w�S����-d���7٥Tvvf���9V*�2"{�y��}�s�!�Ǳ��c�n����������5�㺮���w�������*�xU��p�3&�qMI�M����\�aY��%|������ղ�r'�E"�(��E�t�"A�$����,�zB�G���V1�OB�7��_����p�m� @�����������%;����.�WG�t֬2išL�1A��Z�W-'˨���z����;;к)]T���TbI�����!]���G�LM!vh�!r@�u��WG�o�ě���z�v'l���wA#�|a�Y�������Gew��U�����;1+��<Z�R����x,�1���YO�~��8�%�4���\�c��J\��Xd�X�t��g�����-P�����#��oV6愸n����8܄}���f><9�1���C���Tػp�����R륎�i����7�b�����mm,��~��E��Y�J��B�-�����C_͢�ɤ���+nq�EtV¿��6e�����ld/�f#�J 5��r1�@tlZS^ۖѤ�����E��@�"�O������?�uiq楦KTvH�
�I;��u�tC߂��ju���N�@����+l��^��YӒξ��M�m���cEqԱ�r��3z��o!�5��=��wuu�;�(T��>ȶf����B�ߏw�͚���f 	3mkB����O~-��.�j�kӵ�0��m�'���-�9%��հrİ���pXAhȜD�'J��������F��4it� -ػ��ϛC����W@�h����ͷ�5�%`d��:�Ɋ��%�c�! j�j�k�Um2�j+Ͼ��OJ_d����M���81���Ur�����/}�U�h�!ۗ(A:�@YRՇ��I�%]�ڷ�)J��8S�k@���j�m���ݝ�?��C�����!�otJF�N\T�u��e �N ̛��"�f�c�URV��2�$�_.�MoŖ�eh?��* �}&��L�NBGŃc�>Pv�D��k�&mŌ�����w�#�!+u:s���O��(���7����f�iU�\�6as�8`Z	 z<Ug?N����30�o�tm�&Pw�}!8^Z���d�IZ�;���
�У����S&~�%������v�U���a���$��U�L����Z癌�;)�{���/�?bd��)�p$[���m����l'b����]��=�z��9�OO�G��V�~Z|�O*�t�e��la�j򁬧�wg��Q�;d��2�h:iz>�t����!���Txt[���:�&(�J[Β~6iO>����ì�'py!�7:'��B���w���pN�]���������:;s)�ԙ�-#���h퇙
(6Pf������z�>�@љ��=�j��d�QeX{�ҪWf~���~2��ј%��ܩ�T1�x�E�:��=�p/����)��{q�jR��G�P_*�� �Z 8V=v!��'�ʓ.*����x��j!Ñ�ǽ��8I�{�·H��$�����Z$R[,��Up}�p�|��I��ˉc���v�0Bz�K��{)'{ˁ!O���y�`���c�q���O�G�����h/�����������������%�l��+=4�o���^5��f�<�4çe6:���`!!�u��[�%��n�	�Ǜ�s�U��w����wOӄ)�S�������� �M��.����=$��9�������d�\���1c�W�[Y.ѭ��X����U�x6�AH��M�K���v�,���{���ܜ�������V[Źؿިw9nX�ݮ��r1M�j��s���H� �	ws�T.mz=�,�@��o�~6G>P�0͎!|���A,��9���:��k�M|��=��9Dl���9�7��C#��s�؃a2�5( ,�k+���N�{��[�O�&9E�x�rǨ���B&��%K�����h��aN{�1r�ĭ7��a���_MQf*�"킞�/3症
习�T�Wc���f���	�N��V�����E��V��.7�f4�֏`d-��`��>��S����2Ш����y�|���aݼ���E���G�Z�?���̦�x����bp����u�̳Z�m�՗mBoF�W�P��F>$�7�ҰvmuO{QST�O�1�veZ��:�����P-*��ٸ�3^�o}V��iB]����ǿz��]��&%��	�߸�~1�1����e���U׳i��Q��^,���-f6��� *���/Z:\8�x��</�z�����ﶾV?���5aM8�Pf�g�sQ֯��^�/w
�Z�)���7����K�cۢ����0 8nҞ�}M,o��4]%���,���x5�sBf��q?��}4�L�x��Z&G(�g�sܸn=�߉Af�l�>�!�:6�^�S�P�P��� B��ٗ�"�FC�hV�Kb' FoE8Y�uz�n���an���g�9���������PaBKJ�B"� �EK}����v�����Ҍu2
�9[ g	�U�Qn>-+9vI#���
J7������"ÈIps^��r.L����n?����9���[O��v��������"ڃ[]%���%�C�o��p�"Z�Y̊VT��$��L����ǮzԼ�'��\9k�5�bZ1��7�<:�q�ы1�zخ�-�Wk�c����K%>����Ȫ�Q�^s$ZϊA!*��߽H�L=�GL ���p?�^l�h��}{>׫{N�X�R�Nl��\Q��zf�n���^�@t��\+��9^�Q��ojl�z0y�:��yr��_H�P}����Z (�3�i�e�#�W�hprky3��3��l�dd��]��/�-hg�3��(w��'���u(�>�z�d&zam��9?ɧ�v^3($,JnP�xubB��*�&������!M�w�������������F*NUI/���e�-l�U����c%�Mi{r X���`�y�������} �Ĕ��vw5�[�4;�4� ��x/��o�O%'#/��o"�i���{�n��8`���./�ě[�_2)X���As��TJ�&=j#�⹖ְxc^PL����qW��Y)�̺Ѝ#@�)����{g�2Qdg(|���B��Ҩ��L[�����ߴ�yښ�3pzj��-C6�f��j��(�vx�q��d��%�=��,��\�Gޠ�y��.����g�/r��?���NH:�XV+C��"� c3HSPDv���w�u2��˫�q)1s�5?�S޴�q�KyѬ��ϳK��9��z�e%�x��23���m].�t����s�v�*�>������fh�I�ׅ�{����ؐ�U�3XR���,�|:�u�v+��hD]D%��Kj����k�<u⑂?����Q�.�}~F�?e
;��3֓�����Y��ս���=ai�����as��|Z�)�,Ōpc43�ߣ��Q�:��ht���ftv�^��� }6�~s	��;�����k�s�R��ʁ.�L��j��y<�������*�p5��� �~���U�|\��71.t�0�T���~�A6�Q�-�<>����h��$S�Wߢ/�{���Sª���ЗB�@?Ll�7�
�hP�Ѝ,OĬDE�W�o+��^��('qJ_�T�$�>ȿZZ���r��Cc��Ɩ�w
�y�8�+�Ү��fQ�X������"� B�������0Q�mX"�?~p{iOs��UǠ��=�H��[w�>�aihO�.O���~���y���d<�/K��x�Q3 �F����~%�mG?d��[ ���=�d}�;)J���a�6�_� ^���F���z�_6����k*9��B�s��G��e��y �	���J����=��/p;���cTc q��;r���rLb�ߟ}$��҄���L��C��~3k)�D�ybE����j�D�D�Y|EBxk7�b�|�2�x�) �J��d�at��1��J M84������W�ri`WxF:A�@��X��t���R O
35�D7��{��=�t'ҭKMv
n�imD�7��Y�����f!�W���vR=o�y0�Ͽ#�j9/�#�ȏ�r|>�+��N4�U	C�9SR^|��jG�Ī[�yu�{ =��sm�U��Hگ�6F��B�	ɛ�O#2"��;����Uo�G���b�=�G��8-�l0(啂7/3���7��䄀e�k8�N���Tŧa<1�<�f�}+?�cq,C�I�dF�n��;D���ѹ�х�g��ĥ�'������cz�3�s�Q�wˬ��]*J�wcoo��`1�wJ��py���Y�1��-i���dߺ��l�`R�AS��Պu
T���)tl^|�n��}>v%��k/�L"1n:a��g!~ݻ�4�pw���}�Us|}U8���Y^�r8��&FmG�ҧ�1V�l���C>ccFG�Ko��D���s��H�s�J_�>^U�Sf?�s�u�+zD^�4�z�~?��)oҘ٭]y��Ĥ�G�x+�nmϭBW̴�̀�^Q��@{���^D~|W��#Z����w������w���ԉ�@�ΰ�y��+��u���o��H@�5��^�6ܠd;��@�c���j���[�T�$��g�D�|$Φ}�j��:��j:��)|��/�ڟ�I�5C�uϼ�z��� ���
�6���(P���!�� Կ�f���a�m���U�����g�D1��-��S�B�lV�Ys�;����W��g��p�7���e��Q!J���A�X|��%rT�@[C=da��[�Iy�H���MM��?����.q�uF[ȫ5A�Ю�J���%��S����Y4���@��Y}�G]�J�����`%�-KDzS����O=��*�����A�É�p�維S��$���ə����T�mx�IE�rV�+f�#�G���-����5�;T��U�E=ДH
T/�uA�(k������g��݆7+����ߜE���TCb�5���W�r<��<.�����Z��!�2У��eh��A�J�I��@�[n��^0���z'w/�O�U�d}�­�|��:?�It��INR�w���K��[=����F�آށ�?�/�[�W���;[gx{�#��E�y���&A����淟�`^YM�W�Os��A����ZЮ^���1�mow�jǬn��eЮ)����J�����c*��C`DJ�G�'��
�������Ѵ�!�H'�Oӽ�@���%9�T�]��p.�u��M��&4��s;��6�l&�+Z�3��V/?9]�pC#�)���Z�Va���W��*C���E�ػY���B���"��/p�<?����i������p���������%��a������j�����}K�[����A� ^ z��t0h���S��ӆ���(��{ ͹���W��l�HY��D�Lg�6�LvP[���ډ�7*�h�����6��V/�a�l���%�����l��~a��p��1�<"mјd�}ثкD���Q���?	3��1�Ô��;:�>|ȶ��jVV�Z&���͓2[��G�1���
�{�A$9�q���-��{7��<�M8����9��*|�Hx����j���~�I�F��:'��;0����db�o{�H������ދ��/�;�����C#k�$�Ec��Wh��J�
*�����]~3_��I�U�i�y�
�c�q�K�W�c�4���oN���M���;Yu��>��*a]���l���gt����Yc��O%3��4,j������e��V�}~<+�%]�e<Z'���u�L�tPz�m�������Q��l���ן��3[]ΈV���
6O�_�'Ö��#	s <�s�~����|��H�O�
8�Vq�o
���7x�z�����@��8�$����}�;I�N�qܚ^�����F"S=0�^;싢��;��q(��$:�	#� ����|����*�� �Qf�=�!���i�h�0 �����l�[�m�Ut�4@�@�0ua���.��W"�w�����O�f.�u�t_/o�u����L�9ݗ�s��Քl>a���G�MQ��
�a�Eg�#��?xI�֊&�U^��FM�o��bC`#i������M�s=�L_l��+�N��8tc��T��xl�n���������G��&_����6���cx0r��%Ӄ�$ʤ�ӸL�$�0��ߖĞc�f�.ߥ����5A2"k�Bp\? ӷB���f����B2=4E<w���"�����<����X�������_��^?����kVD������qn|��ɟ)v���0���LP�oZ����<c�!]�rG�1��q�%P���ף ����KO/ׇ��+�M���Wc�M���� 1:�EY��ǏCb��/������V��GU�.
#l�	/=�8 ���,�Ch�*��j2�j|߭���G �w��I���̗/S���o��_�A�ub���mq�E.M� �VK˰�8>?&��T�	G�+��R����?�	�-��+���{�
�Ko��~��I͒	&L �q��=���I}Cg�e�:yN����r�e�r ��V���˚�J*�P'�Ƌ8*"�ߚ���;�so�D�iG����Ja��9
�.���O�� 6�Ť�*��TPٹE��m�.�7����Qqϝ��WH���> 0 G�Z\��{���Z� ���u�hQ��,6��ߠ��\����#��c(a4�uP���D?>��5�Y+ˊ�|��أ��s�>ݮ� ?��8����k^i3�߆�r�g� �����$�N
��_�5.*�z����ԣ�3�?����J7���M������WO�v�p:��0�`^ȫ�K�W�e5�ؕ��g,w|��]<�@�S���*��ߕ����E��0T��o�xj(�ƹI}�C�IN�Zʅ�d�x�O����&ϵ��5����P����ϰ��ӂ�+</�_��U�]���975wE�/�"�(P��PGr���e����՝G�x�ҫ�(q|lL�V�$��ߓ^��hT�q	��,�K��y�^PP�6����o�\3��{�pNg'�!-F�ܭ�Ne�^�fP��eV�QׄͰ�.�肤��ߵ�U5�<���Wg�0bY�U��3O�� ���sGa3�-Ӥ����1�Lot�_�������e�9��M�2+����>}�c*AX4�yJL�A��, W?<+Ȅ@3'S�͡�%n��>L4��Q���������#�E���Y?_I� �����|�!#�0��J:K蟫E0�&���4oZ�4V�ܬ��/�O�� ��i��q*�>m��֤դg�
�0��&��h�~wo���~�x66x�K�-���@<���ݺg��V�*�iq����A��Q�jѾ�p��n�գ�F�#�/�N	���F���O�g~|(>>�� E��0/��������o65��n�#�����=�h�P�V�����T{�굜������Ud�*w��k��::��A��?��p���,rwB%�5���g+��'�ЀaR�R���j��!�yt~���?�����k��pC�QZ��,}R�"��}�g��F�a	�����
S(]A�Ә-��t'�k1,��B	��C��1�\1�[��������I��/��:�=y	j&f��� �@2���8����}h;[�l�hO��7���צZEo�6�u#[�$%j�|�+��?NY�Y@���t�fȗ�A�o��:B�Kپ�b��|�1&ޯ�*�� 0޾yV��3��&C�$�����C@"��6�1j-Ȼ�<�:;�i�ֹe~�}��.~��*�QP
��Zp�\HX�AIykp�4�0kk;�˩����7ˋċ��I��p��-J�`��
�\�P1$D�8�j���X��J��,ʠ�w��;��?$\���Ӣ+r����C(��]��g�)��J�vҸAN��?I�,4%5�q���?|�)�{B��1>OC'��ss���<��\`!::)�+&վ��/�L��O����ؕG�g$0=�*H6��H`]JЎwC�%ޣ�δ��]ߞ�	����ϊ�ɘ@��^�<�z_wj��<�Ԅ��m�@.x�}Syz�>�U�t�3*�a�)��)i�w}-sPkc"��;Hx����P}�k��	j���+hfE]�X�+�X�����\𣯿Y�K8����]-���[�F�ËAܐs��1o���x"�����B�٠�3�mfƮ��lymZ��9]�s��]���g�B��&��D��U}1���l�GnF�j�����q���ҹS�~M��H���K���Zt�;vmL����	i�n��w�Ɯ��<Sˬ~w�9�;�_4�y<��m_3�!�}2K+������/U�x����/\n<[@{��@�:���`�'����MKv���z
�6�(����� ��q]a�7�DZ���苼��6���ږ����q���`�RW�f���}*S�k��*9G�'e7�:Q���3��w/���غ��:O�Á�G�:q<C��,z�grx> ZV�Ҏ�^�������,D�����)HJ-��U��*�2��8~�>������[��?9����R���o-�-�#w����7{��3�d���Fwږ7(G�ék�Fɧ-L�?p�������(��h�?�Ӟ)-�	n�RD��c�p>H!:��]�M�ܙ���l6�b]�i��zj�?3;e�X'٭�m|N�����-���;��eF���$�~�k��2��U�'�2�)'@��6R@;+O�o"�{'�6�Р֥U%��^O�z��9���{�:=�x��|c���)�m�Iݘ�M�0�����禘�m���}��C���;]��ˁޙ��Qw����Ϧ�P�7�l����8������S!���ｒ�v���<.rťn��ߪ�����s�$���\��ΉY"�[��~X���:	Z���l`�Q�.����o#�g��2�4��=,�*��7����q���v��r�Ga�:4��-c�������Fl����z���ֺZ~|)(���7"�����5Ҩ7����`׈���͎V'��쁆T
'[3x�� $�)Dn|�%޸���� |��B��BHy6���m�)cPV���@u�{γ�ѕ����6�F�h=�qP_Ugf:rV8�l����;kE�s'����g[�=��ux��O��be��l>+
��3}:<��?]��R6(���ڒ�k�W�����x=I�%����#KL+K
��@�V�|�
2= �_eCsR��ߠ��\�6��-_I�#7͏y�ǌ�����dɬHNp��2c�h��Z��V�сxM��?%t��0u���	�d)�Eg�5� �h��v6qB0ݛ����{���!�g#��M����􅾟�vZF�g�����ax�������� ����/��,xX�
��sz�&&9�3�C�bU\q'�_m��?Y���[�+���A*5�3v�u�̍ᛤ�?!rG��~��6������;�ia-n��?�V�KV(��n�ƙ���T5����r
��/_����
k�Q��<�o���K��F�T�r@�}��r�F�7�k|����{S�2�-��
L��d��]���M$.��+4�2��c8]��z�S�x�L�s �;���Ǔ��'ofT p�
n?�/E�M�V����ur�w�j������I��v�r�9FF�}�.�d�]��\��CX߄��:����FC��{SF�e��G���*�]'��w���^҇��.^^�X/{�vi`��"��?��#m~q���F9`j��O�������T��&�r��a	q����C�aT��"���41�h
L�ΰ�n�L�	A����aۭ��mz��)���y�k76<�LZX�v���wق�ᩬ&��`��nN����ލֲ�<�u��]�jg��~X�d����؝N���+���9��4F��7���{��@@� �μa���y�&S�s��M�m�]=��o6:��{��#Lb��
�1\�7�I'V��ޡS(=��/y����G]�\C�3֝��s���c$zܸ�7XXR�x�����w��I�c9�-/����;��|����,�6^e��HOX�Ε�b4�ί����;ۣm����K� J�����tf��	*A��˔�;���<��O_Z9:ة��{�X�d�G�F�*}��-�s5�VX)��	�(0;��GE�e~ym4�t��q���R��:�����.M��7�ʰ����'��B�d���%{��*�����/���·����LJ��"�͔��fc�c��)\ZP�)i?t����{�yN�#�i0��U��=��;V�w�՚P��+��w� ���A��r�z�r��(0��Q��[�j߿�/���O،�X,o�=���"9x���zo�]m���1O���
b����*+���f���`���	#ӗ�\c�.����T�rT|�oG�%P�����`j�{�I�E��o΢`�Ƹ��(���Rwć~�~��, ���2^���D�����	������կ��b�A�J��]5f�R��|8]�r�u�d��q)~ѕ[�Z�^��Ь<j���c¦L+LiH��v+�)(����Zq�Oٕ�Q�t�,,� ��|`��]����pWH�7�= ��2/ݒ��yK��(�2K#jJ�' ��m+�{���|p�Ǯ~��MSο�/YȂ�g|\$�~ڞ��14a9���v�^F����ws��=��S�v�s��%g���ߪ�|�2׀����	���ː5������՝�W������&��%�u�o{�4)@��?xKRD��E�vHЅ˗��4O[�����^�o{3��sޖ�F)���Y��4wge(�����Q�Y���nkh��y�u�ja���kL��0UR�7�l�6�I���.b�&�KI��t&~�M�D9,���#�CP;`"��8��WVbhHգ�뉋�y����ȚZ�p����3�l0���۫Ύw6.����ѷ�
��N�#ɂ�JV��%���$~1���z�t����ȳb�{ۂ�SNS����qJt.�
�Aor_�3���g[%dJ�%Q�f}��~���l�r���K� 0.,�5���2}�eGk]EV@y��U�`��C_����o���ෂ��{��g���bDYmZ��§�~̶��s5P��ô�V��O�&5�J���q��H�
�%�"�����Q��(�h(��FW�*0��"���/ȝ�,�=8Y�������sr.��M��7H�Զg4��y�Q��H�Bmj�u=P怳��߁��%�&70Aȉ/�6��_�E?�	���T��y��e�[K�F궏NT�o�FRS�����ɖ�2�����/M��0��K�1ڃ��q����r; *�;p��GN��S���E_f���!2d���t�1�k��甮M���Y��B����o�u;B>W�O�]�wu�4�9��pXo%��>��`�?Y&!G��IZ��۟�ߐI/2/[ul�U� Ќ�,�Z
X��V��>&�9���̳*R���f][%KX���պ��*��e�Dr�Ar�'b{)}�J���x�d?���>���ޱ���;����tZ;q+%�?�D�gS��K�!ٓ<j+G��Nr-���m��T3~�0��� .�W���s[�]f4����r"����Ge	j��-}��A�7�#�)%�����ퟵƓS!Bp.7Uڅ��W��v���y�E�V_�➃���l�ߐvS��
 �>.��.�8{�^"#�4�3x�����Yk?ѯWMB-�=��L�8�	�ƒ�C�B��N������3NQ��G@^��jq4ǃ�ŎG��;�;�dMvh/^�̻qy�]��Q٦W�<8�+5ƕ'՚�1y:!�����������<�<=��a�Ÿ[�6�͎�ԦȸR���7����J@�qZ�1�A����,��.�ьP�]I����9��%_�[���Ž��>x����E��c%��M���2��R�viRw.�pR���GU����<C�szP����[bĤE0��&��k�4���J�=�	ո6�q��ntz�{Q�1��v|��a�ܗ��v�Ӿ�fP�B6Ed\n�k���*��as8bk㖋����鉟�$�?Z.莒�Yͻ���g���_y�<��r)�^� �\d����c�עV�G0E+�_ȥ�Au��~0
���a�f�B�k���&�{m&����Q�eV�e`�9��6��M?6�8�{ЀV�H`�\���c�K�ʣ�6:�@��^=a٣�
�x�L�"�E���0�̎�oyə���h�.<���뜓���U�~{����zۑ��a\��E�S�Ʈ���j�گ�-��rT�1�)� Φ�>�+����;ž����xJ>ze��	bM��Rn{�W�Ao�����r/%� ���A�P�HgL�8&��ˇ���m�ʽb��("����"�Y����X�8��������MFMF���Q��G���-��1�&�N�L��Pw��b��z�瀡WP�'��:/󜭭u��H��|C���1�˪��
&F����?��?�9g�7�~���6�����z����LQA/6dv_o�u�D_c��5�x��"��O�*OV�A����[��RI����Er������K�2�ޛ�?��\���Fi��`>����L��]e9G��������c/����2w�ɡ���>=�T fz�[�}�u�k,?i�U�������7窓2�9��csY���s�ע[R4}���@�%��4:g'F���i�J�NEh�S�_�U��J�!ܨ�O�	�^�]�͔��.S���#!���]@�PʙDn4ҫ��2w���/h�l��{��o�lTOg��Z���T�Z��ZG �K�ߔ�}]��w�d�'�U�P<a4�ݻ,t�|�E��4����7��6@��'�*6?�̟h�Z�'X����BM:ߵOz����������SS�����ӊ��I>�Y>�eM|��M�b����`��C*s���h
�	�Q����/,((njljD�o,��>+^� L�lZ�1�y��K��ߊE��ފ�SK�p�>�<b|�.�NF��pm���AG��FU��ڛ��A�9V�bO͉�1��۶~�ۙz
�-ݙj
$���|�e�IX��B��G���>�%Y~�j8�P�J�}�Ͱ��a��h/h@p��£��e�`��W5n���ݰ���]e�5��7�B�m/%���Nx���
�`�k��g��g�
�dl�:�R���a��\mՌ�{Ŷ��Ã����z�X��S!*T��"拉>q"����bkIYB�FzTM�9�@"y�HUO�g��>�w_%�w����L�/Y��>��-���B�-���K����i(���]���qͱ�d�]k�j�����D�3Õ-S��֡�=n�u�<I�A�w�M��O�i��z�ק��{xz�XR\i�&��f��K�q�b�v�W9_�"��GOG�r�.5�slAҠ���/y߱��������2ǘ�Q���􅲦&
U=�)�ޞ��za �Z�2����w/'C��/��<׋V�̣g >�j�~B���3C�"F"��8N���81v�]'��b�E��P�B=s]��StTe Lh�Ȑ�~�D~�Xŋv��^G��,����S?�������ov�~>+��x=ۦ'��6�f���qK#s0��wC�����m��x&I���f�@9�q�:��K|���t�)��φ�����v�$���ˈ� N_�v�/��`e���87��_�IK4�<[��N��ȓ�&$j9/�zU:]e��}�,��qR���cr*[X��d�
)�/�^�e���}	�nt	�;ʊ���h�DV֌�Zſ���|wG�]Lp�7���r9�֏�G��X�1�!Q)B��bQ��˞�8�ێ�F��`�~���P�?l?�st���nU�����<K�p�x��[+�v�r��iʀ���^��F��
�ͱ�x�O�[�3'��?b�ص�}������Rs��s��raM�Y�(��<��:��֊}���Ux�u���{ vݡ4,VI����fQE�<)L{��|��4�/&��K�������{��r��u��}���P��Pu�9�Rd`�3Z49T<���p�ޒ
L����;����C�a��\���l��+��kK�W�2Ό�lYd^�
��l���fS������ �(�����燏
�՛A���ʖ�J�S�������4a�k�����o�Brx.]8*Y�Շ�B�����I�պ�;���*����-��5P�K/,̚R-�Z�`	��[���P^k��o�����-�oj�z�!�d�đ��sG���p�|o��VG�Dϛx�#B�l9)�AH�tC/��J*&]����S��ns��=�����DD_�C�n`u �ҥ��ߌ�f�t�jJf [���b)�� ������Z��Qщ��D�Q��҈��S�G h�����H�x��ϭc��N�	�ht���Ⱦ6�^>φQ[`���¨�V��X˱|�j���D�JD�D�&T�wI�^�4;2Kx{
��C6��eVqoz��g�+I�= �E�q���ܴ�x��2ň�M���X����+���##��@����V��Ջa5��D���W��8��$g`��ox�����|z�|���4}�﷌��F��#��߶#>�J#6!Xq/��`�p%j�0�]a�����k�цix�+�x��uĊ�����Z�R���H"�A��F�a$������GOSd�ai��R�@�u]I�0V�c�-m�Z'S�� 0��r���;���~5���X0T���L�����E��b�z ,��tH�b�z��2r��`��X���L�;�W����»�9}���HSL�bi��z��U�yɃ-C[/7������t6��N݋�s�h�ƻ�;n�B��𑡖̻�g8H����
��T1Ế[�{��iD�i���rF��?���tg��Z�7�	G����Pi1lH]u}_>�} ؊��
��ٜ���nRg��ˬ�JgH����+���E�DJS�t��3�
��?B��7k�ҝ�:~���ˀ��M�$t��+4h��bp�����(�F�U�?9� �j��c��5�,����L�h>c&3�Ջt�>[ዝ����,Id�Q��#�м�[�?R��1UWMt���1�҄L�Zl�-��ë�Ơ��.�6�#D*pDlK�/t�:R�~��ԴIߋfs�����d�:�_��3�M,Ү(��rK*���2�9$|Ċ;���))����`���<��������j��3�D�8���猅
��`��<J'�3A�ڕ��|'��KH��Q�����_�;�>����6h%�4zO�7���|W9BH��7Q�*<�e�/���J-x���� vJdZ4Q��N��^��ܞc]$��5�{r��L8�H함��V�W���]�v��]���>g&�}��<`c���<�F<��r�;����nt��E�����	ŊW$��t��.ɗ�A:��D`[����=��j��̕WT�aI�������8a�Ԝ�F�#�����z�K�G�d�ʭS7u�|����)`�erc�I��cE@��E�YI�l�NB�1&�|y�굅��T-E@@�Y/w����o�Z'�����!gJ������-F�_���Ӈ?m��C��Y���Ϗ߮r+�ͩK�Q#KL4"��hL_�X�4":~!�H�#,*/vz���z�N�~�[ar��c(s��rz�I�t)�<�5^��l]�>�]e�ⷪK���������luI��2����6���Z5����#=�Ґ�F��~ 9:���ñH��{*�/�ʝ�/n�}oVw�B�s�9���[���_�����!p�6���V�*f���w���jG����/t&̜� �v��sԤ
V��4�
������Nz�,�<�ey˞Ѥ��������}��9E��I����ѻZg��^�J-2z��]&,8�tkt��@k��z��u;��` <B���!y���<�;-�k|;L���`38��-g5~Ղfi�:�7<l�De~������]7%�soѭ�4�"����ņ�G2<��&a:��f,z�9�U��L�NF~T�M��"���H��b���r�	4������>�A����q��~�D��Wb�VTA�_�)�G��?oz�c���m�K����l���,1�����vVK�4�-���+Xq������}X/M�t��`:뜐V@�"��]!'�Zd�'j�	]�I��l���6LA�.���_	�M��2��������[��c���}C#�A����{�xo��8q$�#�"��)b��I$��.GN��'{4�T�1P�K�����7~\%&�c՝���,O��*�o
N�0vyzKg��<#��={�/w� ��7��0%��C�s�4��p������U�q�H���X����䷜6_<<�B�{M��=��!)�u�V���Բ��`c�
QqKV�ͻE�%`z����M�w"��x���R�!���' �.2��{Tc���UJF?��Doo�<�5X���ګ�L���@�]���D��v}�⬰����]�b�;_L�4�Ţ	����}��ŊC�u���ʶ�/����T@�����-��G&��U�wA�_ΰ�yK��`9���\?�������W���U���
� 6�s��?b���D5�ϔ�%��]��;���^̏�^mmm�7��U�i|!�Q���Df��G�/d�xN�y�y��|[��)�Q�q^�8�4��n�	ouq�;!Go�s�ܰ�3!�-,�ҮTl� ;0e,�yN��v9W�
 ค�g��^�I��zs���QGĹ���rM�%ڨ(�%t�EMS�	-�����8u![^&��
�p �� ���[��CP^�k�?	�厩��[�:�<i�L�v6��u����âj��)i��A�$R�X:$�ai��K@��%v�FJ$�Z��C�=������u��g��3��������pk..�|S�?j��✑��R�������1?�H����Ҫ"���i��=��m�ݥ�te#�<�5ԥ0"��E,�z�����y (@%���M�@Q1m�ʕ
b�MxC�Ϗ7��O��iR{��W�)a��E��&�.u��ct,������B;���(v�$�t�������Y��0hj����&@q�����`G�1'�-ޗ�3���_-q�SP8��^MP�V�jF��Wy�p-14%�m�*v�3�!
z	���>zy�?���n��I�.��)]��5��oƻô��?ϫL����^����u	��#h��G:��"��qgC�00� �<}�}��$]a�4�z��j}�>b<(q�	�]=�5�@�SI���7��[ ��4rL�`uiJ�AQ�6�9��y����w�A�b��4I�a�W�f��S�
x��8S���ml��:�{�\�t~~E@�:���wQ~���7'E_���G��.����Ԇ��(��.qϚ*����ߛ���A:�<�l���%%�[M��G�������)�uv,y*�G�ykz��l)��;/
�Zh�9�t��-� �ŎR�z�&=є��Z|&���8�9/O��f�ݾ��7x�gK�x��K-�3P�L����~��Q�xm�Y�a
z*�������^�-�d��k/{�ΔoZNۿқ�dS�j��L�.AN��wn�BxƂ�P/�V=�dw�F<0<u>���=��}J9c��n��HR�?�z�	�w��B�fVMU���	P.�1X�i�V�x�	��r Y����F��W��i�pv����,a�]^r}z��l��=J+����\%�Acl �)��#Q�y��mՃ����w�m�)1P�2E4�%�׮G�thz��S��h���m����L��6���m��K���P����n�kkh��^����̓����(���AÜ}�|��j�14Z��@P�g۾jb;;����l<�g�Yx���8�;�H���ISo�#����׏48C�-�Էozġ]���xU]0
���,S�9D��a�h,E�;$x^����Mߓ�v-�܊�Li��QT$Bssh�gfz��rۜ�Iu����nޏ�����}��@ �d�`-%��u������Y���'@�|a��O�8��Jv����|"}���������g�v���&SS�A�%Mbx������y����:*9L��nt S�	fF�bv`�X���E��U'G�����UN�V ��2.��r�#׮4`ʊ��(8�|t��j�Ox��e��<�v`P��2Q��UP�up�YB�*�Eڥ.c�Y�õ*����j��G�����U��S�����v(��o���*z�+�B��a���- i�����'��<ދ������YI� �^�o��/�dU߶[�T�m�wx	��GM����.Y�t՘��>3ğ+�/8���g��]猰N�]r#�v�7O��>��h��f�<�7�	�e��?��sBU̥_��ݕ�ǎ�Z�v�A�&IH�6���)�|�R���j�20i^޺�1A�e�L-�KC��f�ҟ~�]������7��?���nnKt�`�kh��'�B���/-�2;�,� p���N��=�O٨�c���G���( ���&�2�*��D���1 �
������<b�}{��eA�cUu��>��Ҧ�+S��Z׶Κ����=�*秪=^\�7��
;#��o%lIڨ�7~^����o.[ki��,�:14�����~��}��Jc�����'{t�N5`� x
@�(4��@V�̐	��\gG�ʬbb�3��$�P~C�o/�]��aU{�U�
t�^��aKV�9�[�� ���J�3�h�Y8�{C�yE�V^�n�x�-!0��A���;Ģ������k���<��zi��a���R �Y��k� �g�b�B�2�UY@��k���(Ǘ\W�3�{�k������.��	j��o�򿼠����G���]	d�K#��@�E|fg�O�o�~� �@��E.� %80Z��X�׈g8��\������06��?���S��zy�NsX�1��A�w�l�d/�ju��[�9�C�'�p��[-:y�L�z�C,Z.[����׌�lF���e��sߟ}<<�	�oW��q:�E�M#E,H��|�[3�5�?��%7�"h��o���7Ik�pN��4I4���_�Uś�8���>����^���x_��Xx�(9�0?�������ݡ��?u�lM�t�3N͕�|m G>9��	��r�bå�bn��*�6|�a�`5���:���I����N3L`t<�+�:�^�R�h9�Z궴�x,�, \jdܻť�����'��G �{��5G]%X�$k ~�K�+���&쟬���t����C��Lў��<x��v�QG�H����2�S�r`�+T�����Ѥ�<�Z�<��#�i�^�@��݆�m��V���d�.w��u�Q	�O	�H�v�Fb��UB�g��ʋ����]�Z�.�����~�o��J��4���������%��3CTT#�mM_�
]��Ǵ��u~y\��>���Kdz���i��O̃s�Q� ��j�O"��{�1����=
�1��خ1�.���5]oG%.��A�3�Z�a���6�(d�D,�ߊ��oL����i]��`��%M��&Hـ�@+"�[V���6�̃����SQ�Y�����`�4�ʴ�`�ɠ�*^�KrV�'|�U����'�q���챒V�W伋ײkLh���Q���J�����s\�锗�t<�m�'��������A��=���ڃ��Ϲ�zK����'C�[Y��3u܀03��}�GA�����8y�� �7T���P�Tٝ��8�zEY�︋kM
h���N�O:���h�����b1ɴ�ӻ�Ӫ�?n\C�/9	O��xr��`&-���;����d��΋�/�j$��YJg{7N��V��]�١V�y�dWo�3C�<p����;�c0� p��*$�����r��fZ�_'3Y��+3>s<yw1$�bpn���]�H��ė��l��1�0��69ar[�j}��
c8R-8]a�1���e�{#k�>:���j�V��,��sPhZ����Z��O��e��Ń�#o`�e:UɠH��6����\,�='T�����O�w���o�FZ ڏ����g�y
n?+Ѥ��k�=�*vx��(2��ͤ[�j�����~.~��^�J�����d��U;���Ũ���ҁ���ӌ��d�����vG�̭Ip��L������jW�1(sW�����'���N.��=�T��Ϩ|'>�!���0�Q騒վ �p�;ǆ@Di����҃~��@C%W�l@�N�
y
�t�} #N�i���9=�]�!-��1 ���A��0�ݩ��%������%��/��z�t�udh��I��Zī����F=�m&��|��9������%�O%&;*W�bg��&Ei�/꩕��I��XZ-���Th�fU\���}��)����Ħcc8�"eE(��扉��ʟؽ/�:��)�#�,��RFz�vK�.�lv��a�R4}.�K^D&)�ָu�ķ��|(3S�����@H-����z�"H�c�FS�>,&$�gG���/����L�;L���Wd��"�PV�v�{v�gI��3��#Nw�p���R]� `
��] �2���"��
�������Z�21w�������cM��;��gǃ_"�zۋ���W�h�� J�����]��&���<;l�Fp�Vyre����-'�:U@Swư�4���~�`��W�EX$��HKt���ڒ*v�,>����.�	�'�Bc�2���mF��)���X2���((��	F���ߴ�P�/,۴Z���C$��ڙ�^;5��p�*$r�Ţ"�پ��@u�������T�{Q�2Zo]H�~Ê<�_�>4��qA�Fo"}�g�nt�#Y� ���� B�p�ݩ��`,Ɖc���0�?����1�f�]y�����<����b��`�>���n�쏁��j�(�B/c�3}p4B�E�ԯ*x��;�ܮ޿q�r�R�ݷ�U��u]P��`䄒G(H��������9�:����.	hΝ���"�;��5r���o�y����4���[��3 �a�"���3#�c�LD���Y�PaI�k��z3�V�
�s��C��l�p�h��?�{���~�P�����^��m�����H����VU���s��7G��c�::d"�Yb���d.}V��܀���QԳ���J�'Q�Z��V$x)U��.��-C��7�R�����w�F��ǖQ�hO�S��⣙��n��;U�yrk���u����W���0�*W҆�`�KA�� ��*[SY�f'��t��P��сδ���w�##j@gƢ��v�UH�r��]��_+�;�Q������}A�r1о����gh���4��IJ��7WU�ȟU�8v�]z��q��!VO�+S�>���π�E�1��M4��@���]���K?����H�ŧO������������ݎ{(\�����������T'Ĩ��=��1��<�t��9h,{�-���+'�%�'��%�����*�z/Y���X/�Z����A�� 4���H$�ն�֫��'�=�4�/1�#?��᪯���}��'i//??3�?����wo�Y���p���=p��jK�a~ �~��Ra��C���R}�k�D\��r���(-4��}�/3V�;M���&�%�3 ���!�8��E^U�Utz����(6Y�c#�Nf)Ό�%�<jG�nr)�{�7����<�6�H����K�� �0R��$qkg'ɣ
43gFϗ��"����L��L|���c��MD�;���x�ԕ�e-��Jw�T:����쮵�D"�G�7n�IRqݞ�I#.�"���k�T�|��F,T�%$�#�}�R������,-}�{ҏ���<���d��b�

gz�qo+�+�|�E�'/����`m
�	j]�Gj@n*�-���7�~i��eWQ1^�i��TUÂ��&���f�����%�1?b�R�\��AT�w�sE�εD����# `Nz;����n�?���hy��Ԉ�G(��%4 �gk��Y^�nX���
 Tfx �F��}��}��P���X��L�{O���vS$t~�:��z�<v�E�#����#��9�(N�L^���K�\� E�Ʉ��)��7З8�%05��M������.�΋���8xˁ���[���=g�vA'�v�\"���_r�]�2al��-2p=Wc����<�H��a�}B�k��}cp#�DT��a�8���x����E�\��[C\Ū|}[�rxl�����}$3�����2���0�^E
�Sطda~���l�ҙ"_�� ˜�8�F	��v�ԇ�����x|<p���2����T�x�[Yn)T�%���ϒ��F�Yf,� �m;�ܗ(���$���������CNV�t<KxtL[��Aq��0���lK��sE�9���yE�fՊ[y#���W�A�qe/kf\���������2)7hz��!��^(�Afao���b!���B��gmm���=��t� k��� n���0s_\k��u����D:>���_�x*�.3�X,�P�ZZ�����5�|ԔPS�/Q�5����(���2Zw�2�4��ի�j~B(s���Rx������"��`D��K*epy��J��ߟE]�\.�Ⱦqs:ʶ��zUP���&�Aj�L'�kۯ4��:]�u���0�Ze$��ML
W	mh��b!�n���Pze�M��D�kv��,�w}n�o��^Z�<!'�XǬoH2 A]��1~U��Fˬ	C��#"�H�C^;��
X��a˜t�>��� ,B��:>)�D���V�$O�Y~���ieA�eL�*�^�p����n�X�֟��y��{9^B*���P�&B^&`�u[F؇�(�O�yrY�~�A�PT�粁�3��"$a�-Wi�N�hE���3�V�%��D�K�yЈ�q�'(���[�[O�X�����9&�鿙�z�~�-Z�5k�y��� t8l!��q?��^��aj��A��K�ﻢ��W�#j�x!D�x'�0���}��$>�L�� D�i�P��1��!Q|�`�Qu˞�0�1�‐��Ȑ�����g�}�~�T��Or�l�.���t�1��t��>:s�"a�vZ�������a_�'��J�/�K��6���c���q��:��AJǊ����?�V��wuu�fd$�by ����`���ot�Ԏ�5����[d�:4�����\����	+r�lMĨ��c
�1���-�5^�g��ݞ�bg����'XŤ���5KW�)�m8{��w���9����J�q7� �e�v�)��֬��O���d�@\��,��
��"��H�����?�\�oB� ��A
�X����I��K{X�I ��D	)Y�L�`gTFq����X٬���]�܅�����o2�	������w���駳��l8�mw�>GA
`pÞ��A��h
C٩m�F��vDS��A���~��l8�{��<-�}�t���KJQ��P��~�B�+���� �a!�?�(���~�eOS(�ẽ� ��~�)NU�K0��x+(���TN�l�hYw�	�:`�6\��v�leԾKM*���X�ފ��P�v�9lchX��Ap����Ռ���B�!!�g;h\�n��F�ޮw�?  n�ÅJ����o ml��QW��2�_tT����,d�*LD��*��������k�HG�q�J�y���b��J��7��G���Ơ�tQ� �5L�Ы��d#��G�;�Ao�����[�r_���t�=�n]YU+5��?��Q�<`~���O��� sQŝGe��b����#��O#�tu��z����n�s?�~Fi�=�.��Fm,_�-܆zĒ�5fr����2�i�q�y���
�k}�Tb���(b��W�=���͟�\n@(Zy��*B�n�A�2��m䑩���s	����⃯���/�}���S�����vD��=��ف��|�ұ@���!o�f����m7��ۓA����]�R���+��!DH����c22b�2M�qu���]X�[��վq`�U;�q���1�Ne8p4� ã�m��
��RTxE����ZJvprA�L��A7���뭀���y�qTj�{M��V�k���w��f���|�Úh�S:��
�>l���	�YG�V�2c��򁁦p�8˿8��6�r++����?69?S�ﱿ�n���|D��p(�e�Qd�jW�
/d����|�{8���|T����&�D'����?JW��S�d����A�d�F�f��~c��2h�&��� ���ns��\�$RekKV�CD��O���	7LD
��Þû�C'��i���q��f3�]&L�>�s�_�܀%���m��oZ'����l2�~50<4��ˤ��u�QS��Iw�ە;l���Z�t�������L{����y��;[�"3��N|��O�Ub��Lt�V[���,5-�U<���ۼ�`�Ҫ͞�����׃+W>��j���3��c) �� m]#"�nϊ�����{��ܳ��e ��7�K����59�O�U��\�|��J��>ƀml�����2n���(�Ѓ	�pN9ji�����3�ﶻ��,z��	����������{��8�����4]p���;)V�m�������ZU�4�/ɏ==\,�6���e�d���L�j�������B4���n�2D�sm�����	���Jo_�������ɪ�6�E��%4<BB����<,W:������rӱ��Υ,�o�ݝ�e�D�q����B
�����Z��n����c�P�77�R㵯���&A�Բ���=~�a-ϱY�!P����c��Ќ���������.��l_I)�	�0�y�N������qԜ�c�=�Y{������-?�i%F ����#q�b���W1&Kn��=&7���h؀_ҋE!w�T-������u�(�kY\\���7W��Jg3u������r�s��@��x쨦ɇ7��9,�v�� o.���j�%Y��묶�?33�5���+���s�N�a���*|q#��ّ/p���������YѰ����))����~�z�>

�u��LG?+�4yÕe1"[_�:��ؗ��ఠL��K|���~�����d^����Y${��s���r$���B�8E���ڿ�K12������iu!�Ѿ"ɨ�z�:@ʨ{�C���kK�=3�.�(4Y}'�s��<���ǡ�ǽb�ޒ�}@����TEE⮮�ƛ#Y�00��j�Օh��m�m���V�X��]i�L��VIҺ
I]m� �Z�K�>����Ad^�,�&%/;GC�M�W��ÇG:�v6* ޳\�\�q7�$|F�3�B����S�e�LÔL�+��׬��$aN�+,�����J#֗�~��Ԭ�$������kê�n���jl���΃\[[[��ө°�fٮ��� �N�3��Ԏ����\	?	��@k�&PU�x)��@�eo�d�N�w�W�_�u�(��E}U�VU)�l(���F�t�+{s7�;8��y���x+?�w>%�����C2���y]��{]������ci>� ;a�z	��u}��456'=�����\U�y<���0Т6jtv�����p���*)�JH�ډ��}k�q��F�"Q�8��s
�K��zP�S�1M]*���9<�sx�pX%|8"Dn��}@as���O���A��v��I�+_R�=YF"��&K`0������|�X����İ��}��ۣ� �T�������ak�%���<za�/D�C^�ĦT�	�ӕ�;�Ƿk�G� �%0��C  /��үG�����>�4���y��Sj�����*��� �>��K������r�}�<[��9�s����q�9�@	��� �U~�O���MepQv�/�ߑ�]�#��x_�눏F4�ԝǫ})�B�K,����כǡ"Ͳ��k	/�dI�M��Gv1�Y�6s���߻[gf�7���0��!�dD� jޔ#7�=��M,�=�ȋpj\��ƭ�w��C+�˱���zsc�'�w��Y��?#����U�)QV���*S�A�acE�j����ˆy�ʊL���s���C�J:� yW<����^����{5�}�������{|3�4��]��-(� ��v;ض���j�.괂0����r���2�bG�ř��Lkf��ߑh�����,�	mqt��ݽ��{��]��� Q������Q"��
I~�ZF���l��i��C��.n雅ke��z3ۆ֏f<h���q�ոl��!`p|9������jK.97�{��(KQ�QG�~��b%��&�o�V,p@����>�2��'0UeDp��Vb�
�.
Vcyji�^@D��j|lw����	Ӽ��R�K�\�kChq˜	T��5
�Y�8��[7$�c�zHEme~�2�XT�+U&QPK�?+]8�9d�����~�Z>�B\�a���W��dM[��]񔉭_�����@��=��u����M�+�H�]� �RL�J"l7�^�ť�P�Ρ���ή-
�'��}yu�sR$<��7���Ogee5>�i5F�9e��ё�����A:��SfXs�~�����l�n2W�Y��������ч襵�h�N�����`����l�5��}�0N4&�ʚ�>��y��]�0%��O���u\�󉬫�}nFK{\ָ���ol*�,Gv_1mU̞:�د�A˗�Xe�E��xbZ?Z��[����Y��:�,<ד��7+�OުI|Bo�?�r�������u'�&���J��A@��kw��Dhfff��tC::d���?�d?Y��x�G�i�"��`��(g���.p�{�=m�6.�_űURE��+��f�jU��_sI엖#�,5����d&��yņ&��s�6�y�����"v�͵�A�C�7����y�t�f�����$F�x�Jw	%%e�ޞ]Z�_M�z��X�)�1�|��b��:=t�gC�оz�5��6K -Fﱄ
xmew�5�BkS;;�"����"^Iɽu��\��d<�C��?� �V���A�M���X�ɇ�F�5KB�Z��C2�>W��f�4�TrϠ:�f.,T�o�A��2��w�S��6a2�u/�a�����c�!cG�:�@�4I��M����#��+i��y��Zx����j��o����`�%��:���+*z`������|J���:+>q���mku����s�����?��;� c�X;�,J��������}��:��kZ(�E.N쐀4'ƽ�ӹK�1��\�Xѐb����<{�[٘���=_�s��u�]��M|��*���	"�g0��E]����ዎ�1qu%�[����{�����dՊպ����;����������j"��<�
xbē�닾C��K����cQKKKr���f�(�4��׀OfLS���$�����V1@+���J��(֏u���U�1B�S��"Kid|��^;�g��OAF��Yѩ&Gj�܀a���p�����NDx�9ǎ�� k�l�7k��$���V����D�N�����沖�ӫ�"Cb������9��o��&��E �@�rZZݫǊ�X�P����<N��+�Ɔ�2�
��{���$�'z6$����Uc�g�����is��T����p7��ZQ����]�`���H�0)��wv��HO�1�,,O�0�Х����u'��&�e����C���p0��M6u�;B�X������4߽,"z��l����c��@�2���4\��2����\AFW<X��*�aE�97?����M����ۀ�y�T��d���K(���+�S*�i;N����4��ۭW[�>cT-���=�T��o�QS��ZO�X� �kx�h�|�<8�1��0�+96�D�6b�I���ŷ>�&"w[��"�59���{Kb�q6d��ϒ�v�.����X;������R_�A�I�����"8�5�#ʪB?�Pbb������� �&�t�yC�#�S#6̓2?B��T*o�)�q�ե��`�b��BBo���(��$���r|�b���xӽ���Y�wn��O��N��J	����l+?��Ze�k�P�ǀ�?+�&��ٶJkI�]sU�UV';�5�<S4�	k��¡kmZ.�Q��	6���)�$(�ܝ�;��_%��6��b�$n����	xA�pF�A����|l6��k�˗��R_LH�07`�Q�իY��L�u�*�u[�5�u$�c]G��h��,V�7s��zH��H�6Q��cG�*/v�5$U�+��U�V{!o>χ�z֖i'����J�P�4���^!j\��yD�nE��|��|]���l�n@׆U�[�����o�&�$�x�����03��@{��5���9�)���
�q~)�
����C�W�� ����*��S��_$�Zd�W�;�!)R���٨N'�Q%�h���<�)}����fa�BTqi��U���B�Z�L�y:@�fn��U�y��[�/��	�%PR@�{)�`�\׿>_��L�:�"[߱,G|��&m�p�y����	� ��W~��E}�O5������ȟhOi�6R���% ]�q�S#U����ٷ�C�~�Z����������7���4��)O��Rebg��N5	�G�ޔdhDo���p��)rk�z�2+pPX�+5�j4;gΐJ��wp��%���{����B�,%�qc� �Pd�l������H�a��f�W�v%��q��/#���W�����5u��ҽ��r/"���cM�����x����Z>˻���T_N�ʎ)q���a�8�L�#g��>�É/���Ȓ��<��˄Q7����D,���9��u9�J]Z(���+���9s�{�/��I�
��0]��O^��]Ґ��-(C��rN�r��Agi||w�ʊ�����+ fP[�a]�R
'j�{Z�/)�����R�'���6����Z{-4---��L'��ZUm��J�H�C^
������stx�TVKg�h��k2��d�E�C��}�٘���D8��I���Z��s��1H��@+���A��T�	kζ��nΆ�fkμs��tL�Zo�.Twl+|{[pt=���a����}�w��f}�˅�rᇜ$ZO;M�VBqzC(L��]��G�X��Q���h�`|�f�\�dj��uh�U#��`^&���������ȏ/,`� �U3��F��y=h�Ն�����M��ʋ<��h���^�6:KQ�:j��LG�*_�"��d�[��;�G(_UX� -�}�H��V�;��p�JK���#j��V����NK �m�&�<T�Y�@u,/�0��Q�-*<��5��s�����dǮԺ����-f�U��\��?]"6~�Xx%�/��4�*�A�Rʕ�{�����	�1���{��\�'��Z��"%��X��d, ڑP)2K�]ل�u�s�>���ڐ2��C�܌���nh)���n,��?"�f����	Of6��<���(\u�HS\5M�����hzf;E7OQ���h�1�/�?36��;R���j$�g&-�<��Jz->�_��"/%@%S� ���Cq�"�~�����G�Z�1E3�H���b�H�VE!�Z���Z4c��E�� ����u\�w��=C��o8��)�� DӰ�Hta���t�1�FSl�ң���G�}�����^d��՝�8�rƥ���7S�3�2�J���b�����;��}{�x�|,���C �_�M�0ˍ���ZM��,�V��ǃ֋�Y�ӕ%f��qoVxL)���pf)>W��ш�G�Bє��(i�C<��m�O����G��P̓����H�6x]��;\@Tk�*��U�D���)9κ���Ʀ����B�.��������f�3&Ë���8�/�F����{��J�>��v ����z;*��i&-�qd`�H3�2O��C:33llT6�[?J�!�Ժ��[B�㺈�|Z�5�^^�d53 S5�U3����%(��z���(�2#��;c6�?���a
¸�C�� 
a�/�Cc�#�D���ゾ���GN��6q���go�5z1��C�c�su�����[�3ěE(�]uRE� �����<p#��tQ�-"�5�r�g"��j�iD�6J�$��@���Y%��&jj��^��y����{J0�v�꾂�����%:� �Кs�Z�������!���nbҽ��ISz����8v��WV�<R�K���#-���w�aSp+���~�;!�~l�LAc��}	�6eh@W���S@�h�AΏ��B,VW�4&\�Oe�
�^`��Ku���I�F}B�^D,��%�]���W@��'{�>��Η8̜0�\��;J�g����G�-��9#��/�P*����a�ܺ���t��J�A��`�7�V�*�}����7%���V��k���0:F�B^�ހn^S�=Y�K)��$�3}J�y�5�зRM�QrTs�L���9�S덯`V/ j����l�R�
O���x��������L�Uj���ʪ�vr��f鰚&��x��9#��/�����n������3��:��}����N���i�l��;{Lg���De�`ȿy}�#h��KaS�ౕ�.g���g~�ϛ�5xOF�ޣ�5dăi�y�*��ix�Pv0:j�8:��,��5&��v�.��o&�;�<S$?u �#��-��B���Qt�Q�&1q%�zӈ�о�D�����7L�#�b	�^눂����Ϯ�bgG�Eʟ�x���2��߭�}��g,>֘��9��n�z�Cxu*:O�M0\��*MK�+R?#�N�w � ���&;��>+�p������ݤh����֩��Y����M�807�e{�E��0���Y�����Ԯ.=�&��?�ڨ�'������GJ`�ރf�|�����>K!���]�ֿ�U�^����rQ4���� oR㶫]�[�t�=��r��+7x.�Y���|b�$�KE&o룑�_���D��Q���x��q9ˋ"�y�r��*$Ƿ��3����hk9�N'я/?^zK}Kt#�C���#�e=����_�k��y�O-���̓�kq�w�@Ms]�zm?�)D��:*!@��-~'W>��z���|�KwW�z[�3\�nd�]�z:�y�*�ХQ;�#�	J�q�i7�Ď�B�,�%X�윃iD�^�W!�nW��&�Bg��k��?b{n�A�hp4�i����t[�xNtXU����^�w���G�	�>�����ӷ/��7t����Ƅ����Z�h����@�?�nJƟ���#�묵t<����l˽��9�=��i����r�C�\d��%���!u7I�7��&����q��Ǐ^��JC�P�(�)>�RO
��CO'R=��.��ȀA�=ww��T�țD��*5�2��O�o�|�:����L�7����l��3�d�����k��n�����;�p��:�ّ�g[c���Ƒ5S�O�	�z�7��1�%��a�>N5x̯��0� 1(���
���G'V�R���`c���;���	~���Jn���o���@�����]���owB�+u>�˯���~Zq+-�w<����N�n���$�!��`�\I!IE]}�4�A���hF��5� ��#@��vwc g��_��w��[��h���k�>��@F��&?�Y��p!��k���"&��Dk���'�Rm�?�^�TY����V���no��'�nIO����},.o����~��h���5�����Zmx,��t��_
�"b�Y���9r��4�K0��;;?ЍlOa('��a&668���2�U�\ �/
t��,8a=� �"�����\ JG?5�\;�0��F�g=�ߛ-�䨢DE�y���oI3?Ĝ�q(��We�z������\$�y���;����'���eF}�����qB^qЏ����>�X�����3�#���,@��#|�N��*y�4����D�! 懟T4���)�>#���t�w���eqU���r��|#QKwrQt.9�0p`�u�H�j����EK��ꪞ�t����� �,�_�17�Ch�g� ��z�f���Qo�G�TA�3:����䧽f��b�0��B� �ɑ�F���p�ќ8������v����i��"����,������m��\½�o�1�2�?wS֣�RA���梕e12�5��<���z���6ΐ�Q"5�%x��}c�pz2z<���߭ol�����f7�2������ϰ4���p�LD�A�þKYrn������+�(շ��i��]
b�2��U�ѽJZ���U���U���X�/���g��п"m%�+WA��do�������\����<H�P6yT�Z��e;JT/7�ϔ��~��>�wI'e�7{���j*���Gf�RcŊBd�%�+݀����8�Qj$���k�V�����u3���=��v��X��Y�.�t���O�2*�y����$[ z��s�Pq)}g�Ui����%b0�g�<�)�"����K;�H�'M�>������l��_�:�Y
���r�쉈�l���:T����8�"Bh�\ѻ����4��(�����,�}�w>M�\�k3���}� ���}�Ө��}Ң}�3��z�7]-�J�
�|>BI��;����������~�)x�=�,��d�Ш�gb{N�vL3~�yD����h}��|u�.D�x��y��{s\�uDW\�Ƒ>y���!�A����7���������������7越	����c�Ɂ�|�UPh��DB�"�p��Nvܲ�.�<�� ��OJQy������%E�	��������ibh��}NgG]�� �5�n=��1�қk�VUm=�{��͛�Q��h���j�{O�z�4�W��s/�������\��r0�_���G��y���Cv�Z��|����~��M�Y����{���KÜ��˹+�qP+�l��>�<����rh>��	d��1�ő�i�0�����9��.��i�n���vdH��F���Ҹh��G��;L�u/�K��X�hW�@*u�NSd�_�g7L��mZ�\lF܉(%�~/���.e�����.���H�p۫����1�E����w��+Қ;33#k�V���f����<˄���߭��CV�]���ڿ��2w?��.3����q;��,���ϳ]G���Q�	�I<�j��X�j���c��S�g��K��\T��7.�A���7ܬ��pg{�R�,2�H%rp6�%��e�~mXUڦ�y?���Ԧ�7��{�z��5��A��Ş��u�C����r�8X���"�]
�=�y��g�vh�Y��}��窴RԞ��q� �0�G-�?Q�Y��&�$-�r]-]�����p,/�݊dr)u�}w^�e�]i����P�O��r�����"�����bd�]�v�~�:��|��(�ٛ�3V9�Fw�F�~~~�S�C�(F��խ֛�񪇿U���BA���? ��;c�������T��2��
��$�������vg�IiT�I���7թ]�we�o�Օ?��t�*�/'�n�,C�tq��r��|s��F��]��p>��g��z?c���s��5tw�<���z%�0���{�w���}|Zd�T�dk�dKvCRyٷ�]�5�2�X��Y��ɾC�A��0�afH���`,�3�ߟϿ���㺎+G�u�����q��s��?�T�L �������.ɝ���$i[�)�w:����&�k"v<�#���<E���+�<�@���"ń����]'�2��2��Ee��V��aZnb�ɵ+
vVIt	�wzo��lɚ���C@���Ľ�O(ӏ���T�x	`4��gS*�Â�*�Jj�Z>�������z�7Y^*R&������t�ѵ�dJ�EF���G�N���C�C�EOU1r����Q"+�.�%���;�AF�J6ՕZ��Ѱ����Z���Z�:M���v�r����G�-��	r-���Oq�OJ`��͒�O�GW8�~��B
�j^�g
��M��#׎{oOvXP�|/n_��r5x)1��\J�֪='��#����l�O��7�IE�oK0'�BE�75�%���V�D��K4��$���;��c��z����!�F���s��^�GHKq��Gn����U��Θ#a�?��`�B�`P�Vm3�����Bt��F�;�¡J�7op��b��(G��S�W٩�J&I�{������F1n� ��N\��=,�mt��9�륐�fĘ����;X�YB��i����<�M�/�h,y���m�ݬ\�}�#��^X���J�A������}�#f���u\(sU��`+堌�2�j���G��'"�]9��\��/�����R"�/�z���Dn=��Nӗ�NL9N莁����k�3�]��\�m;P���p4�Ag�D��b�����{��U�{8��i��l$C)��o���j�O'�فWu���湩���8N/�ޟ;a��C�ƚ�"J��-����:L�lu�C�R����ӧ�gK�ۯڙx���i����>/�N}�m
$E���薵�����$KyG��&�O�L��Ծ���3�:*E���o���z�4�ڟB���6�d?�]�.m��)w�W�+�c���Fש�����f�Y����o,Մ�G�C��0P� g��ӣ���=mՠ�����"i��`��E�Q�����8����o���.~EM�ZfD���t�k9�]�SjT�4���D]�l��j�`T�UZZKŮ(W�+��o�#��5�&&�o�������Cl��H1������xcQ��̔�����G�kuΔ�|}X\j>9�{����Ψ������=�PYm��hwf��]���7�UKx�����2N������ŋ��ƨ��6_l��|�J 7.���s�8N;8e}j�eۿ��44\���dΫ~������ �dQp�[~����ZJ�������2[[_Vڙ>���˛P���9y���X��Z�\��˛�;�5[�x��e�J�ͧ�Dm~�3��&"fB��;sO�&�q<�I����0gH����}������ǽw��%������=j_�Q^��k0��y�f�^�m]�j��ct�ˠ���W_��o�\Q��to�'���<^�\A����ثdI ��;��ӲÙ�q�J�W�R0���ITF�5�x�O<����L��Q�M�����3G���4��ߝh\k��d&�MfN�N72EO6NF�w����;�rzNDm��g��3��	��� 3d?!<�5�]�ƹ����ѳʭs�A<�L�Q1K�J��N[�V]��}OI�eߒ�X�b��f�۲��
�u�M�hf���R�v����[\�� _#dJ���$�>��~������n���e��2ۉ�x+쒐`����5��M�<"R�vz��ywY'huZKD��N����ͫR�*�T�P%Ƴu{>����p�혡��RG<=f���6��
E��ƜcԘ�)�x^X��k�8<��a�#��y���)�T�F�I7�7ܥJ'f{_,?({����C���G)1���,:r�r$��6_hV���
\uHZ�,`�13�/h��2�GF=�o˟(���V�h7�*CV���ƸwR��l�FK�v�`w�5�Kz0]+-6���\�}���eN��,���;�FU��=7�)����q>:��ʦ^���u2n�cւ{B��?�I��܅{��`N���g�%�@��h�Y؋k�G�ΓH�1[�E�TKֶ}���$���c1ȋ�!���+'7��+�!���V�7B7\1�-��&�ٳ2��h���#V�U��7����+>u����GR�:J7!J<��a=1�n���9t�����\t�1A2/�D"��w5����Y.�
��bA&���؛�ڣ�a�%�lx�w'�yv�ρ�������kT30c_-��a(�bPC>�3� ĳ$ ���rr�O�Q��e=��ƷZ�(z'��>�Yggר�&�7Y����L����3�7��(%D.���������^	�S���g/�%
��GN�.�m?���4��?1��t]܅71��#���K�8}�r�sg�t����q��됴��dia6%P��������0z�Q�r�so��x��j���I@�������:��zzz�~)`�GJq_�Ǫ�1�V�(�g����egf��Rm��iŽ�mu�7SR�k�f��q��sݝ�@j�)Jy:��Zx!f�
���@�c72O�
d�Ʉ5u��6���繧�a���qLL2�Z;^qi�T�Ԏh-�#7ye�"�|h:h=ݨ�� ��Yf,}�KFA�1g^���F����}���c(u�{d����|k��k�W�����74���(�Ц<-�@�$���ё^�9��K��T�ݨ����ǷC� �(ދ�o������Dey�<	ɭ|#9{HT��+���G3�y�It�|���f�����Ta�G+[c͕��qKV��5?R.�>����陰�
ܶ�p��:���w������t��7���}4yn�����K��_\wg`�O��y���i:;葑 ^1�2Уd��C ��.�����B�<�ߟ}oYr��'ᾶT�hװ� ]!D�(ٕ�n��UTC3��6Y�ut�̸~�����|kp?�Ս�d�y7֐d!H�yP��E.�x��m;\:H���Qא�tW�RZ�S���}���c��T���z�5}�1������v���UH_=F5���:E�껜����
�VםI�v�_[��� ��'f��"�E95��
��SLx����R���_E�:�g���x&F�ly�_l�f�-��R����w9)�+R86$u�sF�~.]�R]`��a�X́�ZeGf>V3?{�Բ����4j�����xA��d����"d�9��c3#�ל�K7�^s�to�};�FQ��z���/�(�K��0(������N������x��jq;N1�ܵO����/�1������h	(�87��qj̦��4q�;�(b�5�f�����[p#F�����
�,no�8��Xd������}�2D�I�b��0�Ȁ=��j�_��0�1�]dt>B:x���S��~bߋ�:E��j�*t��J��$��_4A#}�������C�3�)�)�H��'�M�lKc[��oQ�#˔��Ѥr�M-��c�s:��{w��rbI=�xt�;�%�M�-�9ҡCE�8���ޱ�<"7p%nuƜ��d���|�������R�1��v��ãu�'���r�f��x[=�*�����z�y�d����w���\o�c|�x]��N�(|/���%�5T:q�T�M!k����� [}�Jﶂ��Q�kr81 �K �}��*��֟�5K����{z����F��|FD��fO����W��dmr��>��d'��΀E��*q��縶S��tR�7�X�8�<vq�X�yA#�����z�:�_��,�bT������������r�j����36e�8p0r��U%o����C@w��~Gw�P��ss"�g�ύ������h�2�}��I�ȕ0Л�	T����e��H�"'HH����\h/G�iX{}ߚ���
~E��[�Cڢ��K e-؅�h�]W{�VՔ0��l{}l�Zp��f������X�xwXQ�x�+#�)�^�G����M�ɾ�N6�5��RP��D���[� ���|sTm��������17o�~v3����z2�dӶ�^����׷�;. w�*��:���L��.��i��w�R��ɐ���(�&��?���8gy����?J���(��@Uڕ*��rt��%ye&�<U����Y�Jh�Q�6��[�Ԇ����K���5��.�x����N�>�6�y���æ�L�L��i�I %kX�a��F��x��L]���w&�d5��^���A��t}�3;��(�T4O�4�aF�����n�ѱ2����<�2P_�s�6�s8���4��Z���ӟy+�&��I�������.��X���u\@�{.��Ǐ��D*���O�����PǗPS^C��撒�X�PFs���"�C���(r7��N�����E�v�y�)a�h�\�,x�}��fUc������!&��.���	�j��y�|�x�%����K�.2*�,~�o6��S+��@|��T 4 �ig��x]�]��I���GT"��s�R?JU��@]SF�@���ޜ�����(�|����ٹ���i0���)�J��u(�7Y����PÇC�,j��b��Q;E�|ܵ�<��Lۖ��	���=goܳ�����^��-�w�Y\��j������٭�ѳ�@��4b�l.^�,�3�	�^��&�XX_,��Vjoq�j��q�G��Y���uw&��"�k�6�Q���ޮE�Ꞧ�	)���O]�;o���╈b���dp .�k�5���V�»��k1O�kܩ���k���d��B.���n����^�-�˖v2:?�L����Z���σ>��FI�� i��q��C�E��+�� n0�>��^Zz���}��\17w���y]ݸFf��D��(Q��ت�#�9�f�ߧdQ��ϳ��������FWi�37��O�����0U�^���O�ŇFt�����B��ǁ�9�t���4�0Ͷ���/_J��VՐ�;��\T�!�y��ǽ$W�(9%���s�C@�w��3�ΞED��x��p_a�؅���xʫ=����U����^��4e��"����
���.s�TK3�A���j3ujs�|�QB W���6 mn8U�FRkF�(��{�~�5��X�&j�H* �)%G)����k�rv�ZT|�@��.��q�����yǷ�$��*�,eaC��G�
b�3N�9��Lsq�$
�nP<NwJ�˕�̍{�����k����kd֮��t���v��<�C\�[S賽�Uw�!m�]�R�5>s2zu�W��tܙ�+ļW綋���N�jI����Z[^h0��Sd��4������v�A{���*K<�c�G��+(���~��ڴ.#d2�[�J�9��*[킬C��̪}�uG�A3@s2��+�gc#��^<_.�����3e�ͨ��)Ow\͊�u�t�[v/��/e��+����'f��o'kܲl����h|���W�EX#C�!��[|Y#e�����jA��&99��f���k@TMTds��]PńF2JK6�����)=L�,&��?O�9G=F��A�UPxG�K�sbi����0u�ƕ��BnSvb���`p�`_)0�v�o��v�΍�r�c~�*9C�'gs�����:��c8__P�2;Y9
�1�� ^Q��3�{$ò������G��J������O�Գk����X^�ͬ����dOϦ����#�PF~/����+Xn�O�An�
����,x?q;�̉u6jf�>����e6�#;`z{��ڬ���4���h���D��r��|�ƶ�����'ƹ��b�%�!�o��:�E����}d���GW�����%�r�Y�z�
��`c 1d���fn��n0�6�K�ʵR�xr�)s-\s
6÷rm��1��8��vQ��Fw��K�RRL����>_7��t�k=�I6���p�!��h�Ӽ��>�ĥ�dvMu�\�O�.�|�/�m�i���Uq�7� ����E�pV�@e'XL
m�w�­t�KsrG5���Jv��cZ�����ۜi����'T�SI��]Ґ��P�@��Q�x�yH�����q�V��"�K��M5�=�$"��v�>Y���*�]qj�S�{���� ���%Y��������v�{Հ��q�_kU�E�y��:���^����[w
'��4Þ|��æ��6Y�U���|����Vl��"��H���)g�v����l��8�]��I��c����h�@l�K�p�b6i� ��ǞkP��b�o��9������һ ��<��1��+-�i�W��v�ޒ=F)��璗jI$����Ჶ��G!,�j�_�eX���&���$-E��.8A0BM/�Lc��R�0	!I���)K��?A*����;%]B}�"�D��{����)u!x�*ϰ�`m�v1�9F��i�)��X�ޱ8��L�0z隿QB4��ȓ�.}y�i���m�n(��/��X�	�No'��YY˩������3g6!Ǐ�45jd��� 	s��*s����Z�Mp��~��'���R#rP��#�=�&�rA%�2��b�����M�3����pghK俉����H!t��/�����i�]�:���DXi>�5=112�{��XX��7���|yJ�^����@��V��u�C���]=H_�~��V:�V���"ѼL���į�`Q��$?�ɵ�M�0K�8�Wc�����Ek��{�hSq�t'���@�B�7W9e��#�.�yE�{&l�m�d]3C���쁋.he��O�&N��h�v�l�[8�� =���6v���Ks�� ��+@ZeS�iTi�11yG<-mg�[�e�L'/w1��W/���r��J_�K�哫uS�G�J�'�\��������j�|���.!��C���*������	䒍) �;?,���\�ԛl����O�)�Rm���s��n��Q_�4�y�jˮ P�`T��D���-�4�rF�^�y��ِx��:vgZe�<S�˾�dı7/q�y#\)�O]�zj*��.��E[�݂���	֏O��P�dDѨ�Y�[�%b�8N\j�s�5օs�aLF8!#4��%����ҖF�����G�+/$N���[ފ��)�H��=�:%��?~��;��i�Ӭ�@����=<
r���z�FM偬Z�f^�ȋ�^�qiIc�C��_��~o��&�{y �t�h��r�� N%F��d��ݣ�y�n'��?Ok�\��R���a*�9�$3�4q}�3�j\���GG�����=����{�D=6��$J���?f�"��uD���3gn��L��9b�-%E�Z�G�[�b{Ez�ywT�I.��Y�ͽ�����_q�oiԄ�ׁ�;���0�7Yqo�~]��|��Hcu\�پ��r����61v{h-���x%,�!_�!��j��v�X�h<Ak04�u�b������7��v�.��qf痹�;���Zs1f�&�}�|����"ڡ6%|u��g$����s��������w���{����;�酯�3�����i�$����sL���������N�V�J�s�Cc5M9����ߤ�s�|"6��Z�S�M��SN_�g�sn��߉�:�9����`�m�����y�Q��gB��8+nْ.=��Ҩt��{yX�DE�<��������^��ύb~��#�쨂@�%��G@o=�i�(�t���W^�Yr-��{����og����s��+T7m�mB�U�Q��G��1{�~j�(m���&���_л�(\GY��.�ř��j1��WJ#�']��>��#�7��x�A�c�Q(�w�Y5�E���o�ԴRpi6S+iǠ˻���yQMJ�ck��wJ�_������@W�	j�
�����Т�P�I^��m~<���<p.w�Z���>R�bv8��(G�0_C�l��ecH���ʠ�I�kw��)K�h�aaB�T�~q<��Pj>�/��YH����}>�ݽ�7m-�J.�6J�a��
Q\X���r�w�E�Y�φ����u����6/ь�l|57�6mO��2F�=�����Zo���� �w�3�wo���T^��>�R��E�_+mg��������b&h�~k8�Q#	���/�.��43�0��W΍���O��s#��ʕ4+})�C�����wE[4�Oj�yRQَ��Ou@�t�"��Y�P7�F�����������7��<8&�&��(�@� �+`�k�q�:���D�?�J������j���%s��]��W�
�M�D;��[��T���g]v�nt?�E��p#;��_�$��^��)��?F�^�l|�I1ǉ.i��7�B�K�<�Ry�)"��� Ї�R�@��cd�R밉X/j��%��?X=t�[���������u2r� �k��;x�G�����޸J�J3(9����T��)�Ƚ
���ݽ�n�Ҫh�,����%kC��W����3F�BI��������ǀ�V@�}�+}P5Ȑ�o��Q#�c�\6���?vЅBV�G��j��)�hTy��J�e���_I��;�w��_���EW|��b���ޝ����.7����F��!)f=$��'��<�����Si~���S��/����✰XH�5�Ԓ"��zTz=���z�/��$#<��h*8㼹���!�~V�<k�1��#b̩��r�_���f�
`����A����6��̪�n�������oB�2���9���׊���yl;}����r��a�~y�C`�h��&� &N�@E��|�gN-5֡�1D��v5� "$�����hcO�yl3$���0]��i�޸=�����I�ь����u�c�Ϸ4����8�^��ƻ����#U<UՈ6_���L
�Pq�M���,]N�kW�oQp�rFG@&,�ɕF�o�{��F��l�;&庻�/��O�h42�}�;3jbv�N�8w�,� ޡm�'<]b9��!W���߸��7�4OzF���?�E�}��{�F���8��H�<�Tݾi�iY���j P_4`{�S�����i;OFaYR���GRG7^��<����d���)��>��R~�c��sriMC�k���p�[��?:fq�u��� _{0�"B��If��o����	�r|U,ߨ[��%vd�<8�Ս�0G�fYS�����G׆��6[+Q5B��i@�ʶ�h|��xc����I%�ߢg��T���=l��s/f��T5\��i��z���},	�w��}�d�b�T���D�	pj1?C�jɲ/�=f�ߥ �a�O���n��ve��7g� ���U�Z!�֠=� �Ql_K`U:ֱ�����5�e@2~r�S�>~7]d>zr�㜉�
8t �d�I.H�;�F�P���ZG���e�)�>ɁqKP���Gh%2�L|�sM��o�vI ��[����Ļ5�`^E0�v蓘���& �:� ��N�g�lB�k�|/�ǅ/�mj[}~��B���n�?Έ[�������*S�3�.���k��������Uܴ�^�c���j�qо�?�K�i�� �"�=G,a�)k�������ޟ���e�?*�?3m�'�{�h��;)RU�������>{;�+@���',��]8Du�I#�1Q��f�+�nn6er�oZ,����,Bl��~4�|A�{�{����	��s��#(k��C�O�{�=]�?<�Ny;W���U��s�A%�w�g���/�ܕ�q�G�I���t�J�Ξ��X,y�}p�x�j.��;��Wt��MwܽKN~7ۺN|fq��(�5ѭ������v}p(�I����{)|g���>���<������lo*�4�U�^�3E���"�V�]��3x�3a�-�336���_����?B_U?9���bz�?c�����3$�u�(����^[{of+�h���*�r򅆵��2���Ǝ<8���/I�Ϸ�P�~�(�N&�?��#Φ��s]��Y�^�G��*]���Z-b?��޾�M�֦�3���������Vw��;�?���@a'�u�G�:��x������~�/���)h陱j}�O�,���5)�J��e2�h?�p�������I����T���
�8�ϗ���Pۥ��F-�^E/�\Ux��얭�6�|2�]���ao�����!�[M�������;y7}��'jMN:ʆ��Ǻ~�yJ8ɾ|-Р����D5�}�Di`����[4�L�6�L���g0$v����K�>��j[���kV�w��1�K��K���J��ط�'Iz!��?����P5^j�䋿d`��1U3��yNW-�Jq�m>{���G)yj}~�ƃ�ǖ�'�PI���Odn^����i�Sx��n�w�,�h1���d�X	�
c�`��C�����eghX/D��@�6}p��kxi�)����_b+s�ݟ硎Iv�#�_�!YQ��^+#Ʊ��N:�>����y蛯ac�Mݴ����Cr
ړ�&���T�-�pL4�0�A嘠��`O��!1$ǆ��_eX���;U/��o1w�������`X9bv�͌�mxFf���*�4?���h,���� &�ľ�z��Ӎ�Gdv1Ky'U�#�k��tM\���9�Hw�O:T��m�(R�:�m9�����PCX�l�/6��|�Zn��Νa�I"��FD�\ Gi�� b�l���`�;�	hơ���1P;s|�?={�t&�s�����A�3��ƣ<�}�mVݪ��K���Dֳ96��8�M���O"m^t��X���}z�s�D�ΛJ���@���q
����@�tu�UY�9�zg���'��I,v��^]��wAA�`�h;jx�>���#֬�N+
"aK���	�R��kԜd�c��:�jcS}3F!BWUr���n*�<nH�P���fbn\{Rk�9q�#d�Z��VH$dl��X࢟:=�u^����ˠb�~���!����m��N�OшA
��0�NQU�}G�m1��缉�q_MKg`��>��w�ׇgQU[�4�!�t����&n���o�qX�^�8r�F���y~�n3��P�|
�u�"�|�;Փ�BR�u��r��rl�j�U���q��r�V����p�6���ZPC�ϗN#S
�n�)��߫��7w[z9)n���;�'����'���zv9W���\�K��<kڗ��m|�ܻ.AWlOy��,o۴��ݼ8Pc����������]�h?�fm��;�ƫQ�����_�Z��_O<�Z1�Z?�䏊Ŭf����d>\�\=pv��j&3�3��4��2���z�tFs����J�5��I8���/��q�v+���W9����Y,�ʈ�_΃/�B(�Y��sW }�Ji �<�z�~���`��
��$V+䈭	����!�%<�x�#`�qK��3-��5g���ͪ_f���/	{���L7�0�^��t����i��q�{�����ם�TP�r�t���h����-�r��d�Ox+���U��`V�Y���CJ�tcP�$�}<� -��J8+ܻ]%^�X�R��n��W'0��|Rc�v��w�*ξ��A6�5�֕�/�������
*���f�Ϡ�����xh�C�����.֛�qs�V{���sk������ABXe��幇� P� k���^�mH�����Yδ�o8���|")����o���V)>S�0B9v(Ru�Cqm����_���K]��!�bo�߫�Q&RG���sC�����"�iS�;�z	Ǎ���E���#s��۳o�
��s�m����[S�p��
 P�i��wZ.h&�36�J;�#��)`��ת���D��P��t�o�����.�Z'�rM���e�8Mp������8
u���#8�OX��q�!�M��e��8��G[��y!��B��I*��5����f�i^]�<03������m�Բ���ҫ��Sh�k�F��O�h/�W^�����X�.fM��؅����F�9�|���J'&�f}*�����������9�Cr?d�ޡ���5��zz�f��< hX��U�VG3noM�o�����-c���~��`�^Zd\��c�Te�M'k̨����IQݫ��#��6l^����[22v���$-S"ft?�@�`���΄�"DG���HE�)
>���^,l�T	'�H�2�����Bg͐�������_���ي4�k�B��E���r��g�᳉�GB�ֈ�
M�}W�S[?���sCF�?N�}#���E�� �T�,����T��˂��CP\���*}m���|U~�J���6�z��/lO�|�YbY��Vr�A��,�Db�������c�ZzŢ��i���	�N�_����N��20�Z��v�	��Q˲3��	��*HO�=���ǵ9k$��"T���a�=���)ߣ�3�a�m����T���j�KU�7��E@���l�P8'�g �@r�+�Z+]��%��w��m(V`4�hV��?w�P��紗w�Ka��[�����g�֞W�T��s2۴"��=L�6+�6�:;=�FG�̻)#�h~������<���\؟�Dޕj^X��&�U~�lr�.SFO*O���Ʇ�d{��W�~A���%lt���T�3��#���C$�d�	������U�[@�������t��L��gTL���		�xN��.Xӻ��j{�=��X���c�ɵԦ����@e,��2�55��]պ���<+a���͗��h�õ�2�cp"_�N�+>h�eV^��D��2�߷�A
�r��1#`"?��[��%�;���6u�֜؆
��z�c\��<��ُ��4��?��|r3h(�F>��U��G�,[Me]_\���Dy��|�K��'Fa�l�B.o-�'��pU��T�-�(h̕��l�SN��0(�m�p�k��*�JI�UߋY\�WKe"��������=ɺ���֑-���y�"~.��^�M�4�9��5}$eO��93I~���asm�ax�C�� 4w�V�z?	��I0�;g�y���>�.�o;B!���׏������azz�ٿ������H�慠��������?��fh,�>�d����;!�چ��m/l�)R.�X�=�B5�!����qi�A�{�C͹�����G��|`�z�w����~޵�o�P�MJ��;?<�]�0���Y@RF7�1��|5H�Z�j�3����U���Ռ2V����������L�^h�<Tl��W7��3>.�U�kqJ��~s+g�d���ա�O��f#��4�5�w���d˕�����s&���$�+�~�FI,�W����?���+Mq���J��Y��p��R6�_�bUO� 0����ޡ6q�
�E1�=V��#u�(�wuy�Ԑ4�Ƶ�3��r /��#�rㅬ]��̹:��M>]�T���&Ƥ@����O8ú�Gg�J�G��"z{��yū{Z�b�Ү�����r��#	[/9�z�~(ɹ��e��$x�Ѯnb]�������!)�mF�����C�:|	��;Y�P�o N��>7p�k,����y��8���n�u�Ϸ�|;�Ʀ��Q�t9yS˸Ղ2%��!v�+ϟ��m������c�<+�
񹍄�x��-���U�y9��з�f�������`��p$_e�5��Yy3�3	EJW�^]#=F�X����+!�^(�q�w��{�8^����HO�'Q̂c��`��/S���4ר9����8Os���={e�`8E}�cs��T����5@��wX������EA]tS�^�����ɜa<<�t����f�:-��j���I�<�������!Ե�FI�׭;ºW]�,���NV��# �|צ��[��u\ZdCo��S]���E
������r� �U�泩��af���ipo�仕��))4�j8��P9��?�?�Gܳ�ƕ͌[��zȻ���\r�ɏ��Nj!���~��V�����x�R:a��N�%�]�U��F?I��3�z�dr���n��t��UoWB�TB���,�`��8������<��P�SIp;J��EL� u�xL���ƈ�2���e��ϩi�w�����2|v7�ì�l~`�{h�7��$D��M�=H���dh7��?��J�,����!�;��F�pL�cX�N_P�HݜI��k����R�D���������k��;(�8�Q���pN^99�O/,�0����%��ʆ;?��a1]J	Z=�`�:�ֆ����7�\!�r�Ȝ0 F��5�Q��ŗ��e�vO��/���L<j#����y�&?#���G��i��0p����}й��I� ��.�a��7n^ePLM��}�N��U���;nsb�ٸ�]W�3$�;'_msAԲ<�
���j�D�9=�gm�Ua1pb�fBK�Zl+Q��a�\�,p������d%�qq1����ΐ����<w��#C	�T�X�$x1D'�g@F4b�B����7_���U�ҡd*�0��=B��E13ګ[�<Q�ƪ�%��
�ЧUQ��Қ�_  m�b�����{y	��Ma��By����^�=G�'�X		��5`�����kD��x�&.�Dκ�S;�b�o.q�@t�n$�٠v>� D�4z���|<��P¸����o�x(!-���l�4���(�ExJ�Z�..Ӄ/�O�ꨨ{
#qf��������)E��Ʋ����ف�mV�^��i�"�����=q���{HCcҗ�����W�K��̆e�/��T�6�iD�����	ˡ�_�9�M��Y�xF�p,���-Q�zM�Jbu����A��2لQ�Z������!��s�if�v�t��`8p�����|�H=���v�p�g" ��+'�������Gs�E�̅�oP�!x�U�=��53�=��ɪ���ҽ7E��/��I"�f��թ(�Ь��A�5��O����1'|��PK4[�^h>	��sçL����f$��g��{������W
�{�gbk}�}r8|�d��_İC���������6q�ڟ�[&:O���>p+ �^(��N@��.2��aU�����-�7�5����~�)�?����+-D��Cm�r�g�z�p?���K�!��
6�(T��W��<�{��D���r�V���ڧI��@�69A7æ~��Y���PpI|���rL��H��m�Ԧ5f���٪{h;4��Jٖ,8�dɥ!�9�-U_L���ZT�'�~�\�y�?Ͳug���B%���j�~Ơn����>y�;�ی]��6���7�k���s)�<�m<�5����W�>j��kP�"��;�:�2��0�\�8{��5ҍF�ImV�"�Х��(�V���-坧cq�<��=I^��(y���9(Ym+����z��B�`8�*
V�@��B�ɈM����"�������AZ��lP���9e}�� :X&49P+9�~E�lۃٻ#��SQ+S�Z�������qR:��an��$!�XQ0bm��РrգzVY��\�$��zF��n��D��II*����������*�qE��69(!L7u�*�H`e�k=��`���W��v�\$Q	��`�>�{`�u��u��ܒ�VҜ��q����W%n��,���71�WKRO��ޖ���M��|^�XY�Rb;�d�X�i�lrp��[dYX��3��4\;?�%,������/99GX������߯�Q�_��Y�����������Oo�;�_�?����Y��ѽ��N��?PK   ��!Y;��q p� /   images/e9c16099-5161-4325-9ccd-582d4965bc31.pngT[X��I�i��HKyH����FB�[%��]�%"-�t�s�~�~�<Csf�~���z��{�)�I�������KI��``Pa`�v��+r�5{�x'Q)d��F6�~n/��C����PQ.�p�pV�3uv3p4�qssc���r22�7a�s4K? ��������g�Z1K �1��o(��a�`�G��e<������8$��զ�$�r9�վ�iu��]�g�i%Ŭ� �`#�⽌�cǦ��)�vڃ����]nKIɎσ�~z��;��j�y"h*O��BK1N�"���A���F*�F����&?�I4J�64c�9�f˱�q��z���566�������Vg٪=�of��M
��[N�ނ��0�U
	x���/	"<�a>q������Ag�>]�\�ˬ�ǿ��"4yO�[�-ͨAZQ���%s5�镲��t�y��
�^��N�	���4{z���0\:	&��o1#���y�^�}8ȫ�"�6��w�҈`UZn1}���1��r�<��n���ɃUD^6�Z��g��h��aKz�Jk���_���B?o�	�#��p:�B��ə����L�L���-���DӲ���7V��vx�����}p���Y\k]�.���K��Ta`C{�����t��c��G(p|������[��s����P�
��b�����-�@�S�R�O��S���^Q�CvJo���Ñ]����������΀��"%�!�FZ����K���W�0�UW����
@Ta�I��a��n �J~F=�L���G��޺S,����B�yƸz���b���[�p0t����u�}ۿj�f�`<i�� ��!��Gc��l�r��c?5������,�h��sÙ��̖n�UN��G��r� J��1ip��`N�˲�|ˮ�FL��S�U~������So���`�oA������9d��&�M��
�J_T����#��#���a섆S����e*�����[}�}7O���З��P��xcE�p�
��ߦ۸b+I����R���s�he����t�k�A	��c��P��:k�x���9E��g�t/����t��l��pzoT�g0������)!��m��5y�7�/<ͬK�R.�Vtf��e�w$�\�qS��k��a�fc�e8��-���+4Ğ3�� �B*������DN�I�� �X�* �v����h�_�=co�5+N͟I�$�:F7.\�jL�%���w�y;:)����N��Cy_&ldY�d����*U&:���aw�:���`�;�Dq�ČK/2W$oA�R��|�_���v�Ɨ���d�*�P� ��0Q�/\�S�C�u�� p��/U�	\�u0��f�oX{�j���&�8����Bj�fId�m?D�%�L|o&�˫�W����ϑD��+#sC5R�w��i]�e� xz/�R���v��z	x��G$�����a� ���.�q�A
��,[;��V��>g;&�%�]�u<Yn�����c�q͞�v�M��D�%�Z�BP�v"����T�aW�[d�����܃�lp�4j����S�ĽuBjږ�a� ��]�q��z���dd��u�gUV8�h���	�����譻=7��t韝y�C"'b��B���^N#Q���V�3{8��`i��DM���m�s���8좄�	�*+K��F:ί������fK�6��# Wu���^��vy-\���H�?�$����H�޶"kF����7��^wV&QO�:����5�<�N�2g�5}gE�-��� �U�7Gt�L�Λb�&6Rd�7��J�?��Vc.�}�������|��`��4ŰjA�4T�����=����=2�c�oJ���-V��s�yɡ�{��.�̶���Cl}Mj�4�b\�����"~35>P"�Y��������Y4���=~>{5yA�q׵�?<��dtu��nU������2���l���_��^���NIH�?�-u�?��@]|5��;�G�K�U��}�%U{!-uMLd�L� ��=�!��`#dx8��i�,{��-�'m����(�v����䚠ʀ��	d�\\3����/�z��i��|Z�Lz�$��J8$��,��r&ob��23��c���]b"XJF������tQ*�3o]���b����j|K�K����x5`��E�`����|�O�!�٪/���7n�v�[몾�Z���+y���hf��'[��x��O�޾Nq�Qɳy F(��y#�rz�6��������΢Ě���@*^��K�kY׽s�eб���@����`N�"��%�"��D1!>^.*�6Q��&�;��Zv^�GK�%���ǉ�G>��ӎ�������p��6���6�Q��6�Ф�	�QA�(�C�;dv���3=[�"q���Ů��N�mo���ҁ����:1E�3����5O�hV�F�ML�?tz���S���Tq��:9�ےL�"���=+-��xz俤��v�0��.ʂ�0���'�o�^z�̓������K~��B"a2��f���@f�z��C��<P�����R���G�_�B-XEJ��*�_���� J��~�Q��n}�"��b�ۋ�h�b�ֆ$|��q^5,xR��V��}��gAmb�Kn٬V@;�QB�o�V�����E��7	D�%��{�|`�(���(��U%7����_�U%kL�v/���2������(R��C��HT0;��;3C���\��ԡ2b��(v��<���;�n�O|�')?ޖ$c=��!��L�·*��?r?#���������ulW��\��V�N�,�f�q0�N}j����k)^�!;| M\��	���[]wrI����S}��b���/ȖH�I�������.����k��η�牏Vj-.�/�
�����±���K�%Ӻ&���u+�Q�b- ������>PR<u�HMo��c�O��L�Q�[��	ݝ(��ˀU��!����+�՛s�<�Ө�+���ђ#�9�X��_�9׊�K�"ˡ��6�b��vl�i��yQI�������f�T��@I�B��A�=>ο�a߹�۲N��QͯR"f��g7v�"	j���p�E�ZѮc����iԛԲ�D+������;�w�e>�7p����>Lو�#4��k��`G���ۓ*�AB�!�����J�Q)�'�>���XA{�
[.����Σ����� |�EX��28Cĵ]�����(��kR'��U�/rk��o*��*��ӻ՝��l�ˁ׉K$i�?6���^6�o�Uq�aYQ��{��Xm8kkiwh0e�O�`�e�z�N���;�r� w���U����u|���~ �f ��
�;G!�߻�F�Zj�6'+����Bc�C����+�q	���u�T�� ��s��/x)���o�C	~�Cе^����H���p�8R����2Z�k,T��垭o���*����DX������nC<��/lH�|��:c��U(�.5����������̖�S&����3�{̑�eJy�|���ߝ�g5&�L������Z(gu�<����שNu��}����{�3^v�y�;wrh�d��'���zM�F�'�Щ�ܜ緒������ß��&��e�q�Z(~�}����D�#l{?�%��1���pm�4��,թ!�����vpe������ᯏU�Ώ�3��L�t{�;�MO��GP���3�Ɍ'M5�	{Pގ���k:b�<"O�y���/�G!5R(�~�6���$���j9iv�m�["4��/��݄~�$���jT	����A0Ø.�iI���B�#
	���=q���M2���d�JK@a�����`�Y��+1)��m�������������h]�þn���g<@��TdyV�~�j֎��������+W��V=�fvm��4{���KP�d	���2h�s��YB��F��7��I�!Ԛ�{GCkݙO���ۺ^f)({$��`�~eg�8%���É�ɺ����8������m��p9���k��@���qut��r?ec��&x�,���R�o%I�$����В	C8���	�D�:�� 1��:��r�����݀�%Y�C���|������$'�*�c#j�2I)�GL��233������X����T��ĥ-�O7��ѥ���5��&�H�Q��eY�T�C�Xh�8��I[/蔥h��و� !wҸ�%&�G :�����n�*�|�+HPn��E��_W��lN���5���}jn������BJ9O�T�չa����V���eK|��1i)�_l4�H��[�%��$�=�FNM���'�{�R�cu�a���:�aX'���<�hu�TN=ג>?Ť�X���2K��z}����W;j�?p$���[5^�����06�w�1WJ��r�w�������F����O��r�1KuVjv��+��@����=qDJ��vi��,u��π�2hZ3�]�@c���L1�R
�3"�gqjg����Z1ń�[W��MVQE<�g�|dg|d��|x��� t�b�h���b��P����s���H��n	�K�4v��`�;^
�c�F��?c#�a#:���բAh�&O�F��ހ5�H�
�b��O�"��T��V�@��m�$��	�4��5��a���o������c�����rRZ�/	bGM�X��V�	g#�� �a�g@46���(���ӊ�g6&A��MA)���H����J�`3IdY��O6S�,Jnw��%�8>�+�E[��4:-��b��#��}y�_n<�8�c�>�^���VޢVf�R©b�l�����wSY�gp��F�m&��+��%3_�XzϙxRm��ِ��柮e�"�)�|�B\Ğ_�J�E�/A�T��Ա2_^������}/U�~�|?Q�T�u����HE�^�͜El�E�4=4E���-�I�3����b֥��߂uȨe`���>��K�P&Y5c�����R�� �"�%�#F[V0b1���C���H�
����G9I���,�~��GY���ÞW�i4,l؟�Q�L���B�$��ʨMa�Zq�e�&�K$	������7�JZPR�'�_�yP��.�2<��|s{]T�ӓ�w�LhW!�
���?ڏ��|��õ[ws��-?��/�J����C���҇����{���2�!P#'����b�-�5Exp���D��ۻ�龌���������_��g]0��WH���u�<p�o8�l�8h"�(*yR[ <j@m=�;�wm!���knơ��j�x.�
v<Jd!�6����ݹyQ�!^<b\�O�٧�2�Pn/ 9C�L����X�
�]�a�	.���!��I�n��I��ϞƱo�Z
GH3rɘ#��j6@4��Y���U�b�gӵg�\$�¯�Y�{���Z�'�����S�l�,F�q�O�oR	�<����Qߏe�7���q������fLx��h����FpW{��^��d�lXŃ[%mn�z¥6k��0v0�����L�#����6���C8 ����ѿD�UԤ��ѻ�17Ȱt�	��%%�ŗ�*ظAՊ�jc�_�g@ZS�m�i�-oL��v�Lծ@2��h��Ѥ;�g�����S��
o)l�al>��!��wޅ�a��tc�E?X�1����*�|inm��`4��U�ڜ� �X���ʲ9v���+������H�o�2K�2�^ʥ���l%�z��MV#�A�zS9��m�{�4�>��_"\�/iz�'��l��j��3�)x�l��~\e��\��s�"q��8�-5QQ�`_F���W1�ق3���C~��I`��T�"!#��k@�>>���ښc��h�9D��QǳcTvԞW��)��'���\?.�7p(�����Ǘ���?D/��Ut/�L8�*!u��
b�C´;	�_/�y
��iND���+��f����"0�-5S��V�e�e
2�x�����:{:k�t>62�YL�e�����@����߉(�U��R��Q+X��*��Z��t���W�L�)N=���M����:]%��u��/T�Ub2���%b@ɏ!e�ɍ+�5�Q��!~
��O�0~��g�5���=,)BI���J�(=�A���"x�/����bb��6Ӎ�+�V�*)C1�W,ե��BQ��G��l���sc �DUkK�w=�W���d���jw���*)��h"�4�M�����J�r}�t���k#��g�K�fU)B����Oc���-"���m�������W�ua�T�I"��-�ڼ�^�G�Y�����2��ix��j4.��0�)c�h��b�}|�CC��L��\����r��浛�|F�4n�a5ZR����/O�rz��l�9(��Iu�ϖ�P��Wi��Z?��L~�|��#����?y�hR� `�ð�ca�e��D��_�By�R�pxu�b�]�3��0Jd�ɹ~n|�+z�������΀�;dVƻ��IT��]�㑸��G�V���$��"����YC����\1�^9�xq;=�?����q4�ê�r�҂_� K��4q���S��3�UO<R��9����bF/�:�d<�7c�vIzEό��b�&���N ����`�~���������M�P���X~84s��
���И_X���_*o����߾�y�®�d/O�K�[q���+�]�V4j��iC3i��M�7>��צ*H�����!��]k!A�)��u�sc��s� {�=<.����K~�s�
�-R~��Q�TXh�d�.I|��u(q�H-E�8a�7�7T#��n�4a�(\%�����^����R��P��U�"�W�<%Ƴ��"_2���62���C��M)xQXY�Q^%������uצ��3��߾�gG9���Í�5()�ҍ�Y��
�S����Y�)Z��w7��8�E�
�t��3m][B���Men!L��!����e��Wԗ����?��� �u�$,�R�>7r7�P�b��%��6����&���/��C1��ՇU&�����M��K�bv���pG~e���=�E�Oi��*W1�vtP��$<�h}BX�&<#�'�f�T�f��CJf�$$�h���b�g�\� ����VA>��n��hu��"]�Ns��;�����+O��U��̴��@h�b"�Y@r��fH��ëiP��c���ǂ�h,L��<3߼�X��L1��GP�.�A�_)W��f����a(�U>x�;)4m�U�7ո�-�W���Q�����g�"���0��b��*  ����^}��GR`��(�ZfF���B3�P�فR���אO��-�M�vp%YN~�Nð?gO*�,&N��G�Q�1Z�	��MXz��� ��+K	*t �s�,	7$��b�A�Z	
����w_	7��!�=�h
�fz���Dvl���#<�F��t㩿���YM#�.��Ѽ.O�e�8��C�ݠS�=�m+�AN7�.|o�<O��V,�=ᢷ�,*rȐ�HADD�W�"/PK8LҢ1|���M���I/�_電����$�]'=k��I*[4~����)f��A�=�ظ\?�3�*�Tͪ��ft�d�I�������7� �2Lm9�2ٸ�X�$�ч�wI���������&�0躓�%�F��çѳG�T��Y@ec� yD��\*�r�+�FQ���ף��OM��8���n����o��.Ĉd�4�?�afy^\g�)vA}�J.��֛�y'&��Z���U���D��� �E�B�����_|����!N2e��ʤ�F)��㜊ʉ�y�Qg�	'�'��,�[��,"3R�3�|���FP�� �^�DL: �(g�2W��/E*�oS�E�2C|���Ze�"�~+���VL5��B{�5V"�2.��.�͑t�Y�����)�]ֻ���8��\5��V�
V�z��@"}F��w���ܷI�9�/�)�ns��3�T�թ�8�(��SkN|�3��͓�]>K��v�ҵ&CU������H�E��ri�v��x��:�:��~0HQ��Ah�BLq��־Z�W2Q(&��@�S$��}O�U��vG}��|����Hy�u�-�o�##ƌ�`�k>>�����n�^D��(�
}�YL9��0��Mr fэ���լ����_�+���zhC%��gGt�-�O/^um٤9-�J��y|-9^��C{�����U�!�����<5�]�$�ђE����$$$�J[�@tP;-�P�Q��M��}��Y%�.c��=���v����\��tt���T�`��~��Eh�|�Xƌ�b#�=�ˇ|&Vx`�֬]��"�����!�m�����ȩ2�Dy���T}��G�6�]�o������#��dw7RGG'S�c;;��ꗺ|�{*�,�S��\�Ή���:�8�˺Ka�$�N��|6�נH���ݲ�{����p�ߕ������ơ��L�S2�D0qEy����7ttu�ř�2�d�� R oz��̨Kt��^��@h}�C"T5<,��J��tdK����&��9U-��{�xI����<}G��N��i��-%�Cee��u]����p�_���F_ȹ��|�g3uN�W��XXϸ��j�䛧�d�3ܑ���R]���MU�Q�q�R����>O�ϖd����X� ����;����6_@�� ����Uu�%����'s'8J� �Ϙ2�����hJ�"u�jD����1嗢)�"j�A+[�3k�O�2�<J�?���#�yiYzU��W����cG��!V�u���a�\�tZ4�;�i�rD,��ཞ�qv9i����㟑������W��p�'�M�m>��v���	���o��SC�L�T��!����}�KjJs��U���0�C5NH����m�$� I=g�O�k��u$�+ry���U��Id-f%�|Fd���:�'�sT٤�6���A�*x @c��~��nA}��$�J�L�!&+ؚ$C�eÉ$�������;���W}�ka��&�8����I'�Mמ
$��k�=.�I^��X��4���#e;r�_�O�	��s�g�ݥ�Ѯ����a��n��,�S��3��l(87��"
h��"��p�1YՇ~5F0Ġ^���U�w���@�+Z�ᐱtsTH�❛Tb�@�p��?�j��J:��pЀmZ�5���!�{Ǉ����?��
x���n#�Q�L�ܯ?�;9R9������3�.{OGO�#e_��|�tr�}���v�zk��~>P^�pz��.��A��+���B.�����{0��f����'���6���eOv���
�;��p�4��x�-��j.��Gc�uF
�������
��8[Q<A���]�ï�G��g��Z ���īB�Z�á�?�X��9�W/z�����F7+�S�t@#-A��_9=���� �z�z]A�:qei��u!�iZ�?�m�&��\d��=�W�V>�F<VLBK�(d{��{z&J+ge��n����q��v�Zjxb"�J��q�J�Оp)_��-���eI~%�/V�˜:�n^n�`�s��6Tg�_9eb���	�/��m�)\��N�v�������'����W�E�B�-(T��.jUګ]�f�@R�����H!R�'�?��|�~�+�b��=��Zs[��@�Ma���Y� ����%����gh��Sr�f�G�̌�}���˞�FX`) ��g�Yݘ�C$�%�k$-���n�F�r6��a(㇄�~�m��቉7K?��?'g�`!�=Z�l��+[h ��NBQm�x�W�ZA��@7�"�@H��!�$���eC�T��.�W����n6�0ڜ��?�g�mUS���i�}(:-�F��G���	]���Czh����x�*�+9qi޶�a���LZ0bZc)�h�D|E�o�xMk\~+~T�Xv)x�C�	��Hb��R8<��X�4������c�ς�^��"�S����~�=ݴ�űi�%�ٳ.���󘹓�'���ܙ�BE�� �D��C�5�_*��8Hѹa����%��ѽК���%����~R�"�(�%I�I��ĭ��/�s�����G-��B��-���� �kr0���kFf;��e���U<��u�F-;v��bG���-B��l�U��ɫ!��&!�\:�p�[ �2(���	�/b%��r��Օ��~�Ͼމ�.UZ~O�Dg1�m>��1��fd��������wyO�K" ���x=�Hd��B��yY	~��}|�:j�*Cť
��?xuv#եע�9_�7uY��f��GOq�dY~��,ciб^�n���$͂/Xt���@K5����e�����o�1�32��&=gף�w�2��'͓��eH�lQ���'�ە��qv�&$��W�<5���hOE��^A���4��G���)��G?�'�)��-����<Y,�HW�.�7r��I�/��R�b���yU����˒�#p\1���	xNp���+Wz`� �H�A��E�O��q�|ON�#�WҿT���Ck<袟���$��C;������{!� u�b��x�N�?p�%/!��ʺ���6|})IHh�g�hG��~i��'V����b�۶��ݭX���R]凓� S��r�rv���i�[��������_O��VP����B�B��ə^(��/�dw�ئ8-�/,}�Y�RH�8�������"'+���!Ƕ��%mi�����j}-_J->�|=���@-�`bQ�٦P٢����`#m�%��i�`���H��5�T�I�
Q��뙥I���qJ��ES'+�dK	���v]4LP��Ε�_�A����cף�/�����H��C����,�����.B����R������z>5`bd�%H�5�SJ�}��Q+m�5���;{��8qu"̚|R搎}�6��;��*K� Z��੩1� o�,��a!$��L�Z<k����j��@�+�������'ʃ�tB�����xK�l`�g ��W�\��m;�Ӵ���)�i��k�����:���������(}D�{{bOw~��D+�E~�fn�!mz���l�}�g�"�W��sOdb��!��v��%aF� �'�U���7=�����f�����B����e��N����7����!��0%BW%�e�G��h&�
?MOv,{x{��Õw2��p��;���Vv=,n��u��6���QBG���"N��Ӳ����qS�l�	ԀХ#/��ђ���yR��v֩���G�Od3���&-�1je�Â��Ro�{MxˀӲ�2@9��t�+E	sy�^�e�ۚO�Qnu'�
{�`�	ᰂR[X��1r���v�,ТѨ�G�־�{
_�ڐ�B�7�1�v���!i����������k�b�n����a�
N6h��2�J��_qp��U�g����L�)�<L�u��6� eԛw����E�{�l���p�o�w�"��-�����Սk5j����\�&� C��9�F-un'A��W���T �X�^�hYf��+Յ��þ��
dڛߚ�v)H��T�a8���3���cz�fK*M3ຈ���2w��h6��%}�_�����oq��lԛ�� ��q"�W`�m�ӵ���$�y�TۭL�*�S�^*M�oŜ����&���b� f�����AI�^�MY��A>
E:�i\\�䷌jg����uEk&���^������n2�+]k�� ����<AK#5u�s��e'��|�(d�T�Vj���rY�4I^�����ŗ��{��R?E�?�"����;ucQ>��b}��S�`p�2S�25�*^�,K�.K�,E�.��0��6�p#�x��+�^�3��18�������A��)Q�G�������|�+f�Ĕi��}����+����8@�&pA�����)���*�e�p�_~ſ��I�L��ǲ�*3�Z�iq�z�E�â������(jX"���U�\>�Zd�@Q�5swl�"{R�a�0����enC�lT5��`�O͂��q���1Z�r��u� �����w�n�5}ǔ	U����"L��g���i��a�'AC��~�S�C�a�ץ���T��93�v�Q�U�U+��@����p����}Ħ�o:����X���'���5��
T�=*���8��0U�0E`���x?�Y����g4�*u*�[�=��n���)ý��tx�ޑ�� �}�q4�~����~'�¹u����S}��F(t�m��'�{1���G=����J���Ƌ�ۙ�b*F��������9�:e�<��z�g�O=]V N������Jd�_��+�)�@�b��ێ|P3����ɔꦪ�}��q�ZH�ؓG��پ�~�u��]։�E$[�7I3����_\H�X�˩-�����g��hX	+�~�$x���ֱ�uQ�`԰��U��b���'p��g�Rb�ba�hs��-E�=o�f����Ys��τ �q�r<�\>|��X[h���~x	��V�$M�!���<���?�E�s%e�s��ִ��	�ic�>���0���/l�%�cnE/;�k��(t��X^tg�I��8U��7:A|��������U.̤���f���l�t;ZyTOz���Pފ½҄c7���g2d,*nT�H��q�Q��Ԥc+K���J`cn�Z�8U<�D?2W~g�Ud!�ܲ�/IqMÆ�et�8�o�I{�X##~Z��B��L�`��������W��20j�=�͜�˺���ʊ�33�.!�ٞO;M���x��Oe��S�BJ"a��z޲�I&A�TA��m�fn[+��`�!�Vq��kP�yu�-�{����_�UX�J��L��"��+�~Ęq�˃g[���D�����Qa���&�WG�XML,c�u�9JO�L������K�w�� �v�K���[����O�=�z�������Q�����l���R[�;��bE��VA ���)z�R\}A8t�b�}�&�nI���J��X�D���0h!#A�����%tb+�W�<�m���z�zf>ABQ�+�	��{��+Y g��oCc��s��]�������scS�\���4i��}'1��[w�q�i��"�D
&��8b����?����B���w) ��Q�"J��p�.k���Ӯ={<8?z*&yW��f�������G+��1��X�T����荇i"��.��l��М�e�]�KrxŠ�v|�C��-Ĕ���m�:^�ǨW���{q�V7-Pv�y\p��p�5m���ȩ���"]�8}���Ȫ�i��?r�'K)1�P<tl�NI9���/��"����z�I	�I11�L�0��ޚ�=$�����%���(1E���L_�LT�>��9 z��W;�G� �o��O6е������D�JU��pm����?�����\@�?�݄����ǟ��I�%�4R'�@.s������+W�H���L��qA!7��3�X��M��2�\��C���DF��н �m.0A���r�dw�W�.o�K���)|��7C�?��BE�%�?��T�Z�ȫ{,3�vEܭ���՟�|��/LH?n�_mŚM���)?��UL|���{��{{b3��Ѽ�v'�_^�w7*���d����۵̢�#+m�ro��^��%�4�t���G�Gb���A����FUQDx�T��=��킩��Ǽ5�s
��_���g9��i�	��6h�0U�ɔ��	�TjdPZ�iǎ�M11U��U����y_m�ҏ ��G@���H�unf^�'���M6=-��t��o�� �����.�Mf�p�9
~���
ǳ�&�8RςeK`}�_�#�G��M��.U�a)ʮ�Ѓ 8�?kv�޲�
�Q;��	�v�ńJ�D����S�?6�����>�8깲���z�`���4�%��2�L�t��f����w��
`,Ə�N�sV1O�w�n��'lw9��h�������"�K�!���$��F���>sK�^8R�hB��C�<*����D�S{���r9���~�I�	�i�i_6If̱�Y���׿��t�@���"���w��N|��K@@LI^����]���,�ۚ�����p[EN�B�(A��U�,	��ʡ?q_L����������r?��p�[�~�'���b��I�*�'2+dDyq~S3�]����2r�ЦF��{խ��t�w(~�f��2[$GaU]2��ڂq����<�^>0^���K|�����p��V� ��?}����퐉�ڍlU��0�*��˰}���=�n� �mOf�st���I!ʼ�����V=(��/�p���;���^��E�~���:�t��$2L��J�O�s�3��Y��Vv^�^���a̗}
+ɛ�A�@��)[�!&!ֈˣ��=<V��/�,N]�Րe��E,�a�m�CS-�O�yi��C����7��q��Ԥa��sV��^�E�5��騼8SY:.�n��:�V�le�7\FIj���w��r���*mG�RFM�rc���Z�cF޹�d�LS}I_L����`��4�@��.m5�-��k��6�So*t��.ޕĭ�Q�3Lr�_y�t傎G�,[��Ι�ݹ������e��:\�[1���t����;M8R{#�Te9��i6<����0����m�{����)GZ~P�#�l�~q�
�*���Gݗ�ˠG����Њ���]�s���m�6"��G�a��2�&$�iTIs���-!`!��&/v�[bFMg�_X�͕k����_F:*%c#`̕�P�'�L]�v�6n�Y��<>�0~�^��s�>0��"P$��j~����(�H#�x'�yq�E�U_Lή[��٨1�W.t���q�M��Ic�'?�,S���&������;埪"i���Dzٿ����<'o@� ���C%E:�Shos98����S����ą1< ֿ����*%<a;$q��D����2��M=FD��/�&�F�;�V��_.�Թ��Ԙ� u1я���I&�A7�M�_vn��yU��t� ���p�:媽9X�[�=�Gg�G��f���!]��xU�;/];��U����#�}�SO��?���� �wJv�Lr'� �V��խ��&5T���5f۟a �7v6)((��a;�u���H�4�f/�^U�Z%�+�eA��18L{Ö�CX�����ߡC���l��P�?���L�2�Y�ip�XC#uȐ�诏�k4�rВ�N.)k9@�*�MDL.��m'�3����[��˝S � �M�x?薗��>��vFX��nn���M������RA���B��+Q)�n�Bu�t��ܽG=
[6�ӧO*���KҎ�Gw�:��'&(�������b=��m͑�-��e����	kv�OV�3wyO�26�]���|6��W��5���f@�h���-�@Zb]پ���Ţ���I㟵 �Ç�ު"��`!��D�� ������c���tm�#�-�c`4D+���[�Aw)�A�d%�u��%��k���8'E����|_��|:�s��wP��-��D-��\�A�Z|@q�N�6s[ Q�U��Z]-v��vͻ��^}�V�֡�7�r �Q�#ppJ�*���j�u��bL^Ě���äʘ�9 ���[���U������*�H�����Ӻ�D�̍�]q��3U�T@�������M�\G۹r���=��J8{���޹����	ٮ0l��
|�J�sq�b��V��
���x��(��ӡU��q����<>�8�򚏟������'8��7Y��t˧';���[e�(G0l/Rz�7RX&�]+-��}��t�b۽�^�	��F��d�p�����l�2�Hgx=Wc�,��Mx�!)q@��m2W�E�R?��e���q�	��T���i���K4l���
UTԎK$���y
󔆍�v$ڿ�fLs�2�19�^��Ö��f���g���V}��W?7����i�)x,��ޅ #�l�M)O�&�Uˇ9C���~�)�����;�Co#��
���l�W���G�i\el��{�׌���nc(��|��U��~hu*�y��e���H�0��AO6d���q�y� n�����$#	9׋Y�d����˻Y�H!F�S�m���r��3���G&��E�۷Շ�U����(���6�|�u��(I3m���.�}ܿx����ܓ�*Y(�8��Z�y�.K=�s}ļk��;�*��c=9�#x{5�[��Aj�~�R���d.�;L��e,���/x�kImX��a�����'��`��@@?�:ù8��@gg�]Ǘ��#��pl�䟃��|���=�9�ч�G���І������!W���jȥ��\�༤ay����b�F�����)WxUea��,kho�����'&�X%�4*�aO���s��.'u:���r��z.���'�N���d`_>��K�:���)���$%��\9���c�p���jr�u�?��={xGyg>=��>��;TA��JZ��^�U�e�����WL�.K�n�t�W���}KLj��q�]�~)�Ek̿��ՍW������r7>|��·��R�(�G�3�a�M}���*7aa��)u���&���P��C~﫨��c/��t��-����@��}p�:�l��}O�TU����Z��&�9�M;�"!�nϓ�+� �		Q4����f���~���j���5��(��V��O�Z{1#v4����#��NRej����5���mg�t�Vr���#\c�}|�Ӌ��K�+ᷓ�9>X��ȓ�!EB�sj��;#�%��^�ٰ�����QqDM�0w� \�� AB��\���kp� ��݃www���}�w�<_/~��U}j׮]�����x��L�P�=2;G��g��B%�x��.��Nl��<&rOfsUS��WVcm�
lJ���v
ϳ�W�q�	�@�Pߤ��9��r��X��E�y{�)�3�m5QX*&�WΡ��޳#��U�c�[�<�[A��b���c��W>�oMy��|�'�g�ql�iw�}L�k����L�ɬ��\��:vO�f��B�]&^71" .�Ĭ���Tgd+�)�LuaϲR�}P��HG�og�Y���T����IЫ7�ؒ�R�i�b	8��A�9��XU�-����K �I����/��b�����{�+ �E����I��}�I�^�����'���[��ͻ��Ϭ�|S�����K��d��~�|UŪ���)z��h$D:<<���'}h�аx��Ȩ��ԯ���hPN���}?��e_���uú#�1��
 Gs`�H�K44f��lD��돳��_������Q�{��f��#�O��i{���d��t�����xV��Sf��J�tR_ ����'�t�w��:�j͜�*�Sq�e�,�5��gd�4��@�F�nuٹ��G
&�� -qVB6'u�|p��z,-��<�&�y���*��l����:y����ӪSa�*"��s᪟���~.g��i����������C�¿� ����wߏqtX$Y�X�L�w^��I�2����XB

)z��'~������5��!1�g�VV��Q#+�f��,��2�[!=_ly�ly��s*�U���
ݍ��d_"�����=[7�5��u��I�>��M�e]�i]��*��.��ʼO(E��\���X���MGSL����!�n�~�+{g�i1g�?0�vg�%D9�LJ��;�>Ȕ���V��G��^�����u�ʂ�Ud�sy릺��`��1��͊E��ܬ�]c�%c��	K��
��V#[������v��z�į���ʊ<�:m�C�߸Y��&>{���SHte�!�&��?���T:�z?������.��|����7��~4�򍄢����;�0� j� ��r�g��\���$��U���r��@���N..��U���b��F)��#��&&/]���jfQ-�3����۰�a�$�ի�x��hI#;��B�I|E0�bT�}{�|�ޑH�f{b��f��u��c#�1x��$��j2�U1�Iu2�4%�N�7t:�y��k�`��"�Ѣ��X���3�&к����r�� �����w�&C-��Wo������SR�L�0V�����,��>��7����"���*U���;�%,�xc���,Un�e�r���(ԛ*	G�=�F�<d�c�h��bԸ�t;..�:\�!��mb][ܹ�0Ҫ��q�갆O�d��J��H%���z��ߧ�?�cwJ
�W�.6���[&x�jο�r����ܹ��:X[%l�Ϝ}͛V#a�fr����*+B�uM?��Xo�JU_��G��`I�D7+j"Q�ݵ ���Sc���K�P}V���@�r'��dg�3�!�.d��]���B��B�Dz-��;��F1�O�4P���f>��_t��"�_'�g[ت��:f�8�/u�*F�\UQ\�Y-ߞ#�{�����9%qD��%&*�㾇4�ј/���Ve������X��l��dP V݅Pc�Q�6ݴ�9Ȥˣ��"��f(+� uC��8�ps�Z�r�ۂ��N|d�/��YI1|L0����y����2�]��G���Y��+q���.�
P�	eb��"e)F���Ј'|����v��9���A�sj2�SMc�m^���Y���p|�j�h��b�ފ��n���+*4��L/S6��/��埍�@�'x�'����
4��+��o���_�s�T1��R�w�]R<�J!U���(W�!�~u�|���W����7���:00Xw�<t�z�TW*�l�
�g��}�&�L�r��i�����|��򠚊��<��yy�gE@<��!-�[��M�N+r�9U�I6�ho_�`��T�L�".	��g1��7'b�#��a��*A�aԺ'z�E�T_'L�3�io�؛�Ԟk��T������jgˠ{g��;.��5���%�w���-���NAA��_:V��]}�}�<*,4��%;�Y��!�T���?����1�D������N& V)�����z�s}��Fo��k�Cj�����:Vٜ=��O⒇���'9�6<��=}��>��|<#>lR���������?��L/7��;p��G9A�#����s>O�z����a*Y]}�hbY��d�Y�/��K��<%5uZ���):X��!�.&�e`0B��JF��?O+����VV��K?C��F�C�T�?r&Au���)E{�I�}S(�̰?�C��'�t�ak������yw�Ƈ-����i��}�0�U%u`t��)���˒]j$8Ւy�ZKl�(��9[���crPW�i���D5敳��Q��Uz�}|v@�7�}fz�`�w3V������2R��;���'�]��/����c���_���o?3��bi��Tx�+��G��� _���v�,}��&��J��nc����E�w��U��$��
4I��
����kR6ܪ+G'��*-������B��Z��h�=34�Q���7��S3�n�R��K+�YW�HD�\��8F��h��c�X�E.�K�e���t=�R����/���W��q"�M&+^^ i��8M7��d�6J����c'��7��2�7���C�Wx��[&�R�u[�j�o<���>��K�h\]��r<��h]�B��n����H����L/�̉ۂ���U�vpl'Վƙ�|�al=�b�h́: ������󩌻%C����V3�!��q`�����n�@t J^<���s6�{-t+��f�)�d�a�Q.0�m|Qz���:ҡ��q������Jܫ�
��q����a�V�@�����2���pشN���2������ۇU�-����^�@����?����=�*��쯒�Ȉ(��2����`l��,�O��i�H7�E����$�^���#{�����q��x���a@�����a%RES�pm����\�ƻ��(�2�膚��tP��]$]���Tb�њ-��:S��w�S�����<7�C�Ό�U]6��!���ո������$�,zQ�ۗ�)+uQ+s>7g����Z[�0�V"��M���S]��My��5 ���A��������xW�F�v�����"۾���Ư7"O)���--�xV� �	�k��İr�ּ�b��2�%�z��?~f�ݬ�ͬ�[�gQ_3�TI��p,�U��V�5�zˇ��F���'��7�oN��pl�%9�Cc�@2�1 C�.�;?gf�8�PI�Z�[2��q�&���l��#���0+�Q���dK���#�3�e=$*�������$��q���X	�ɖ^X��$:�1c�6��ڢ���i����N��^x�'���r����a��i���b�����oPf�ʏ,>	�Y�wc�Ie;��?f��Q�g�{��>�.\N���9|�֤]��(�`:d�5I�#܌|���$�{�ٛ.�*0	S�NQ��_e(u��Y=b��/WA�u^��-�϶��}�6�>$o���`I���W���u��j��զ �	�P�唭>�n>�/�I�(ڨ:���셍\q[亽�E]��us����%D����=G�-�(�}��dif��@��zɯ6�����g�<H&W��x���?N��쀖�t���&��O`�ٴ��,`'~�d����tw�a��J�r-.$x"d�+r6�ն{�9^&����\�ɂ(hqr2����i�O�uӶ˪m�S� [��Qɓ��C�$I�������/r'����}Q���c�|}9�I�A����݌�{L��?��*����M��f�
��2KѲ���ci���w@$:�?���t�O14Ȧ)�$+V|U��C�q��ĈK!f+gˮ�����S�L3_ݫ�+j���"�D�\�`�y�6ߩ�,U8N?>�����w�=(e�h��k���<�{�H�nZ�?��ڐ��Yo� 0XN/'-r�K;u
�&���dA�Z��.�V(����0Y�L@˒���tVI�������6_�/V���sۼL��H��R.��gyy�el�\����;@-=�M�Yȟޯ�;4�*�a~��H��]�'�|}BR�a7�?j�}�Uh�;��۸p%Ei	���6���ќ�!0?z#��[�)G3q�� ����)���^��U;����{���5H\a��)��ڂ�x! �dcB>**:�Հ_�t�'E�AA��,FJ�.���ϚN z2U��Z��(Q��3B��AhNIj�y@��LO��Q����|�Z�����9i��� 6@�7��NR;43��	q�Z�O� ����&[x�)C1]=s�n��|�����ڱ���O��\5�4�R&�k�<eVq�N`e��A9�;�4u'��
������bi����|dw�	���O�]R��䰌���YN��Њ�y��6�6^a`�_t,U�<�h:z�p��!~�,�`ѣ��X���DP�\k�e}�D{ =88f�ۃ䩮�����iӥ����|�%�k����.�I���ls�W�/����&'�%����Ebha�`\5�������VF��`�/u��	9A�3=V,䜫�(��F�S=��Ut�dz�V��q^��9�o�y��A��OQF�y��F������bsvɸO5��\��
��Z8g�r[���g�c>�"iU+6���Wr+LY�42+O0����H*�m�e�	�=+a�t�T���p.>��R��r\"��*r��pJW�.k�*C���VQ�l�j:��D�����'v�b���7/��8˙4�X �	'�`m}f�)����t�q����k�������ۻ��pi�'��K�Η!j=��Ob|T�ye�'˽����}�e�ع�sQ���:�ᦡ��������oǶR �Z��WM;��$z�j|��/�O��������M��g�z�L~�����O�A;�,�Z9�V�v�ʅ���ɫ����0�u�j͎L ½Uy ��ԭ�;��n�fZZ������6a6V��F�<w]E������d���1��V�_!�@O;*��jϱ�� (j������ܼ��̒����T��_핞�vt�a��Nsޙ�q79.Ҩz���~����M'K?N�"��]�ՠ��i�E�>���g5�_��^/qv�-�&}�~�B�$(����(=�INS�N�#1�G>�4� ���'.�����'��c.�A����V�`(r,�صU��
�{��#��6L0�Y0�l_*1�� �t��ҽ�"�@��M/��%<��2,��R[�Xid�3|QD���}-��S1�{d�����|��bQ�6> �Qs���v�,��G����#�
!am��Ǧ������+u D��F�1A�`�1SCّf.i,A�?;Ց�B��=����������H����aA�O�}*���n���}ff\�0��F���:͐��5�x���&��J00�*_o7��m�P�>ӱ E���8#�
+Qn��,�{��?u>ܥ'�B�E/D�wБ��J�N�}W����aެ�bD-D0�	oI������hՍ����X���ƬV��y�B���R��V�3�|��XO~�4r˥Ǉhj4��i��M�ңIǜ��^�&~�w�X\��jx:�����7NP����@z���jr��L������5aM�0�#���­�[�TE��0wo���N͘��̢�8���B�?|h�˛$����,����l�E�FZ�h@>(��>�]n�*@��쒓S�����Ø�}��~�Jٰ�<���e��s�KM�P�d׌�=y5�QW_3�=v���?c�b~A���T��$֩��	�ۚ�[m���-P��0wr_���vf��5��ws���Ԟ�*[��7�,W".CU�:j���r��#A+���_����W�+�,�i�b���yyS��ߏ�g�m�#~QB�����
��(�@��h���Gể
�|&@��	����l�m��+k�9���� xY�gY�������8㏱���q�_����|���T���z�{�B�w�wj�~�x�Yf����.�/q�s��X�`�,r����8���zb��p�qErƵU0���K�Z��|��������a2Y�2����h., 4(���T@�[��3�$�����Mf����|ƿ��ؤ��q��R���2�'b�+����>)T)Y���U+SRW��5D����%}������� ��T�rPn!u_T	)��1)Ij���b�=���{���?!��Y*Y&H ;T�U/>�L����17u�^"�!��7&Z�3<�0�h��n0�`��<�-O'��$���M��Cϖ=b����oJ<,�׬�v?�E~���(c���񭄊���h�ܤS���xw{>t
D����5/��:�0p�	VVu%���P�B���b(6<�F#cQ��G0��F%���X>'���`��u�^4�fl�G;MHWr^o w׉{SV�h|���+(�r{�`��X~���Ͼ���WCe����o"&.ٝr�%k�yd�#��ݔ��O�۳�-�X�AG����򮅬��]�AD����U�+��	�o�f��qdU�[�c�c?��dֶ����Z�C�@��ڪ��=�=)Y-�@)I����������O-����A8�y����v������6��`2��lN55���*��gۺ��2|�p���oJ���~VԼ��DC�}�4�h�z�S�kz�KkC{����P����rK'w��k�8��H�C�[�T�Z���30��������N��"��U�Ye����C`V^�����{%���Q���xg�r���W_��?���T��(�cS���
)+)RD�������5Ξ�+��9i��Ѻ��S���G)�'���
�q��r��q� a�`���r\r "��=�`̏��N���vd553�]T��_}[�D3���&�������&(!�a������\�Ыst�H��@�7��&$�{�F��0�Y�q�Wz�f�%��9�	{�mR��i��6�0C��OS��<����ߡ�81]!�_����V�r`h��ʭJR����D���*S��mGv��t>�fN4�b�v�9�B ��XS�B�ˎI*������[��DP��޶(�����3�Z0�֭'ƻ5�|q�����кD��qx�"�a\�!��Y~�yw�y�;˱>�·�����/;"	:��?�q�����16D���W�7;�}*��.���=<T���.�"H�l�o���DHD&A�ݪݤ�yf;6�}�_fp�e���+���i�8U�>����(2�Or�81�b��OL�%Wo^r���mR�D }��Ǫ!�^��uM�آ�	��2���S�x������N���Ch���P��o�%�[�����Uf�9��{g�>�b6�����olb�o�M��m(Y�Å��W=�͓]b��h��ɐ��/`���Kũ�9*��(�!;DN3k=�X	2�|��'�.F����yВ���M�>KK�n�,.t�
9v�4����B�tQj5$�U�$�[ywB��h�~�����������dƲB_&:���Zơ$�OY�H�I��XJ�M����%&;��E�\M˰N@������FO���wӛ�C�޿�iRv�Z�
��j��{�X��c�"��d�Z�s��L��H5����%�����cX�Y�k����>�J{Y�9^�t�`sf4���{�_�Ǎ�[�{$z����Ӷc����bXB�*O��@r��ݔ"q�r`b�)�5rљ�$�>�����)#L���#}�����o�p�Km����"g�I+�����o�sia��~��������v`�NO���m����nՐ�N�M��+/����G�'������=^&@ۃ��`6'����
ؖ'<k� �Ҽg쌵k	FFΛm����b	���;��pI�7�8�z�3b׷��d��5����O�=�������Fb��!Ƈ����/����������,�ļ�Ր��ܿ�?����sz\(-�+��������b �w_ �:��J�ɘ֢�R�V�5Rf���*z����{Ǉ�Gw��ώ�i�;��A.�"9���={�J��R7�������^����h0���csQڣJ�Ɵ�I�����f�S�l���cbn��a�������v��ب�(֍2�����=)���ges���sZ��7�������h���*���m�E=�x����?�ZJ������>ҴH�)�$��d��	�7ņ�[�����_�5�CS��zxY�������4�K�W�v�\KU`]81�T�m^0�� �Z�T������Xe�=e -5��_m�o?��+�X�d�a���ߴ�h�T<�?:$�����eƩ���;<��z0	VX &̭� ����I�Q9ȿY�8ű7-~�--�ҌSa����@�������c��+��_�����L��pOqw� m��g����V�2��w`���4�7��~���L܍cZ"�e��U�l�}:��_���M��VS���K�Y��A��ٿ�4R_�o抔���qH9�_u��/���Y��+Vy:���c�-�؆��.MTa�zg��h��g�W���a�z�e�[�4~Os�Z���K��pš�'�\��B*x�\�w�8��B��j3K���e�48u�y�@Q�!����rDD�,�t��]�;d)
�I��M�̠|��?�h�{7tc�ɑ��<7O��_eB����79���w�!�փ0�dL�̥�Nb�"]�2]�#�u���X5�:�G���̴Eg�d�a���jQ����I.��8D���ּyEї=N�Qu�0w�GT@%��n�P)Ũ��z�&LM�4�?5-nJ��0;�Nl�1��������TX�>h�k33�aW�h`�V1�_Z-5	��F�1>�"Kf#�U��y�>g�g�p �e݊�Lo��f�j�(�����<��=h�z��j�{�u7(��`��ғG6�����_�S�@��@nq��*(*�j+"G���,-%$���D��_����\�N���)}�خ#=8f�m!��*I��������N�_���%K齄����WA��ʹ?��{�C�TW[_ �@�dwߕ�s���w��c�^�Pd�v��՜y��e^/+���	
Y�kOԷ����Y��LR4t}�z��kw�r���8C���l�J���u���3��Z��}��D&6V�����L����-'�Ƚ��ވ��ő�EI��)�"6�`V���'ќt;�l��^_W�l���n��t��vg1>��\ޖq��&A�qm�����-��]���l�ZM��ԗ�EFɚ����e��m�n[�,�`v��1�a}qӄ��y�77Uc)���M�JU��3��.�ы�5�p�x5f����Kw�6��ֿ
J�(�2�,iܿ!�;A�H_��f��6]�8�.������ �ܔ	X�����}f'���s_)���+�7��m��s&�&e\g7�#~=>NJJ�F#C)�A��LUy�G*�Ƚ��ѭӚn
鷻s�~�zK������^%E4���?� |��Pb�3�I1�۱��jz-)r04�<��>��=+�������.�[ot���
�ݖS\����vص����2���|����*���	��do"C}���(���HJ��������_�z���%��9�:v������X���-��H�0I1�p4z���׵��kI(��]D>��Q�3��4y�>y�*�!��-���H8��2�0�?C�ݠ�+
>�����CE%m?Z�{��z?к ��ܮ���g}9�w���3��Z��5׉wYee�{���>�RE�޼8q���q��7�w��>�ۏ�;4�^�RGI�3-��9#*ю�=�V����o����^4�d1v9#�w'}k�DJm���m:_	�,���A�����.�K�P��g�E;aD����p.���Ƨ_�/����&'򔂔���icJd�ɜ�#�Z�Ԗ�R-�t'hV���u,A��\� �~ ���Pd7X�����]���]\!����T���;�^A��z����v�W/�顊�����W�����,�EAV�;V��*R]}���������ˠIX��oR�|�5v�R�m*K�d!sa�_�0q�@I�`n��/�NT{�|CՔ�;t���UoI
ۮ6��9j���j� /\�R뙕o�9'��·=Qd�Qd�y
 ��Hjks���EΫ>��B�x����p Y��*����7�d�qn.t���0}e�eK(���3kO�MݍD��
i4�{^P�����1i��zm�Se����+���P�Vk)�Md��PL��hlX��g&��x��Z`�-���Vnt���]���mB�;�l��`_�����E:�PiP�*��]�&�[��+2�k褤��M�D�6=xB�;`��}5J����8��c`�1%��k��#���с�J~��I��*gX&���(˄��D��_��a�/�t�������/e���e�z�M��"+���8�=�$��+��j���Z�s�0��j�� �h�-?�x�%T�r�L����΀���1*�LRDH��0��ԇ�s�r�wa��)�:v�Ё]B���"14�=������筠�pTv�pL�2a�B&�/�"���]�yi��������Ĩ��)?/�b�Ri�nY�Y^��� ܻ��l��J�`�a�	��K��gv�aZ�J!r6azݳ�OhDD0J;maVK��t'�>�<fq����c���S�p��,��qViIF��2-Wɥ�"哢��q~�����Ĳ0[�(|� �T�ىmQH��E�:�S�@!�ޢ��E	<^8?)��A������I�0�0md��O�'/�; u6�n��J|}�A�E��5r��M���K����pj��s���2�>�[�]K�Q/.k����,T)���qw��h9��ƾ���\a!H0���w�32��$n4�g�&e*-y7�'��@����A�z �4�[�A�8yr���
"�������S�+3��_cD��� Q)6�a�Oc%l(���_��iF���KW
d:�������A��� ���F0���^�AF`c�����ջ���8Ǣ�j(���E�(��`P0``@�����b��{�ڗ��x���ǖ%�ԉ���(�D���_*��E1F8_/Z�[v ?�m�,���͡�����R�
�s  }=2o�t��݅�6U@x��(U����~��qV� < �������ÃM�d?��,~M&��p����I�ۂ��5` .�[������+ �*��M݊x��8&<c��=f�]�կ�b�����)ۑ5��2�h��J}�d`v$��&�:qQ��Q��\	��ʖ/��BV�]�R�e=H䯝��R��(�(�_�R��qgtx�St�2�ɻ�>������h�<O�&� �}2ϛ���]��S5�8���S�=�����bZ#GZw�[OK���,�L^=��"@�����)[�5��:<2�����c�������4zs �d�g�yv���9AFZ?R-w
�8��pG^ё��}�(�x�5�#b]F�_m<����(h�}
��(�����r��lڏ<��s7�ot��/����4�~d"�Gb0(��W�K��J�I��L$�_n-�����m˓���2�M|�4l�����P���}&W@�9��X��^�jX˒��V�ß�_緞����^z��Ij\d�G����It��E�rDb������C���K1�(z)l)��:H�HLJ�j��VtR�p�ʃ?����ty�l3�@UG��Εi��;�h��/슐�6칊�?�BVcB���њrh�����،�Vq/2�������_I�bM˺$�Cz�E:���=�?��ő�p�kM�
*�,З~�-�sa��.cv�:򑅆�F�-K�1�MMh�W�������щ�C*��lС6��q�K��.�r��$$�$\�(��:�0|/?Ϛq�����q��8}�	���8�T,���^����+V�JwD�������iE��N};,vvvlg��!�CR��͐v��Q+����ε��4f[;�V���/F&|�t ��:�d��"��ϧ�(�������<,-YR�9!�y���8�;����~�A���!qK3^�N8����F�E��@�R�!�|�;��Y8ܥ���/Xv<���
���V���Xn',qLz��6��s�\�8/Y �Ue��f���1z��/S:�mr$b7�%7K�O�b^N���+d��ʹ�`�".!�#��Є��Ɉ/���D^/&��_����3�h+N���H~��4�]pph���-�6=����:�Q�� ` Tl��BG���q7#�z"�G��̥���[V̯�P���T+Oӿc��cP��`�EH�������a�d(��㞭+�����=yoU���������$"S���%*��#�#�w�&���{ڹ�-�@�@�02���N�������Z���a���ז�^̱�\]}�s
������_�z,Us1((���� _8dz$#KQ�L�?����q8t5tk�I�O����lcG�<!�oz����0U�Y�9��7��cր�]�p}�9_ϔ���[*�ohA/�Fj�}w�9��k�[s8 ށj�u���a9�22�[�`�&&oA��W:,�9��.���j��#v2h�����V��e
�G�H[x��P����(H����d*�陘dz:�S<�(jm�:��
���Q�i)!%��-�	����Xy^��T����m-��o�T���F�.�όU�/?ͩ/[��{����q���(����l?�3�Tl@����'���������#�.�F:i���/��,<�)���zQy���g����gU�Y]����[����Bs�S�Q�����x
*d�/j�a�?��:�Aܴ�id.��	��٠��m�Kj�^�\��k��F��QAs���b��S������3^0�;m���rw��M��"���L�&��:bI��9��m��sr�7��z��'gQ�ez�ͅR���痓�֝a���N�D(�t�����Hg�@����*��X�_��;ܻ�8��^�Dֈ0��e'̠��#3q)RI)SS��E߰�9g'��ҩ��5���+�l�a�l�U�C��{
窎@��� ���oGG'ʟc�����Ŀ��>�q�_]�Ec�5�����G�F��~�ֿa%1uA���Q��t���&+������r������|vC!�	��[,�Y�=u�B���B-�v-���ಐ��{G�7|�K!��?
�<��k��#��nb���jIY�]z�R�Q�4Cp��i78� +۴��3J�0�?w�<_�=���t�
�m�'�Sf�L�-�g�<��M�k��0��1�}?��,k�+'��v��gc�>"�m^�;>��&�A\\��kk�5B2g��h��pr���AK��o�޽9 %s���(C۽g\9����2y�!C}an�>k���,��C2����iw?/ƇqO���r
���t��8��@~�ݼn`IW~���5u!���Wr{2Հ>7�}���`5 ��>ЄF�1�<���7���njjf<�����&��_�l-���S@�4`t� M�V��ZZ�¬�=�F���SqvTn�����n���Ke�'�_<�CX�
�RQs�خ����� :��C��+���=o1=�ί�JO��=�g2�05QLnp��nEn�7��W�<d�� �\��V�/���q���ǧ%���g����C�d�y���~�
�e��%���cg�y15w�r�w�/cȾ�����6Ed"����BM�Lˏ��+�0�<�]Y����c�1'��xC�ǣ��n�Yq�\>A��q��>p��ed���$_�!���G�q��'/w��,Ys�|��qoqe~� ܐ?�k�x�Q�����e�Y?�X�My��{{��QS`��<�L\�c ;"()�?I?uݕ)������-P���u	��4�b
�b���N�\���G8����sW�� �����eG��NC��t�MC��@���y���?�Y���zb���M�v�]k�h����4���9�G�0ֳ螑��T��~6�,��
=�p�-��=��ܬQ�񼅶<[[���،bh-Ȼ7/�{u�:�6��k�t�6�7�i����Ub	މ�ޗ�x݌��ا��ί��W�w�lz:���t�?�I� ?)mr�UL0��^I��wN�M�@���K"Ӵ��2[�較�/�A���9��R����W�o���1�Δ��
|2u��P�(�`�WMw�Y�dd9�?P�.�1=�\l/=�̴���b��D�_�m|���' S�]*�f0�6X9a��R*\��#X���1f������`�~s�S�G�"�79�v��l�?�y����'�}2�p���D1)�z���){d��Ў���N%?�=�ά�ќݢ�"O�5!O��H��0�H�����Q�X��W��mظx��ǎ���k�.>����������D̯Ã��ih���a<����uͰ���GqTe����v��u�&��ceߡMcZ���<%[���u��n���}��7��!$)�@����eT�x/|�Q.t6��y3NW~j� }=^}�v�vR����"�@&|uu�L��y3 3i�Zs�B�=�ܛ�&�[��>_�64w[������-d�a��vc�g�H��Z�tEE���R����K�/H�bzҒ7��q�]�6s�co㪠}]O�D��,q^u�ǖU�B���23���4�`�9i�aocQ-1>~��2�i�tQdF�����/J� �|_H����֓���-�FO�K�زJ[����UA	Eִk�C�WS��ϲ_M�p�1�r�sG�����$�5B]��/;�m�q�B�_�~i3N=8煔�3��!��,eh[x����b��9�4��n�DAW�s�W�=���4����S���S�����5���)��K��6Uv��۪�鬳�ͭ׳g����s����z�p����G
�G��,��D�����)ΰ�J'�X��Q�6=W�(Nf��*}�H�ćr|�3�?-�?��?��Q&]K]�����wR5�Դrm�d{���ڍ~���yơ��[7)�Hu�{��-9 ���oZ���%��7u��/Q�˩��o�FfӘʘN�㦫-�m��3^ ��+�:��=�TH��̹�+ ��������i�4����Ǆ�	5,+)۸%@_�]�â�ć��ӅMw-tf9Z�5?��g�PU�E]��fG�
�2��*��E>�2jARk_'�۶\���l�=Qd�X�$�g/�6{S����W��:��r0:���!�i��N���tG�^�Ս����`�P����N).7�	Z �y�l���g@!F��*��o���Tc�Q������*kZ�\I�*���(��#�z���=��+;E῿n�H/ۿ�&1Oy�C���/�Յ~��U
LZfAmK���LJ�r#�m��4����>�q׉B?m�𛄄�ctCq|��J���D�`M��Iz��V�0�/UU� ���ͦ���Q]mz���0Y�1���;(n�����u}��yp��N�&~M��5�U���� ��Qh���p36���!!��4����WY��������e��:�����`�3
tO��U���T��w�?�9,�w��~q{bEo?�L؍�j8�3N��U�j�D��!t���$L��׶���yR�j��2��������Do�t��1)�dbe+�q��v1ۂ������ji)$ؽ��cII�Yo`iIy����IE���kE�7��}z�z~\{_��P���6�Ą����0�_����a�w
>�,��[1�i߾��Hf�bC���N4�f3��m	�� ��֧h;��fO�U����M2�,;��-�	ܰ�G�D��)�qԩ�G3�L��;�mp�H�����J�c-uM>�{��l}#W��,#�����x<�wt�-U�Y�����4�1�g�ɧ�ͻ�����-���끫%_Uz^gg�j��%O�����]s:��.�S���	����׈�+�!a�ja���]#�-����e�i�I��=�u��T�n�k}�`5�(U��5�(�9F��gk�Z8�ꪅ#�p�ov�;8�j��� ��>nqä�~�IQ�Ϛc�G��PG�w�Ŷ�p�0��Tp�h��J6��eh�>�z6�o�5�7=B���ϕ\��iT���!���J�l���9+�Bܾ8G��H�c��i<TtT[9i&cv"�ԏ��s���@t������Xn���O�p�vq�ui��^�[�Z��{�,��C���-&�q2�4�[(�=�@� Dq��>��9���-��zf��?;��bx�N�BVm��	H��/�gU+��3KOD��Oa��h�r�\�92����="h�/VT���E
�l�<�����,�Vz��QC���M�t��ovFT>��D��xq̽�p0BGIU?_o��D��:�a�r��0���m}�+S8xHρl�N�~,05�@M�)X�d��lqk/�,ޥt�.)����T�x
E�qZ ����������G��5��x9�+����]3NbK�Mz������?�?�'|��V����p5]&�-�÷�!�}9❗.4Ρ�9�b�c�bD:�J�i�r�ʄD�"����SG���Ky���Y_�t;����C���5xpw��� 8! x���Bpw��^s����^n���CwU�]�vu�ӓ>������ל��n�EJ�X�N�/��������̛�P�8T�1K,�8k$�/C'.NB�D���T�
<�3����xo�@Z�� ӥD��gMt�y�%Byy���s��V�F�t����\0_���[֌����5��Cd���*���Z�k5L۾k�N��E��7�{� �{��oZ!�|� ��������_O���M�M���a���<��;��%Zb���*X�>;.Yp��8 bH���̮���%؁} ������J�Y,_�5w�AB��%eƚ�/��r�bF1�"Fo�b��8y�BE[����R�����lĊ �͔�=�oI��E��K����~y��`�))3al�������q-�#���i>����{�p޼X��椔d2L%Yr�aBV��Qz�h�ɹ�s�:m�@(/�_���W&�A����%���y��}K�ʾ;h�{ϔ��)FZ�[��˴A딷�bKM�ʸj��6S�:>�8f>�J'�P�q�6����U̵����ǥ {İq�ص�4�_�:g�s����$n����<�N�vP���G7���7���d*J&�ν�|�%��������r�r�� X*)���of)�&�E"-�˼���h_�i_�hO�&n�u+6E��R�q��4�kk��`�����	�?v�|���t�5� a�G�U�}�(P��}�+8R��6�P�:��i��'!J���MiS�r����:�U�ûI�Ϛk'3��yc#�n��O-8B�.�๊����0�����ŕ|+Q�J ����g�Zx�ذ�{�t�Ȑ�y";>�1k�H�>�8*\Vd��|�}�+����U�Q�|�v�|���j�[���{<�}A�:Uv�:7Z!�ΧB{7��@5an-���)������p�'q�;������(�j�n'�>u�2�O��h�#JO���QË��x�Jd3z����&���eZ���8����u���
�t�o �N��^���Z�XNw|�r }��LY�c�˅¶Y���^�zI/�C#���o��YZ\�3_�Y�j��Sld$�zǚz����㰶�.9�ұS��@��{�b/UiR�`e��O�Uɘ���=�]%}�]�H7�2/�I*U�4����a�m���w�ƇL�,P�ۏ��gO�����x�teR���իG�wZ��ņ+����m+�T�[��5�kw�(Y$+�B��Hh�����3�"P�q����9!�ƨ���}�S��Y-��f��ʣݫֵ�9�A#�������.�D�':�SO��0*��4bd`�_1�Ll@<��iG���Pg�b)�����r�o�/�˦g�^��Rci��ѣ##X�q
*>��{>��R	Vo�anH+�v�[�f!�;V?��#���#y����mp`�Z@�\]-325N�z���Ի��#��J3d��M���O^����7�ٻ���~X0�|�$ %'����;U�v>�6K�hR��5JB�`u�h��nl݌�/ ҕ���q+�U+�<O������
�c�+���F�g VPv�����\4c?�����6�x_��m]ᐭ?�[�C�>�Z�?�4e'�*��x�рUj��b���;g?�c=��Q������'��H
pլ�`3���Z���w��]��럁G
�q���Ps�ct�Q�3��y�tn��o���Lg��\���<�<����_	Gq*!�X!����ԯ-ɟw��,szK�w\:���㨁��N���)����J��ٿ�<����u�0�6��n�$����	 �T*�+�i������ E��J�h2@6�Ue���ڹ����w%3��\{5�9��m!\٭�u�G���J4�@�m�gB�F/�f���z�`S�Dˇ����\�m����p�:;��T���*�m��JvMGΝ�Z�n�z����s�k$F+%*��%�+�;giD��5�ʙ��^�ŖR�2��|E~�C�zX��RWS҅����c������:bu4-��T7�M��nڻ�X��B�� f�g�`G^Xo3~�U~�[:��+~m�@y9׉�SMr�����7u�v'�<��Uޏ��[�۳��w�<��x������0���;_��x�?���yw�a�E���F�gXWA�o�,�|eɂ���ʩ+���f�� �Ry�(~�R�p(U��zXE;*��>h�=�� �ih����OV:Z��Ƀ`l���R"��%k��ˌ��'���8���/��^�`"dd"�Y��M;u��)!��c�0-Q�#?c������ĨL�ׇщA�lR1]ti	.�Q�:�%�*{Yc@���NT� �%�.����n���ˬ�l#.G�
�N�ɚB��wc��*�hփ}#�B����?5��zDF	��$���2&�r�v��T�{,�y�TF�y
�C���Ă�2�� �i��tߵ\II9M;4��P�z5�4Qv��/���̻u��Ϯ�=�Ɯ����.����J��s���p8������UpP��2����)��w*C�e�f�In��2�t@�؎������}Fօ��a�ó!M��
�Y��?�?ʛ���V��_K�t������`��}�g��Lu)Ɠ0�>�'�I#�e�z�X��Bh:dq�c��x9��̼51��f|c�՟�lĪ˸o_�z�C�ӈ	�J�	���xI�d���-�}}�[F��8�"l��h���{����-�"�C�ٷ�H��b��z`�F��6�� �s� W�o�9�IZe�/�)��9�������@ ����Ug<ť�뽜��h�_U�YJtJ��ל@g�����t�����Dn��S;o��f�+�%��]q��9 ��=�Ex�]�s&\�O�+�`	��3�x	�x7�8���R� 4�{6b�{#�s�R����E�Ҏ�Q	NZ�]��#��8=�5�k�V���Q8�%��P����A�Q	GJ@�w"�q�I��Dr���--Z����L�ʕ@�]����i�,jHP��1��ӧ�*xc.Ƽ�q{�������>�S#���Q��:�pԣj��##��N�}�8�JA�MA��N���ZsX:E�Gs���U6S���0<�<�hLlZ|e`�%9�m�t�
:�4�Ӏ�T�:3�3�Be�D�]�=��[N}봒>�{���*��kv��@�q !�x�m�-�,�쫓ۀ�z8��B��1/!�jC\q����߸�>�� ��X[w~r)�<��l������`R-��0�U��"��G�m!󳼰�hl���
��t���b��b��b�2����,��f*U�i�L��i>�s��2D�v�ҍh��{yKI�'/�}Nl��>C��Z�?�".�_vJu��A�?�u�PE�}�
7���xgzd*u,g�I!t[���3�=�{��⟬B���j�11H_��l�$�Ҩ*!R`���&(8��y�S��(_�B�L���o�e|�;*,I˄�a��i��`,�x�x_hA��+�gZ���G�F���1%�r��������̓@L?>�g�$3��z5��E��%	.�Y��|��xH�TM�i���z_��@�-�q��N�(*��� �MI�`?ꠅZ��=����X���&�p�Ї�	s�;��e�;'_����:�츏�wo�FӖ�����tl'3Pd#*]&�}9����*15%�T�Hfu�^�DƅeӚԫE��R~�&��h��$�
�$m^�wk;�������)��od�a�Z]�2e�Ӭ�
T��/��\�Pᴠ��,?�0й��jx/m�ɫ&c��bo��<)���[���p1<](|'l���x��X9r��eT"֟r����FS+�a��P�pjaKn�����%����nd���*���O����ȳ?�(�I��-�7�꙼?���&A:��J7{<��) ��_�b�u^u���؜K.9�x��������êуo,t^�d����2)�����=YȒ�lj�Y�>�W>
��� �e�AEK�\���t��$3��VeI=�'a*�.��X�Gs=H�,�\�*H��=T������ �|��tƫ�n��@lZO����>���Of�b��.�
K�5��r�f�a�+�2PA�����,_X`[��g�� 5dC�털"�a��}5u9)���������u�Tbu���l���E�^Yj��Ckl=������$o��z�'�]�*�`4�{-mè%vc%��&���w�0#�׀����I��n��f鸍��+ܨH5F\\���̎[xǪ�&G����%�nZ:m|	q��gZ���~��j�J�Ԏ�;g���Y��)��{�a-X��A�����V�`ߪ�>;x C��Y]���>[���U�a�%��M�T��emĳ�l�Kޟ���h[$i\� GW7�M��(ڜ��E���S���_lK�f����^�{�9(ĹSCm�W�8�тĴk*�����_WVB�uˌ�{T�'�
����f=��w�B�;;s%w�!��Ӧ쑳���3�[�~wb��{+@Q|����p*����d�49��E�4�yx:����Z�*"��`��dv�Qe���b�9k�td���\�IM�6��������t"�Px�1���9(��e�4�̟�(*g�+;.�;`G���l��V���nʝ=�}ϵD0#��zu�HW��a���C a��eC
��3�*!L7Ny�
e>
R��B�nF�T��[Ǟ��{Qj��*1��;|;籂Y9�v%S���?r��q�e��Y�����w�̬R��0l,��F :���&����0P��ibfc��$o�s��leV6����%7�ӥ�*�{A��P	ԃ%>/�t :���v���P�[��G�����$$0�G��Z�xFM$��km��ב�a5/K��$n�q���l��U�S*Ț�q��匮���a��g�*�V�0����������֚�a�Ǐ��^ ��n�0��Z�� ����Q1Y �U�B!������͊�dH�������ڮ@�2rp�-q_8���\�y�9�~/*�/*V:����uqֳN�K�_z�m;�l�A1�؊�lP��i�c�vE��W�������2K�_�S���S1��<��r�.�	 .���g�X�z��Y�
�5�H	~m&2
��]z�d�9J)Y]ќ���U�;���Q=�Q��_�cn�@FG�ȿ���7s�!�|����w�o����/�2#�h�_?�������]�-�H)ɢ��'p�vw���u�p��0�a	vHO�,��Z]ΐ{�;6܆�f�~�q��紡#��F�$�-��w�٫����}��^d��5m������fTI�07���szw�����[8�� 0��6�!�A��8^���9Է�ɋ�<�TA�*Us$��H��{c"y9�!Zv�S�3����I��ؒF
�6��q��d�����ն��n��O�c��\�In�˦��}��JG>�X��ܺ^?"%i��l$.�Ȩ�����ɿ��C�M\��Z�bÀ�B���|�a �ϣ�a�7�EU�R޼����Ux������E�*���'�h�<��"Ӕqu8_u瞴9�_G�_wfʬ0��?o:�$#�����e`��JϷ�hBR,��C �f�l��;��RBK�؅7/f߲�m��+B���ͧ�2d��^�HJ5�R9�&s.}B�'��tK:���9�x�@k����Qi�.�<<��R�O&�&��I\���p���e��;)��,$��m�1����?��N�7��£V�������ϫ��������@�t�;e^����-��W]�L���#�wE��2�e*���2�k��O��n��p�M�I�/-5�������9����ܿf[��)�S�J|I좔�"�����I5$&��G H�nD�}3T���c΅d4�͏O �/e�$������[�`���k��ԻU�U��RRJ�:����2�A}�������\A"��É+�0�wO`N��5N�#u����,h�K��6à��<�M!ϥ�����Q���n�M#
�+���q+����)��a�:�O_�)�y#����	s�2�]&�=h	�OA�s�[�B/?�1��GhMcgm�O��}��������U�6���$�	<��[Ԑ̸̽��U��@J$\���]A�������Qz��j�f�z�w�:#�DI(@X�W3�Ua����>j�^�Y0�`S�@��������p`WHiR�%�#
{�4����-���7�x�"��F�����o�|�w~�7O��D�h��x����k<����VJE�m������Ω���2ӼD�p��E�A�,.ab��}ٔ�~�&<��V{�H��	�CM2��x话C��32?��3j���e�ڮ�Dn��>oI�DSz��k��(�\h�k�𴞥{�J�DU�R� �ap��5�Bii�^�-j��x3g��XuK��*4k8s��M)���3#;}:��Ƙ��:�`�cI6��:�8/��#��f�n�R
7W��d�n��྅�KYą�8~�84������j_��-����ý֋�/�݄tӪ-�04�_���/��М��N>�O�@�7�%&�!��%X����_�z�ʊB�z|jfe��构4ڸ���z�#������q2y@7W%��V��8~���pF��Z��'vl7�O��x���J��DȻwY��[��|)����0�\�5����7������L!'�䥁�33'���W~���ɋ�S��zߋ&���Z�M|�9�T��N�d�u��k��ꊝa��ӹsZ4�����4�>���#��/��u�7����\xg�]�A�o���R��%"鮥%b�_eL�N�\����뽜�����\B"G�Q��8�;�5Y�M�z5����B �K��/�7mT��{]r ����q�b�
�R�I�]3W��r�Oc;p)�v��A`U��$s���q#�Rf;�*RΌ^��,��y~4� }��@���w[�������(�o��Cf���W�%m����:���z����*V��l��G�r�'Ƹ�Zr=��^y�����fÅJ�U�S��nR��#g��^��T���
�i>�ny�ɒ�r �1ݱ/�|@�L�1����j���AX8nF֧�<f���93.ka��<�'? !|�u�I2#'3�w�sA�^�����! ���8�D�L8m��40�0����u=���g�����M�r6�Q��g=@�r�!��Ɋ�PPcf�S>&!YLԓ2�?�A������a[t��V�,����ˋU[�����#i�����T-��3 TSf����HD(�C�rh� x��y�h���@p"�W}�7k�깳)��D��8��8�0����.w�Q^M$�Q���j�K���ӳ��
�:;0��Z�(��U�x`Y/�N?�����b�"b��,������{?�є���Ю��=�CC��[��0�,� Y3Ed��d�)ʷ2�6��urn�8�|������~�����U1�s����G|��\�c���9B���?�t����j,Fw�z�|Φ��R��f˗�m�D4�1&�����������.��B��>q�*x��Q�y��=$�zLo���J�K	�d�:zF+.n-��3$pu�"+>�"�{ZnB�� /�_�"�e�z,�7mM�`G��(�=C�vh-ӿ�7V�Ito�2H���O	�V�sI�q�	�d��tH��_����H����S�����./��);m����%���MS��G��s��"Ep��0v�j���fK��yҷ��\�S�_}�/��V���_�N���R��9C�Vz(8�Wjj��m�f����͌�G��~%ݍ簺�s�!��3`(���f��e�08VV�/�k�4P��@�p�WGc��"P��H�)#�8�Қ �-X"
��2
ǧ��}����G���b�*U"WU깹�pM�h%���Fsm+��6���$�H�B��N���-�����W�wiE~��,�����4^q ���aF��l��r�모/���
&9?��0�Z���P�H��N���(,}0�*3aUk���l�0R2�7��[������h�ؘ&�>h��iuMCɥyf�!s&�:�4��@���,9]?���!���6��=�c���Ŕ�i\�|��'F2�:KW����o�9�����b�[z i�M���'��ƌ�E�TRīܳ���O|ZzzK����ݛ0�#h�8�F$�1��lH�A�D��� ���cz9?��O_�>3<ŗ�Ś,�T@�AO��
/.R�NM�Y���Y����.��3�\o�e�I�đ�$%F��iA_G�S�I«i��^G��D�䝈^t5#�s�&��Y:�$�k�PA���akg�i>a>�.���&�a��4]��`�S��w�*0
 �h�~��H"�(�&U�����1s��mg8}�K,��C@O2qr�j
�(�av4�J#����N�����&���y�=w�m$��!�T~�@�ڸ�t�����P�B��y�]Դ��qQ�$����Т�\���%���qm��?�t@����&�LLL@g:��-��>�	�K�Fk2�oH'���d~��s��( �Ȩ^/[�YS�NrrrF{8��Te�YI�&K�D���y���Vbs3�y-M@�Yx#i��\�y��y����kk��;p����%�JEq:�i��5_�D�Z(�>dt�JY��l���1O�aԓ������ץZ��u��mK�%4�H�rS��+�DF2 W@��YJD'�����r��iE.�c4ʄ3�E ��c;$�؝�	�qZ�l��D��L��I�8R���2��4���,�����Sw�>3�7�>u�i�ri�D�!0K]&�uUR*p��A����A'ͳxd �
t?��/�5�%:w��HQiI1�1�����z�H�ԯL�i�\狰��3��%��ئ�
�=�P.t!�R�
�G�����LH�N-tCGwe�I��I�68^h��4� �ʚ�Z�2f��y�,+	|��TJ�0��UI��#Þ�y�a���&��9�B2"d4jl�~��*�hP^��=��A���M��E �@zE�Kx ����v�*M�M�j�:�q�4<TD\LD<�����d�OU �J~��;|ܠ������(��c�8޼����0╒��uR�g�I�偫�(،���a���*��V�������|	)L��G��7�cb�HdD���̷U՚މ��IڮC��&y��fMbN�f%2��|ײ��zWÔ��
R$�N1��3NL�H[qT���
�w3�c�X�g@ 
�8��}6�Ai�]����0F-�DJU���y���2�%~/�5�侹{Ř��&I˻��1�"��՝���ƾ��ԣ?�[8+�\�KZ�H/i�7^�f6��0U<��Q ����|��W��p��3����/�4��
����kX!��م1��	VQ7D��r�YZk�^��E����V0n��lB��L쳜�U'~]��&�w��߆�Ƞ���~�� $:6�֛�JW3=�e9�x��05��]X,����y��F^t������h��Rt��M�}1kOj�}1x*�0��C�p����HϦ��q���{���Ui��VF�[���c)����p^;�<����r��W�g߱w�G� Uh3wÓ-͞�^��V��_~�*3�4��ʑ7�Q��� n8/�$�0g��+X�g�Ӱ����K_2l���f,���%�n7���>i���A�Y?`ԏ���qUBO�u�22�(P ����-��g1�����=*��F��m�;	�X�1K���!���J��rIq[>�)
}oUD������wm��T�p�8J:b����\s�d��tH��Xݠ6^��0y8������o/N�����	c\3�5���5��d��E����8֍����|ƿ
�2��r�CֈLQQ�
��$OU;�%ީwV��^�"v<il��AP��`�w��Qr��� o�TƼX�,K����R��X`����W!A���i*xw�?��'Z�� �hE`�ۄ������A�ZΑ�"y��RK]�jֽ�����>\��=�-<�~e�{��]������Uo�`�G��"b��Re5M��q u����*�Py��Sc�^I�Y#�����D�u�d%�cdА'�e��ZW���u�"M������2O��f,������ܖ�kJ
�!h�S-�A�8�W��Zw[�D���9$��<�^��/����D��}�h�N^��?��1i?iAm��9޾ ����|j�Y�"� ��F	<�\���*� ��˩���W�>�����`�|E%��먣��@�J	�<���CG���|�I�q޹_��S���1h�3�gB��3C�eX{Į����ih����{*p�]9�;I�?7�D�>\ɕ]�^�D���%���ٌH��$m�d@<����^h��c�$�S�Z�Qc�^��	����t��i�R�8g�ۋ�������7[+���`�9�?i�=�pY���le��&��������@|"#>�YiĬt��,��M�I�p`��d�P�����%>���gu�u�y�r�(�S�&�������O5�:�cRF��.�V��p�X�i�nw�$���V�Y�?�@��03��*�^�ş˜����8���1�x����"���y6^q�f��S��ƇG[���8η׸l-\��#z-�gn�1�+��	XLue����c���Ė��w�����7��_�s���Q��5� T��t���d��$_�ɸ辶�c�����\O��f _�n+A��Ijb~[g�G!�yZ-;gfÞFnR��|z���nBST]"˝ȡ���@s�p��r/���.d������+
�E-��$�@xC� ��?��eԁ�g^A�"'7� pE�ju��^��J�ߨ��㨥�x-�	���������bY��Gu	������]���=f+}�%1����MX�b ���z�Q�-M��=9hS���DX�C\>J�X���u4������7t��J0�&��:i��ǖ4r�+�A��"��b��
Ls���B�v��w�qT)�D��{�y	��/vZ$�;�Y���a���N�������!v�ߗ�U.1�aI�`���x��"��������p��tn�Y0[�q\��×m���=|V���#�w�~W��m�c��g�@��s��k��\��,��k�Xd���=�����g���4Nd���J�y��+�jI1���).���iԈ.������#�!�����}�[̍Λ�$�n4䷐s����BA���y�Է��зo_�	��__ Q<�a��7���{��s�Qj�� �7q6'~K�B��@��5�q�K)���*�=�r�*w�0�qU2���ɧˋKrD�����O攼{	���NPMv!:iZ��5�? ��^�'F��TO~��aw��y,b��I�D �w�زz��Z��=���H��oY$�tEO�AxN�����?�4��oa����O��O\k��ٽ�:��־Bp���1(:z!�m�u��,��d��t!h6?qp����lq��ת���:�(BJ��PK�!�M�;sn�����u���D {�SPD`\ޭIg����ݶ�ђϨu�Ҋȷ'���*iz����98S,p�~�{c�㱓�!�,*7iX���`��9΃JϘ>���?��j����e��r�z�6bp�LHNo9�����F���o�I����X�ڠ�T�'���Kʗ�)�/�B�c$)���Ԓ�_�tA~�=��od_0���h��Qk�(�(��9��OkzL���-��ϸz���O$����-�1�
�u�
ՙ	cA�,Y��k�yK���#��v��B��*[����=����Ϸ��Fz��p���E�sơ����P�ي�9��G����\
r��:�)��N�S�6j����C�S� Ӂ���N�|r2�&Z"�ps�ϝz���s�P!���Ùٵ�q��� `��G�J���堋.���3 ��W#�{�]��i'��u��s=�ѿ%Z�ǺՕ�t���0���N�	���N��c��3��_y�H#���Y1�q�U�{�NZϏ��I�-�@ Ğ��7��PUV�p'Pz��Q��Z�&勜^�'��x�gC�!H+.0�5h�OҤ<|c�Tox,M�X�q��2wv'�s��ik�ۜސ0��,%'���UPo@p��@����-�ݧ�lM��Խ+����Y���}7#'�W̬n�O;t��r!)�O�f�o�?(;h�H�'i�]��G�0�c�R"�vA�\����vs]b�yV�k:lJ�p>������i���&Pz=�y�Z}�z�������^?�0�x����P�-��@�m������rkjw3e�bލ��ze�V���z,u�������}�|C?�EZ�������4LzPf: i��X�~�P���	�\���5�	{��{K�Vd�
���eq�b7�k/@T!��� 4���X��Ӑ'c���F6��׊���M�2� � U>�K����b3�Y��u�����M�����5��U��4�Tko:���T�~K��8]�h�,^6�ip�_RS�GE����Y��VS^�/R҇wf��!� ���E7�)%ߥT���(د������?U�����6g��	!�6�,a����՛+��괥��O����M�q�}��q�<��@��(��aA��ŃN8b�~�$A�E�uIM���5T��R�_�ִ�Y?4Ȼ񳭑�'C����Je�W�D�?O��dq�6�=5��P++��:n���<���O"Y���OP� $��U�S���/���
�nͯz�\F�
�yAY���<�.N�T�;`,Ig��ދmo@>�iJ}�uǸ~�vMG����M�5��]=�FB3��H+bGk��%V#+�CϦ�0��雙��MTb*�
���i�ӝ z�e�����Ol{`�q���n�1��6�SC�!�~Wr�^f]�!`�3U��ȟAs��̺�X������I�N�Tv�B$�� C��T80�%��S}m��gu�{v��ѱ�A�$Y���K��j�q�o�S&Rd��.���=����!��#J�i�KC��.`J����M�Z~c�r�I������B���r���n>Z��-��@n4ku��Ϟab����Z�,��ES�Y� �۫�A��Y[-O�����ćn04S*��M=y��j6ݴv�~�^��$�X��H�q�f���?�k�=�r5�;6î������]m� B>�������v�X��-Q������9�W$�@%Gp�ꅩw����T�����+/D��'w��q�8�r�,_���b�\Q�X�-�NZ�7G6@���-��Oj>����s���\7�Z��d��Dq����,҂^���|7������������>��*uAZ���a�V&����뇁�̳�wK�w-�.�!�t���L�=����u�NQ�M��k�cU�L�y)�Ɔ�x8Ӱy~xm����c}�*�?�~N���~���Q��d@�2&�ᮯv��c�=p�������Uv��C��2hi̭=��]�����H�l:��4��M�/,�P��g�V�FY��nO�#���_�<pxoL%����|u��h
zH�?5^��z� .`�S�����j�^vn���-)$����RVKى��u(��eMj@؃S�\�������j�l���E�@���J�Ex�N�D�p,��ޝ�hp�x֛O-Q��ql��!rW�xX� v7���8����!����mgԪ�����i�.븧��@J������v�h8�a��tiN1��]�qE�l�3��_լ���7@.O��g��&�hmy7)�~�|�J��`\5���l�F�~������4���]�[����z���*B֤��4����?h��%F5�v�n����扞���tV�R�e�i����˺��ˍ�	�;X�j�|�zk����)ET)��ն�_���Ԋ`̨��w��	��7�gW���ԃU�A'i�}���I�5��m�Z��~	N�����"Q���+�����9�Մk9;������ǣķi��^yM"kn��������ڲ
a]B�>L����8R��y���g�bP��n���A˳|�Dg����8�# �9����R��/��A��<�����w�	NBt��p��O����\}��(X�/L&�h��5�ߋ5-�7�7d|;���$��͋�H������FWui��{Kb��ԏ{w�B��`��eCR���q*b�X���W�mu��C�1�F��E<L�;�g�o<�<�	h� ͳp#O3�Z3�p�|��qY"��	%I&��P ����uZ.��!�ͼZl��a������'d�1��`�?�9��?|vDugU~}��y������]��˕̔��0��&�{��|K�h����Tw�:��׻�P�en�V�?ܔ�7'����P=ݖ�C~��8��߳L�LƏ���� K*����ɛE���/mcxwOz�}i��Jo�p�[��Fa��@�]U���r��ˣ�4|�[����[Ch��lO���z8n�6�������F�M��A��BL��j�+{m��X�����<���	f��޺���#k���c��K��:C�W�Q�}g�N{^������D˲;DR�c��������?U"�J��s�B4��'|ð';�wTZI�{�/�����w��u�r�n�;`]b����*��#�7��׽E��V7=��u%oW	N̶a�%i�)����߇
Ndb��	;�d;4˽+f�]�Z�7�HO$u>͊�Y���dGl�C����b�C=?1I�����[���@�G��K����T>[1��Gο��ߵl^)��F�w쏌<���o������M�c��*h�|Tg���1y8��[��7���d��h�: 6�d]��� �����Q1؂�#l<J����W��������R��8G��ٕ�Ƌ� �J����E��Kbg7��9��}�>_��vZO�q@`7�:wkQ��Z�)����Rw���{]�s��g8�����O��Mm���u�5�#�CxoֶF�·����D��A�B�����ʍW������gb�`�C���y֯�D�7*�g�i/��� ���]�#~����b�;���l:~���!��W���":���GD�G&A�tIc!o����G�d�g uHXdڡ.q�*i��Tw�b� ��Jx���r��N$�����$��u�+�K����Ū�_5���+:?����(R\oQe�:n<�l��5�(�y���9�<JU_���VZ�)�p���;��&%!��`�:ɵ\�ʳ���s�ox.J�����1��!Q�H,�0�p�56�$��W�8�%��-�bPw@g���7���K���] DƉ���|�����?�f��&����o��%�N��Œ��!MЙ_b&�"�ewX"~P;�k��k7�-**$>�����"+%��=d`^%{V��2�{�J̐""�#���>�%1�6�ںrȣ�R����B��_ϖı���b�f�%���+!bX����ⳕ�>���Z��N��3{�������1;χM���iE����R�؍1lO݌Z��B�ө8�(�
l2\�[.j̟>�F�z���hY��]Bb�X1,垢ŶV9�X����p����\[ܝ��˝�+E�r����o�PXg9Z��-���ag]�Xft�ƃ���\c(�Q@Oy"hg"�<���A�M֟����¦��ͷ��ܠ<�����?B0����[ׇX� �-*ߌXVow����߈Jj�Z:�H��9	b�]��#�k��K���:�tՈ�h`-�GFrM���D���i���_�>Sΰ�8�GZ��2��������"���yV�:D�5�x�ކ/���l��ĚZO{{�"�ei�d;�]�-�^����*Y������TZ�ŉ	���.��
S�K��cd��P��ĉȼ�1^���i��^r���͔Z%���+�,&��HG}U���E��Sr��.P��'��b��yX��װ��{�vډ��'y�ݩ1{�ip�+�+ɯ Ū�H�m\�l:ܶ�tQ�i�\c���K.���}�/[���j6J
��i�Ƶ?2fO�	M�=�O��b�쁍���ۣ�j���Rx�IS��Q�g�we@w�E�U��/L�yy�'��ǖ�EXYb1��4ЌG�o�=�>�7��Q�ׇ�,B���r������kQ�31�������)H)��dЕWC�p�������q��{�W!����w���x�~z�xX�')~�N(��mW�:�k�́���M� TeI��i�漏����%@E�9M[�a�:GJQ��,՚���_)-��@���ǽY�dw�t+���|x7|x ��x'����Af�|/�[r�_yZ�?m�YI�o��t���,^�Tb4#nLx'�萲�~�&{�*���/���̨����r��
�SIûj�O�ep�����q������,s��Se��W�!V��=�/�aֆ�s.��x(F��c��9h�פX6-��-Y�騫!���䍓����I�{��J���J��]��������ß�<��r�ODt�1�GҙKaS7��	������&�������<�޷ُ����Q�\,������&hf$�B�+_\|�m�Y#P��-�6f���a���Dl��3V6�}@�_U4��?\}u\T]��� �Ҡ�t*��� Hw7R�RR
Hҝ�R�Н҃�t�3�������᜽�^�g��9
e���e���ǌZ?(*�	�/��$�N#���q�1�r��\���� ,d���覦��r`��c[�p{0C����]q��nr�470���{ U�/�T��]2$J�6����H9r�U�&*����������?nӠ8���@�,s��d�`��P�6o��Џ�q�&��7�N)O�rs+w�(){.fY}8�x�Xܘ4�e�o���x��U�� &$�'�rv)�pqUQ�)��5�/��Ά������3��Y!&[�f\�pj�&1�}������+S'�5M	`�%����I!,�8�g�k�U=T	0�M��>���U������2WS�vHq�du�?~4�ߑ:�ą�0D�*"�����K4���B	6���a7�Mr�$ͥ\7VR�ӆ��|*|'��Y�w�������5Ib�u�[�Փu{yM÷졿��NQ�I����gf&l�,�hAƣwK�z�;%&LU��W���#�$��ê'xT^�<טJ@U���tp�-�t.���g��\s��s=��.�w@���!���I���a�Sop��p ��L���c�8K{��V��]�ʲ�]>�9�n����@��
��o�p"���$���DG��*�P)l%��Y99U�����z�L2�W��$�*��_Q��/�d��F���!#����H��4��:�'�>Y�B����+7 В�D@M�:,��s��*t}�e�Gd���anp��|�k�*nTz���Bf�x�]Ǘ�7�_�9�Bw��$n/6��Siy��9j�oO�+�զˬ+H�n��uzcH7�I;'.��%���.�D��'߫�]?�*��f��|�H�s����z���0*.�xKo�(�/v�k�ا�[�{��TZ��ST������Sx��������p�OFI�7�IDԗs��'�����9Ɠ:5}�F���-�,��p0Hi�WWW�<�}�i�H�{����k�|�%�F�?�gDe�j��k�͏�Q�Y��S�ϑ����d�&�:�ډ8R�c�I���{q��3�$t���)�9�}��P�<���;in=zN�ıOO���v~Hq�m�����p����Dp�8�Y-#O��AK����l�Ϲ���|��E씜<#�+���W=�!��z;����F�a� ְ��C�9��ph�S�Sքn9u��h��eV|�8_VЭ8z�Pp������D]F~Z۷�ǥ^�5ҽ&���q�1�Q&L1�����5J$�4��S�ۥ{�f�ĥ��H0�xؼ,P�h��~�-�o�İi���z��u9'ѓF����?,�k���
�D!����^��D�T}}�b��c���E��~$�|i�zC}CS��_�4��J����Cp�4yz*�U7��T�6\����6�7��MUBI����X�r��,�v�Ir��8PX�S����壾����DTi�"��t۾�"--��=�7������(��:�^�aDyXٶ�6n�H��#�=�V�c��N_=��k�E_Y�m�ZU��>��FРa�@b�����kצW�m;izt��'����O_[�[[�|�a��4(����q4cě�!����֤�`��9)<}tﻮ�I��j���XT�d[sH��9˧�/��q�F������)��L?m����E,V2�;*0ff�{0�%'/�H�|�MI�i*��3���@�A�怐�qf@�����/3n�Ea*Qo�5<ʗ�.S{����2�ⳡ��ن޽�'�"6E6mj��|Z-��Y:ԥB>wT/�$>�o+`���K�ӥ"�2����H���S5�7��)���k�Xab�M�Qؒ@gl؁�ཚ�d����ގ�I�r����&O�ǢNE�%�B�dR/\FR3�b9�T���$M~�UW�d O�%���Yf<�nzn�ޏg���Q)=Ksz�a�X?!����m���J1�ͫ���=eL��8(��>�*���n�d�}�/��Q����k�<���+#�d˭�o�Nl��W�*.��e�C8�Ǜ�\��ct�;D�b��Ӵ�"ð	h\����=��\3L�s��GPtۖ�O�q�?�/�D�2=�X�
�*�-��]�P�{vݙ�����W$��3�qbes�k7��ܪ�R���"dir���H��&~iV�7��xM�1$M�8vQhזR���׾8@�M唈�: � JF�������3�\��,�۲[u2W�=��ޘ�`<�|����%��S=\8�W9��e5t�����<z�)Ȁ���K��P,�#D��,������m�Ȩ�[�(�\��Wf#��Z䣧؍�[v|�nkۣ�HI��/�P	v�OP�6��(S*���?�{�0�������n-HR���N4���(5$� 8~~Cm��l�G`�n����0r��
��p�"T��Ǯq���w�(����I�I�ׄ�"sw�c��uuspC���i�b6Z�8�����Mb1���R|�ln<ז�mE6�~'�R/��~yd��N��tt��$}����^�]��x���c/���+0�i��_(5�/螃./��iص9���B�qw��;�KA�}��0a�x7���a�9PbR����vQ�~~o��@	���qt	ɚ�nn ���լԬЩ@��ٯX�W�5�B1�e��BCuS�����GF��7�cz���e��ȵg�T��E���uR�Y7��e��-�b�C��(/�~�o굒�n�E,��=���\s���lS��ɦW��D���[�'#�dʾr�9�����,
wBarWs����0NY���'g`=�?�ż��権8 �Jm�M�@�<1
n�I�y�K����=:����2
M�@R��d�@1X4�8g(m@ܷȜ���^壞��O~F�<j�Ώ������o���+AXԦ�i��l�k��͎hî�B�?~3-�������SR�L/NН^J!����L������̓��ވ��{���ݐ����Te�������R�9��,��ȸv��~/^dzz�[�پ'�� ��Ŋ��ȵ�)R&��O�'�M|����ϊ6�|&Q���14[��?9����
.�r�qK��CN�ԯjt�{S����A����� ѥxV�AI����r[a-�T�E��b���1ed8?^�ddH����߇���<jvJyD>Y&�=��]n=(�xC~�X*IHjM��Z�W>����x�=l��>���Խ�g��`��������Qђ���� )D�䑟J���wn-o������,~usx�T�)ܲ��blլ��>`�d4an~Y�Y8[�0�9�/X���{x讈I����po>�L�A�Ғ��Q��i��{J�����U@�<[�(��wy+ ����ʢ1��7�ݾه�{;�����p3��,0T�{�뿽 ^���+���'�����$wݳ9
��t�l�.s,�b���~h��8��N�P��7D�9j�]!�T��=*G���moT�9��0o^�(�����T�����B@�ꌨ��F��\F�-�v����c��pȥ�7-���J��2���fi�e5X��'0J|M�ϕ�W>�c��9"��i-��h&l�L�;��/�HrxT	v9��g�ʧ���MzMC�B�㗺��ج��/4�B�E�*S4�te��?��~ↀ楢S���bg��4�ME�\�|�t1d�S�x ���šqav��^�`�����e�+� ��yAR�Bc������ق��;,\�՗2�<R����Bs�2�sF���M��]�6���]���j�-߷���9c�x�.��& �t�x׻ȳ�����W�E^�Q.avv1�z�e�D��9y�<��4��r�rV���?US��bG�god�����dE=a�H��T؈�-�?I�(M�Ǒ��4V���>Ϗ������U��[��p
�b�snL�IRb���Ŝ�/,��M�f<���!�}��d��g!C������k*hٕ�򅇞��M�>M@cK������Y��!RqX���vp�B��Syw6"m���/�׵	o�}�a���{'eG�bq�-�5L2<D�u��i��,�^yo��PC�jc�Be���Z$؜U����"����>���~�5}����^ ���ܛ� !�r��bwFo�e���9k8	�鿢����߅�W�~"�ǵz�Xl�#��|��s*n?�"��M�*zX����׺<�1eH<eO��>��� ǜ����9PJ���6��b��O���^�v���w�S��)iG�aY��o^�sSy���ܵ8h�%�	��Rm��)<,�@���f���uj�^�ȉf�_����4a%�N�@�as�Ĕu,���Y�������J�u�R����"<l<ȧ)�G4��K��p�9����)ދG�?y���XԾ�[�XY(�Xb T�D/O��=��g��QFnfT~!�!`Y�eѥ�Z'�H�$�ݖ6�d�M@�}{����6���S��|{�&Q�O��uYV���{
u��,2���e.���z1��}���p6��e8ʢjm�#g��@�wk9��o�\�۾M�	2�g��A�sA���YsR5����q(���ꃏ�f���;P�k&m#��v�,t�8�_LU �<�q�A \b6_>W���dQ�-���)@��o\�Ri����F*��y��%sq���0���:�D�5�3��ђ�*լ��u)�ȋ��b�a�U-|�����ia�5]
�|�Ue��x�g�{�a��ԏ7�Y#q`\�)�AS�L��\�R�zTĜS�f���v��Qɴ=zm�衔�T�`� ۩���O�۽��ufPd5�>R�\�çZ<,T�^8xj�1���װT%k���ꊭOS��K�z���@�C�Ȳߪ�D ����=�y��.��� 0������2�'�9C�?N�r�zѰ�C��}����#���]�kc�H�A���"�F�NH�G��2.��	�+��!T�`BǇR��ΑDJ�}�W@�2Ê�4�jP��-���~��Y�ؘʦ(���!0u���D-��'x����8b�����|^���d�]��e>i���[�ǡMWN����Lx��sv��*\��b慚s���p<�j��eؔ/$��������]
�hk֡H���yԣ2��<V)���vI�y�j=G������mE�_���V�&��e4�1�H�.�8@���&�R�:�׋��*�C�zNysWa��{���ڂ��o'%E�?/�hM���|m�b���o�^��S��~�&UF�xσ�hG_�C�� ��t������BN�������>�ȓ�lKO?C"B��od��Ļ��CP[�p�Q��k�j��?B�ͰgX������t�ո����ż��iۺ���M�@�Rɶ`��4kib /�_5c�P��;(�M���-q�5R`} ��#�9k�H��k���1�V��dv��[��]����>'*E\��t������qG�S�b�ag�b9�F����W���qIע;����#�iGX�j*$�'��y�(��M~�
:�En��_wA�2Ît�r8#����g��B�+�v���BӶCJf�����P�ġ��>�5����8��!w8/�w�X�Y9����.�%�q�>�M�M���hR}P}z�[Z;� ��/EO^��<�,>v�p0x0�}��%B���螺䜽��#��0�I��[��4� ��v1T�Sr2@�t��u
�8�M��Z���0�q�7'o�m��S��
#� �X�Egy?��x܊�h�!��93�Y:� ��|�3��AHW^V���!I�գ�:twn�y�]�����$���]|����׬q���,�{4����Ԇk>��B���z�,.!�.��]�d&ĩN��:�{~e9c���;��T�&T���7���k��#���h%��g���b�Zi��}6�rF�o�'��*j�+�}��d��i�7X9any�(�������h��-�ٷD'��6>�'�5������gEMWe/&�/��q7$�_���w�����Xv��	��F��mH~o8CU�n��B�F�V�0C��ۼ=�1�aO~nq/�Tͷü��l�p����#�Gl��;��Gl�Bc��+u���w~y5q���d�~b�v���U�bCtҲk��\|Xۑ"�纓=�E��&v�6���w]�9�$pю:���0֎����s$���&�@��H��/���B8ȓ���쐞z��r���8�T6Bwߡ��`.Lz����7��@�����.X��9R{�I��ًo�DVЃ���2e����;!�ʶ��$��cwφ���!Z��=z��ϺH�����$t�~)o���������'�7��ۮs`!� X��nBs4��p�@��1f��q6 �J���w��������^o�M��PWv[���>}7���VGؙ��D��:��'U�����U���Sts�s��'��
���&aE�X�����C���5�:*ס���'�&�Z�ȆL�X�1��KO���õ ��mi5����0��uO���@،�Y45������m�\��h�G�����8�ǫ��E��,Sk]�5����uޮP�p#�2�nU��AW�s����MnQ�z��>\�95�t�w8V�ن<�
;���^�b)����{n����ċ��;�I��7�fK�p?��*��p2,�㘥��H��iG`�*I�S�S�,��V`�yL��0P��q��C���6���HM[���%�Lq��z��]��"/����f��
)�F��~�K��%"t�$o��oa�ѫ׊��X3��0[R)�@
C�&�sG�4
�S��l�C�j鈿��7�4�)ZG�WKr������u��0
�E]�w�;D	Ui�O�u�]q�3`4���w�^�Go*�ł�d+��̬�z�`Y���`0xL�ق�^����nh@" n���Qd�Sks���D��|^����_B$KC���~G���7k�G�7)օ�D:�o0���	�m޵K0h�,I��0�B*}n2w���_l���1\�QM�Q�5Kq]>��?.�����t�/(��Y�8�	��1�W�?#�4!�D,|!�S�k�	�5a}ږ�0P� ��?&��׬�k��K���5nw�#�eLDg��2t)b�4Ai�5<$��F����V�G�]uŮ�3
�s�:QY|,d�
?r,�_�3��v!6���Y�ޗ��� +�v���26Hw�I��g�)j�/�J��%�9d��G�<e��Í.�P|OKz�g��+n����@θ+�	yh��P��0eAC%�>rw �������er�@|�>��_�9%x�D<"���voIA��+x����$&(4s87���#Z���t�����o#��/�@���	�?�:�+�JIu�\W���>�����pt+n��i�E�jy�Ο]?Y�	����N)C/Q:Bjm��hh��"ˤ��gmE�[N�2�+5S$�}�t4JĐђބ��h�Ǯ�1X�}�c�tr�b��_&W쭮n��A|�*3 ��H1^iߍ\?F��l ��(1�b5��Ų���NrE�,�[r5Q��#h����W蕯�o��3��~������
���X,�np<�za')�o՜�.jg\g���~�c�0��sJB+E��NF�r:[G+��E��+�o�kU{1����M����I�ŠD�i�(��L�$D��eW0_��{�������q�|�e��y|c��c�8�[�V:j��C�(�.}�Î]O6�k�M��p
֫a���x�+���[r��l�IӼ��TLp,�,j�B�j�ė�q���`9+���1;P�b�0��I]�@�|S����ʜ]r �.!�	Ƨ�M��q6k�B�Z��i"��k���@~?QS7R�n�f�g)��=�<�H���yU����c%}hb���*Gl/hT���EE��H���Gu��+q���.���d���kx�k�R�G�g�M�����ȡ�������_g����P��;��f&tª���esF��Tij����Tj"&�~��h«�?����pzcν�I��K�-!?�Z�����b�	*���8П4��q{��G�@Nw���t2�lkZ���<��D�F���b1qS������!M���p�n��'u���k�O���r1���������Qa6=�sY��;˩�ހ������,�[YO����9��+�#��i�����z���y�U���RY�4����К��Jf6!��ŦOB���4Z���}�eJ�K�R����ەHR��;�C�E ���	���z6�_S����$���v�nYZ��^�%(·?�R"=��ňuQG˟ :ٟ��;9�}L/b����Xz̨;���Yh�a��]s%�3G���^��B�"]����_����[��a�����,���M��O��n�R�H�?�PBL\���������)�1!��te���H�z�i���'(Sb�[���d��������`��9y�.���� �eAϏ�s�oy���(��t��cp���]^�uA������&'�ڞ��H���}*/�ϲ����wE힣���Y"�Jg!�2Ju�@���Š�[I���K����(L(�Ɠ�g�O��Ox>
o"��y5��I.�<��r���"�н�4I:��o���x�����u&��!<�������L8�M�.�4���,K��_�K� ���z�N]��k>�a~�'%D���$���:�@:o<�mIUGG�o�.f����ѳw���8�oB9�*������ �Mgf��
0�N�����`j08�/��"���&�R+��;+㿒�l���7}��G{w�`8�}�A��|�������x���g�����D�xqW�
�*�q�/�_N/�/��J�EIAL:�r��	>�Zד�����X (�Z77V����&jV"
�������^~a��c��EV�6��f����[2�.ZR��7��[�:�G���e�׳|���-���rR�ե+��r8#mm]��J������ퟮ��نVXc�z�$���$=���)QJ��l\�"�h-&ɢ��HϠP}S����Ԙ'��w�*�������Es�-���/��s�'X�_�pn� d��e!GNC{d|l�&򤪰�?(F�WÀ�+�Y4K�ˀ2�e�oD+�ƫ�ꌨ�|V!�ұ�E/�Rv�I�Q���t�% �}O��1G\��Z����!��C@;�%P^к<���6��p0m���ayg1��?}�80�ZI�{��.՝��Tf���y�$��0hx'}��Td�������@���0Y(_�X�W�m�'����+T�^����Mp��=Z�A~��d]_��Ss��.�<��/��:ⅹ(�������[�IT��?#&��6�yx�����>M�?�`��*�Rw^î]��rvlݡ_����x�Z����5W��bo���Z��(�G��1Dq��y|"C��d�c��kQ|���-.�۞���	�z�`�V0�a��ɣpH!�E��YV�@PJ[{��yA��в@r<���.������@�ic������\��Jқ*�Ө?¶����ۋ���*j���}�&�٘�!��JF�n�ß�{�즋~C%�w�t~{t������?�媭 L4�/��:>X5C�/�_�V�n�a�Ԓ'� ğp��/4��+T�rN��P��oK�t�,Z�z�R�TV��ӧ���:9�P7�b�os�w'h��r
�����V�S�9��Ք��J��>9���z������% �B�!*�����ˉx�x�Z`�ZQ�m���zYW;?���< �l��3��f��E�H�I4��U�ǩKY֫�&� �vV��̝�Ib|�&m��_ r��g��R.�Ӷ��d��&d���"�O��E`�x:�o#{���pZ�V�_OL7\�| ��Iq�]7J��yb��	R���oC���86K��[�?t��D���Oh'w��%}*b�c���Y�@	�4�4�p��DX��ܝ�	�0�# �s[���5*S��e5�E��!�.iТW�Z%��v]��l��� cDe��N�ğ�$~m3�]S] ƨ��ǁi/Z���x��P��E(�u�0��S��?%+�|b~�Nr%��TNW��%��r_?��6V�旙�!��qR��1R�����\ǰ X�=9�i;�#UQ����oS+}:++�`E4�l�,��&�P,bY�r���imS�s���a�U0b��b�����Yc�����{<==c�yk�܁��N�u0�ȼ�+|\WP��U��,��8Q�٤�B�E�~����b���Z���"R�ndt�{���V�3�mB<<�Y���K[gY��?�An������軇�������������ň2w�[?����e[8�~˶m��� 	!��Dӂ�IC8�4x
���'�m6Z�ORy���(Y{z��H�$�I]��X`�O��y��A+z�f�?4ǣ�f{7����m�-CB��G�	ux0�H�����(Ê��d$UU��pC�l_v���Q�W5�LĲ/���q��r���/��=&$}�vW�ٶ|�%�EM����Ӆi�F�����z)3�a`/�afa�I�?c�c(���+ҏ�X�W5��x�1��	yv��j�y��~ڼ�yS_�5�wK����bDE����	[��F������O�o�+�%e��[<LG�%� ����#��Aú���̔ca�I.4$r�`벝6z�RC_x|ԙ���5�c�:.H
<ut5i=1)z�Ȍ��#�O����g:e�0 D��{�Y����Y�i虇���'}	&l����e� �Jrst)N�2���M�m�TOh D���\�?��&����W�~tȀ�%o�!���h+N��l�TG�L�{V����UR��E�}7�\X
=l�B Ic��l�3�I�i�e$ \t�dW�$�$ ��l�H��CO�T%�h�O�x8(I*���*�c�:�P-���:�%C�8��J2J��Y2�悰V1\�J�e��Ŭ�n �������zm�`8hS;����T���GF:��TI�I<�]R"87m�;j?��YJ�=�(��%���}����k6P߀e�	�}q�8�D����E^��@�'F�lY�T�=��چ�c���cѢ�N'S��q�6)	rϋ�Jʰ�$�)DRZ���2���n޷L3�Ȉ �D[�=bMS.�.�5-a\=�Ə���s�B�6��(�<�Sb"_�u��n���]d��,k�+Poz��,�G ���f�yƜ�[�DX!f�@V4���B�E�HV���na�-[8�<�1���3#9�##�"��w��R!AY��@�r$ X�g�'�l2F�>V�9\�#��{|'3s�->2����[�Xc�9n���:L�h���h��~䃂
� �i}R��_(�c��=@tמ4$��0Վ�z.���78�Q`�#}]�4k$Du⇻F��&��j�,)�-����	�/K�/�ΰ�lp��(�E��lu���I�2��lč����2�ܨ����^`�ר�3�����ڶ�3�h�B?,}�������<]�L��|��T��Lk�����4�#>��ʣ�tdD�E�pc�{H��|�,`�y�}Ԫ��w7(�E,y��%��u(�9D�94	�R
x�]�S�=_�J��`"^�b˗iې	�n\�r��q�o9�	��{��Ëz�1yCq��\��|�Ly��4�F �)���<ܜ�{5�+5z	��� i�����wl�&��nm ��{m�c8�ز3$�9bd��#�80�Z�~y���;.���"�ˈO���؝�ϵ.o)��8�ʫ�w
�gEGGG�;M�J� ;���V���tmz�)�[TC�x���j( ~K%��Li���(�8�n$�\IП�5�K㋊F��+VΣ3�tz�A��f�һd�䫭���{�����7�*��e[�y�@��C�����VwD���/O��]�U�#%�TÌ�����|O&��|o��J���o����"r��[!;f^��������;yb�-�fc�Ԣxۮ�'��S(�Jq6��\�gMHO^��Z�d���1��9L�y��z0]��0�B���-���N �FiJk`�.�,�nY&����&#c�0q�S:�0��tq��IϾ�ir�.ڃ	��XuRZ$2#�P14��U�f
�f�߅�x��U������˹��\�Sq����v���^�|�t/٩�'���AKc�݂4Y��k�f�i�a#6D9�/�+Lj$-"�@wb�WMl2,ԅY}�{#����?��}��g)R�~.?�:������U0��t7H��3�ז7���ɰB���b��4a;�:�"� �ns��� &׍��U��7� ��(f
���\�vo5Q�vzȮⱶ�]`��	x���&��z�;�~κ׾f�<^��Ru�'�����_���-�#W:���eNd��� ���*ְ�$\Z��.����*�k!�){\'G�oɎ�dܥ�~0(@��cT�j��B^~�V���\VQ�m�5y�[�XX�[�rT�J�!��WiH��o����{&��m��Wv���'}A���35�	��RN��(������π�}!����\�QQ�_���,--齱q�gg}�Q��{��~�y�z�v�G�������;(T�Gl�m�;�U��E!Y����x��I�2ё�p��?��0C��"���AYa��[�[+-|5��n�f����l��I��;G��>LqJlq?�뗴dr57��7/��%�+��.c�~;]��-���hi��[!{{�#��l���BL��e��#������vB�P�P�`��]>e@�e]�3^[>�y��}c��F2H,�1�kԁ}�?e��J�f.�x�X��x��k%�1#r��oō#A�5�X-1�x��'q�? _�E<�4c3>�[�L's�������xb�Ubhϴ-���:�l�pyȦ�l�^-�u�2�mW�S,��#�+{H��l�9��U��@vY�j?�aoAɌ��g���|6̓�����eʿ}�pz&'=���{>��*��װ_k+m�{_nQ��ZɄJ��FJS���-uBb��R=ߐF�[AG��;6X�\ݤ�j/`0������<Wb�����z���;y����-��)3�A�@�u};�Ϙ�+�k?܊o��o/���F�k�����R��:�V�5���?J5{s����f�Zc/��vi�� �U�냅�#W�S22��"��������z.���9���|'DH�j��D�K[;��4�X;��5��!zĪ%w@���"p�]Ano�'`Vk(�x�����/V�i��x���zS4چk�!>���OB�.��"��SUMm`��9n�L.N�YZ�+�](��<W�M�5=gg������{W����oL�Nh���^�Kx8p���n��$d��	O���\�}Y�Ix8�� O\�>[!�Aڭ]���I�|Uk¼|75(�ɮ2�P-���Sғ�}"�Ը�n��C����Iٮ �!��+�-����}��W�� �8��QK&�?BL�*��è��[[k�r�-��|O牸�<~��pɰ��
����1�e�iB^^ټ8Q���|����I��M�2�e�&�w� v{�
���|g7�9Ϫ��כ��\?��a�´��S��|����?�c+3bSbH��)*�=!K;;_�������ۭ:� ��$M�������fq����W��Jx�_�@n���^ΐ��I2�ŪRgmBU��%���.@%B�j��4���^����b ���=li���R��8�7���p�M�J��Y���Bw�������A��@������ַ�]+K>�����8����!1���ا�vfR��p��O._���W�4&xp���9��`9���w6$\&�Ǚ^lO���a�/��n!"BZ1^q��[Y5�����r�8��4DI}n����.�*�P��X��)�>���_�H$=^Ѱ��M!^�'n�'�r���hx(�Q���[�J
_nF�Ŕ�������{��n61������]�����KC�e�Z�Kn����?�*����#�n��?	��,,ymp�T�r̔��, ���N�� �OQ2���{:]�k	�n��\��0sm	��
���kˏ4�����I�%�����OsTm�w�5Ko⸖�gsA��@����5���h�o<��U0,��Ȟ��^I���a?�q��o!��a&��������+Mkm�_/_M'��wkF���o�7�M�,�'?@�<��?���)��ib���l�j����Fkp��� 	6��t��a4��s���AsQ �O�J���i�?ӲShiAy����~t߇�*�Y�k>�o�Z�%Cɀ�.)��R]�5���5;Oe��dYA?�j���1I%:��'"�ħ�ړ�P�E	���������UO+�壨?XNY߃��:�w�TH�,�1��@U����s��|�kfyۋg%�������MŖ�gP�Bb��2r)vKc2�hcJ��2���g�D�`.4<��h%VA��{�3����|��B^"� �o��[�����^l6B�8�s 7�����^3��%*`@�kb�G{}�S��"W�vf-��A	��-�%Z|��-�bD��o�s�[_7��9{f��}� �����}X`n��(޸���2���D���d�,�^�����&A.n�j�#;R�_�:��*U�ی=������-}]��`�OP}��[�|Xk�^��kbR�[9We�Y�jK���l'�'��׺��J?K��|�Rc��_�m�\���r��R���O��z~To	b�;+Y�S�*����fj����埀�Q�.0` ��0���4}mW��`X+�{����;��ˊ����C#˅w	������5W���4�#��p {Iۺ����!�ե��`�_ �������hۣ�6�Ӥ�FZ�ܞ� �λ�ظ��靔��[�hb�dX_�+͍�ɔذ��39�4��4ݨ��'ں|Zm8a J��+�$�6�X�-�w�
ߨ�@���Щ��<�F�꽦(h$���,Zp��٩a=a�*[_{�([��IÏ�)�zz�4�G�-=QR���0!�n1s@	�`�}��c`��>�B�(o�xAI<51o��2�öEW�E�$���ٔ�ˠ)��C������c�g��L�m���S*��{�b�ٟ� 
�4���J�{gDvR���e�/�����w��م������۾��D�+�B7uZ�a=8d�rG�Čm����.6�+���̑�H�E��P�Rߨ��f��&�-�Y�4��X�q�7��_V��W ���u�h����p3ʡ�E�&��?�v{�@������������y��O�~���A��ނs�ڹ�8(vyepe��7#�|�������:���ɍ�q��T��Bq-�׫�����2W��f���H���A�#<A ߨ��$�?a�hG`�
��2�^A�o3+fw7�����|.N��>~u���X�J�q�U��e^n�[�?h��'@������_[(�X݆�4��(%�y�ެ�F��C��G< .�
���8A��l1�<�GBĳ��O���-���q�0n!�o�1�������g���5����-�liz5B5�}-��!4�l@�l���J\L�R�{���Y�&[��zܗ+�4�����z�Q�W���w1���Yݜ�4���{���XL����9�G�ߺO��}Cf�y�y�Y���/|e6j������Ӎy��%���ޟ��aE#v�x! 'ɦ�T���jx}{�X�t��D%6nu"���B�EhU+!Fߑh�R ��I�p�k�w�w�k��.�d�z�2���j.����ٝ�Cԡ�N3�n3};�*�hD�*��'���z.Z�O�87@���w�ϰ�������6ƾ�׫�����pVp�s;��SH`C�s8��K��c'�u��:��½=�b?���|�}fY�mVO�
޲����TC��4Qd�t�]��#ΰ�(���ʃ��E���(�M��������7}��A[�2��_��дjfN��i}�,���Te!�&I�����w~���ig��L���Y\�M�b�n���(
�C��?��L)�S0]9�s�,�\=�]�^�|X4���z�F�~��t�j$�����T�HHl�F��m���ki%A�AR���I<ͺP23��}�����iR��E��>�ퟳ�N޾q��|>��@ �/R�N��|Hfp���ȇt��N-�e/�\� ��͟�JW����g�s�s�d����i����ڶ��7�]=�q�x�㥥k��Ns�X�1��ہvK�Xk|������ⲽ�ޯ���i�I�>�Uqn��]����d�g��A�7��i36������?���{��j7����#�F���Z#n���c&I��m?����4Y3����oS�~�}3:D���]� ��5�] �ч��H����Ɍ��ݐm�g����؉�Q��F�-�Dn��I*P� �ؖ�Q���gU�W'����zB/A�q�Z�~w�KY�b�ME�̵�ms�_^N��@�*�ٛp�T܏��۸Wo��6<�q,��_I H�Ɵu�������ȿ j.��@w&;f^��݀a`�e��������:X��_�Z���3ٍc��2R�y���P�A�-�_�냾T�����mh-:p@2(G��am�-�ݢ�E��>�t������~�_�(>]�
܆�W�D���$�o��"� �.�g�^��22�6���2�W����<��4�<B�V\�s��΢�a=��_a1��a �|T�^K��#4��QZӭ4�������m'+���^v١���vȢ��Lb�bs��Y";_���z�Ā�Ҩ�B��8,���������ΰ����(�<c#H�6( A@z�3P�ދ ]� 4u�� �.H	z�&]���A:$�Z�w�������s�^{�{�k�u�9��qS�++�o�2��VI�Z��p�K:���j���*�n�h0b���7�Չ��ސ����:e����S�� 	U���+.�Z�\�n���B���R��	6��>S��>}��
�>ڐ�I��f��c�[w��ּ��1��n�d�s�Wt�7�;�N�B��?��g(����5��ԣ��,2L�OQ:�\��O-���c�pх�Y<)<ZƂptɄ���������=��{#�#�.)�M������1,C���8�N�-���ٮ�M��r���W�_<( �2��=���H��'��f�Р����J�bA�%�D8׻kX����PC����gӁ"S=w�����}��u�_�Ϛ/C
ځ��#�_��x���K4�y��*�k���H�k�\�	�7\�ѣ����n��o���~�/�,׸����_!>�k�n�>y�#ݸ�d��Ǡ���>R��q]�T��0Zu��֐�j>5�'{�Ҵ���Z���45��:��߶T�%Cj�������{Z�J-��;JsN�d_7C����$�;�='F��G0� ���;��o_���^k�3��,^�H*�k�򿁣��?�t�os��'��,��[��ѽ��Lݩ�y)ڦg�=M61�L^B[�m2�ޡ�͢�
r��Xv��{f��z�N)cK���P��K}"Dx��K�Jqo4�x�T�F��B���>�� ��\I�c��t}»Pv�\��z����t�tfJ?.!�L�	U��j�xq���ׂ�W��/�}D�'�n�+c<�2��p�sE�������ω:6�����aVu�1�K��nG��0�l�ǎ��m���okn� �﷟�Zt~�����"+�
�!�z�y��7����nd�����Y�R<�B���X{�r��I^Kq�"{T1��=Ϥm/>2I��L���Y�FJ$����%�_��t�����T�����>��,�Eșx�ᕩ[ 9�x
o�bT���w�3�������]L�0�[ޒ��:�ۉ������_K�xۓ{�N%�c�l��ݥ��IRgp��ELuJ���G����I���i��(�M+kGE��FB��fۂ*f�AB�+�u�C�,�bM"�Kua5|�ȓ�Q�z������(��]�P�	�r"�)�_�1�G4.�����Vʝ�]?//5N���}_I>}�:������u{{���"�h�ʦ���P2(]/�E��Z���ZG���Τxn{;Τ��G�k
�8�ǘ*�T&�tޖ�e���ы���\���@������D�QL�^�+x����gř��-��1�Ek�Dڭ�62"�4�S�gLX��H��nmi\_�ɚ6�!*W*��P�н���e��Ym/;V�B}�V���"�ڝ�՚�����~=����w��+�R�g����F:�lK]��(C�3��/c��do�*Ez֮ED���Xz�tڜ��5�t/ 3�X)8����z�T��K�5�R���Q�X)RA�`>rL��5uM�����J��3�2}�U��TK���~vbD%8(wל.t�M��\h>���B�E�RV:N�c�ņ��oF�OCƖr
e�GH�^�L��b[=�fi�k1�qࡐ�Q���f�@ڋ�A&�����3d�9�g�(4��a0+m�`ܵ ���i���2�h�Ա?@�晖����WG�μW�d-Q'�c �r��l%�[��*]R
㜸�q�-�3/��|�܃�F�BI��@qה��Y�.�����Ev�1O�4��σ'��x-YbxU`��?꿎�c��\�|6�R_W,�Xċ3(o\,A�LY�!�B ��O���{P�����AK��x���|�4�����l�)d�u�@��ޖfF�0s��������=�X�F��E��u}~�B������(��5��QމBj�;O����jAB�h�,P��}�XN�7[r��a���f�?i�$u6XN�0�m�D\��<��_�R�w	G�o�i�f��P�ZM]1�_���$3�����Ti�e|�(t0-�ۘn� �(!BB���`�rA��*t�:��g��b#l� ���s>�I������X}�YH[A@̖N3��'5��w�߸x>�3�Fw�Ϧm�x*�p��-�s+�~e4V嘋4v��z�h�����R���e`Q�>�PӋ!�
�O����$������}����3k�VGF� I�`m����F�㠯�Ѩ����ʸ%�lT2�N|q�������T����t��r�c��K-�;��,$%�HMƑ��o�82��s������KK)�ݪ��4����]��m��,�k�@ ;�|�n�e�p���+�7ΊO�fU��J���]Fhӝ�Y`�'k�'6�f[�+^(w3~�X�����[h�c28ޯU�f�h�m�� ���<�]o�
��-���ے`"o]���[I!�x%['ОRR;kv."��@���r$J��+v��c�8(xhpc+u���cf����y(VT�:�Ί�5b���ktnv���^�g9o��F[}Ľ�#���]RW��.4�P;�y�{��RO��W�8�B��P���Jg��rP������>�7A�W)je�}!�
�֕t�{�U�	S�q������}}�;;���C_����Fnh+7���q�g��w��h�f�Q��B��l�oVsfI�E�u�r���*�#��pU���p��v9��v��_��,�k�O�gΊ�h���`P����`}wB!�(�p� ���y*����� ʑ�*��N�'��XiU��f	DW<�ޚ�����i�!��ڦ�q�&R*�:��y,M���6��1�]G����e]ei���u�z�Z`�K=G�"[����T;W(� |�����_$50ɇ�zm�(��;q`���|<}�9�tn/)���|���R|ovk�M�3Bt{0%:��ˑ�>�;v£�Fh�UV˽��)t��x�f��U�O�%k)�
܈����{3���ҏ����Ԝ5�?R��2���[�r�Qj��(.�4˓�Xv?�o��pk�Φ�F�����n�ՊEX���޻�ez"`m%,�a��b5<����<�1�\ONDw2a�L��"C�=��n�������P8��>>�?�򐽐Ҙ��#X`7�X%�h�b�:i�^�q�h~0�n�F�̔73�N���XwI�V�n��6��� ��Jp��"�8�e=�%;��o����; �r��`a�����K�
�~=��s���m��M'�[)]��:�1��04��c�c�x�*#P���(P�N�e4��;?n%7�����T[�m�65�bNT痠�唫Z��-.�S���X��22���Ւ�:I��%���g�'�Ʀ��K�^Ʋb�nf)mӔ���Rb�q�RX+����G��s�@4ٻk��!u�6%����q�~4f�H�`�fUuJ���,DZ���2��s]����
��롵�ڍ>��tY�Ӂd���[���#Җ�y��p��B#~A�)�ǩ����5�O-������&�»�[Y�����Ƚ��8���x�\�O���h���?"@8�7��(Ne�7>G����Ǥ����>��NF�B�����a��E|�Хcg�?�xJN3�B��j�z�tե��C�E�O�6��s�[�0<q'��D[�N���t�>�C�*}鸪I��&;��$�Y֥O�z!:�]%��''8���VT�����іߞ��%�P'}�S�e�2�:¬\��6���z�%�"�U)^���2<������xu�^����EmE]�eaD�~��v.�R����r�@��A�����7�'Aj+�},���u��F��_Le+?��nb7�h�wиYo�����c�9^���pa7�'`ҿ>N���SW.�lgĉ�v�Q���Ϗ�������m�#F�<�poe�����00t��8�
���No}�,!lH2�@��
!u���r{��QG^t�p��,#C�7����@P�n�����J�ڍ��@X�4hk���!����dqi�Z��M��Ym�*�����(�����i���I��Iw-��M��a��X��3�l�J�՟����R�╂�@"���+��D;m����ʳfQ�� �U'��d�{՟l��bY����b2^]���C�"<��t��Ic�GލJ��o�c��%7P[��|I��0|։��}	t<wK����:�X����P7��a��_�U�lS~��L�J��@ތ���_r�Ȓ�U�C����C2�$ooQ�J'�:�dT��^���������� �5�1�l��4D%��3�ѭ���=!���,f��?͕�E�3VԼ��y�{] ڍ~.9��4�ggsK�紶���'���?��%�7����) �MK9w6s^���i���ܺТ+#�љ�l� ��.[�0|b�zP��$��=��82咯L�%�o���{:���k���F|e%�[ �S�q>&)�`t-�CS�v:sI�z(C$��z�h��>��q�о�����PFzs:��ܑ�g7�$(d+�Ҁ��@>�C�!�����c�f��ˇ: ��N�:����eP�����$�_O�٪��r��l ��[i��q�ٗ)D���w��W�������^�n?�.'�������|;����' g��LrH��=�¼ ��C�����z��?��WW�V��ti������U4�7}ޒ��:f��|����W��x�����,��3(����>5�;�7. �Lȿ
�Okn�ň>��YÜ��v?���\am:qe6�yX�[��xy{�����]�{_t�⯟i�t��+9��>Mn��	��������<4vJq�߬$2�@Fش�xL������&���<�����Љ��
�~��#�Yk�#���/))��|!M
�~� ��3�E��%H�������FC�Z�_�&�z
�u�k4�)�H�&3�!\��ۇ;_4�\zGB[�����T5)�]Y��P�̢P�,=?y�j���f���q�[�ŵI�ૐ�{�B�PÍ)C$.���s1h0��W��D���'��!�CCun�3���򤌭���S$67E�>�2v�����6�a�;]��0��{�mi��L��@�,O��2G��&O����P���hÈ�_�rk���j|���w:3=��Gz\�3?�}��pHKy��"�{�ėZ��\��w�2dv�Q��t����8#��8o�fq+Gg�^�^jZ�b{rό�\r��޼�N��Zy</���D�Mf����������Z]wXB�W���=.�1�_�m��,�4<ӂ��x�-V����E��*�p�$���ˍݖq�O�kN�γds:��K��-�Q�N��v1	erk��1ȷ����iP@)�W�代�Q��a��5�iW�f�eX�����SD<Y�C��CGG�*�#��W���le��"���� 03�&���Vi���LLg*��}{ć2�P"	8XIo&V��K�U�
���\����^h�"�sK{�6����N�pH#/��HK��;���wc	Nh
��>�T9`�f�tC+`B��8�{��Z�T_�2�p3�pe�y��}���I�ҳ��xuuy��H��V�J�/�lC�����ޏہ1y�䭂 n�JC ]Vx{�ъ�s��e61QE�q%���]|���Qo����H/��f]�(#>ƍn=.�B�`%���m�7o��U�z���yP�|�}C�}}Q�[��L�z���#�+�z�c?]؅(��M��)Ѧ�+	�c����eM�p����\���m�c������8�:���������+�,65�(��G����Ծ��7��χz�¨l�Z���֕������4;���@Z�F7
�P�G��阢�Iof�4|���k4�q9ܼR4_!a�=�e^��q���si����-:���Uq�&N�ח�d��%.��1M�3�c<ɸJ.�`V'����[����1>=�6�ڵ^�y| ��y'?��eh����vnI	�������1�j�2�Gi2����d��z^��6����ˁ��;L�,����I@(�����z�{s�$�#�0�G��( %�L��~&�:5 �f1�?b�)+�܃���W-c{�.hKۊc��R�r�_���jc�������o�>U%n��Z��C&e5ns3L��K��3h��YQ�����*j�,���^?w��*@*-r��"�c�
�u��m�ٌ+u�B��{r}��̕�+��%+κ�imT���̏3iQ��P���?�Km��)z�ޔ���*j&��"1���+ Yɲ�\��Hg}�Pg^g������;�O�=6ַ���'g��=ˡ��F�k{w<�7(�{������2
��Rމ�� 1�o�x�!۴�̙�aҦ|vR�Y�3V*���G�����GB�������݈W'�=FJ�1��>���܌����#� �opr���?�IKY��a�Y��V��8HΕP�<�6b��y�w����1�U�&poN�}V�?��y��Zf�1O?���HvhG���{�����63�"���V^�_43���\�l�M/TC絪"dװ���)�΁��MXEe��e��[�V��a˩�Rs����=������7��}i�s�v��MY�ܔ���)#{7,l �:�8��Ɗ6,Zf�ۨ�JTX�s����D�o�&����d��Z��\�[͛�l\(��V�HT�r��?�q\��[��x�9�r�/�g�b�̛1��b9U_���IX���n�d�߸��
8�,{)9�MP�#�s�+�5����<b @=(�+f���}t��A�}��տ�|�%]w���=e{�p+�%�o �@�ur��l ��M����Ke
q��^�$��Z���{�|y�io�Q�fP��Ñ��(���8��doa)a<�Ec�T�O�
DU��v��%�G+.�O��0�
mm7�c�cY��X�.�'��
��(�o��e�JCǢ�2�v5x�s��'��׻-"^x��-�$
��(�=u_3��eW�j��&���y}l'�v���:�=S�$��x�����������s�f��ے���A�O��<Mº�W�ܒʣ	��t��Ӵ+��3�-����B
wcc��Z�X$��q��oE�ʂj"�r��瀥Y�B�,q��w!W�G��D��<>Jb �d��s#1u˭q_f��G�V�L%$��L����,ZWw���	"Y�����o�n��٨CA��VDX��a�e&�}��|�:��	�ʓQ����y�XПwr�,Gꭊ%Y�4�
�3�/mX��r���ߜk���<#�uT*�v0��g8/�s���o�����n�VB����E��R�`|�$轤b��SGi@�Q^|�+��6Y? ����7(Ԋ��=��W�rpp�c~����]}��"�[��<��K{��.A�;L`{P� �Ҏ� �C��r�C�a�u$�tm����AA����H�g�`WӮ�FI���
>���K��y~1�=���S����M�-�bYמ����x�Ϥ���(,�?~���=���>�g�r���X�4�b��rV�5ߕT�n���l鏔6e'�f,A�1�1���R٭���M�6*�����y�G�$�G�֜��a�/U��i����D�m��-ɖi�dHgW�ˢ�6T�tj�'��C��xez�}����F�+ҹRW�
sp���Tm�������r�߇S@Yo��v�� B���W�`��d<�'������^��M�����ML��a:9)����e��t+�ļ���>�w)��JI������7�p](�_ (Δp%���G}��[|�O�H�ؠ��4����PS�2�˭����{G�!X! ��&��/d�����c{0��L�T����%���U8��w5Ɩ.�2��g%��?>��=m$aU�^�D�8�VO�~�M8I^�W�����.U,8��x�y�o�������d���Zt�vr�{�U$�?|�맞t��)�"!㰔���j�H�s��G2Ҋ'3� M��VI�=$��7��W6G�`�`�/4lr�>j��*w�a�O�i��ڹ�#���w����Ty�~dNN� o��O?��� �X_�x��Y�7�C�k{���%�(���bx'l��_l���U�D�9��	�~��u^���7�.�ֶq�"M=�.P�60�j;?�9��-ض8�2}��D1G�(䷼��]�M����,����k��~|R+FdI�3��z��Hf��(���S��;��B�����A�9S2*�R"�ȏ�V���irl������x���|M)�4�H������z؉��Z26b��u(�H~�e�u��Oo����T��HoD�n��{~^|��4��y�_�I?�'�.��_~a#�ۅ�����'��}�xϙ���:y�������;�v��]2����;U��v�G7)�_4����!��eq�e[�2�i��#�0vJbt��@%�P��������g�J���f��� л�;��Zr��jٲ�܎?�=��~3��	�s4C9(�;$I�=�˔�g`����ȖXj�y�q� ��{�b�xtoך�FH=_4Ё��&�@�fk�tޅ�׾7*eէpn� $]3�:����(T� ��r��F�4S����b�qy[!ן�/t4 �"���1�����40kП�a0�hZ7&k��7��{�X�ݔ<�J�	�@x�m�s���dҮ
�.�z��F��$���y���r�1p~TP�+2�A,(����Q|UV(��y��I_���2ʿ�2���V tQBZ�2�?A�v���_-�ѩ:'�$J��&��|�{���@�y���@N(��\���p��� B���W.;U����<��~�z�*��o�A_����]�Gކ��*�=tSsho��6�M�Ǳ;"x�d6)�{���NW�g�_66��l�+���I��Y�����<�;�~�l��<uu+�u�AH�����@��Ʌs�V�v	��/YĮ��[�-DRܦ����l���8Q��%��um�Ջ�����I��[����5S9�,�l%n�ċ�}����}}�8`3��<��>�J:���-��>��� �(��̷�ya����n���t�6�Uj�$ß�P;�L.�?����̠I��u(�S�"����$4X�ɧ�h��k�n�Dä��,f��& )Q_d3����E���w�R2���>*t��륷�=�������Nzڋ0��T��v5,���'���� @����|�ʒQ�yR=��G��m�g;Or��Y ���PZ�jf�b��3 ޡU�����W��Fc�J���X;:9�S�H�Z��w�6��ꁽ촮�pD3�Wx:Q�%�޼6�yЮ\a��.������kLL{ˇ�+f�O��IK�	*o�΂�w�Ν���Y��Q,;l�����MC�@��<Mߚqo*I�\ϑ��.jG#�ʗx��6Q������Y�f�����n��>|�'[���2�m�c�|}}v��e���}EE�cҙ�j.��a25�e�*U�9 �ku=%n�ZdŬ��:��?ϙ���̄�V��|g5��B�k4��lnI�I��X0��F$.�})I$or�9�f.�Z���do l^���:��_��r�r$k���wյ�Ϟ{h�G&Q(;�����#g1.nRU�S������t��1��>c�"�к�$R��0�c����m���%����O�t����e�\ğ��3(H�Ͻ����h1	fM��ڣ��<�� ��<&n��N^��1�S ��F�><'���pN��]�D��^X��*�*U+����	G�l�lmgI�,��'��@>S��h(!�;@������0?�i��{I����~��Sk�������1.	Z��+���P�����n��^^�ǌ�U�U�|)�d��P�7���l�B8k�~���I� ����D�*�s���{�J;�<��e[L	�͊�6�Uy�y��cc��v�H�2&�،�<�p���qlͷ�*&y��r�pVh��M�f{�UIu���;�ե:�$�b'�	w����WZƒ'(�JH+Y�S�d)�4���%���q^!�E����	؏�,敦����Zrc��ފ�^�d��ulb���a�n2צ��Z����e�x�@�mY�Y��8���u�uk'7.� ����I�鉳�p[���h]��2�Do�5�������fC_�cB��ŵ��unԂ��?W�>G���#�r����߱�)�й_�{�
�5U�E��ڄ�W43�W� ��rF�=��W` �O"�@��cr'��}��m߾^C!��9��c!f�9^��?�z!Ӎ���/R�#��&;"���O����d����6ʷ�w�2�O�+ՌQ�ے.	1�㉓�
�IQH�������9�7a�3�C`=7!PYI�? y��X~���z/�Q5o��v���ט�Yl]F-|��.������y ��tw�`�-6+ΐ.��H_̦���_�4��y�j�=g�t�̸�u&��摟���m�s��N)��ڏ�E��i9�]�����7���[��m_]8����f���:�J" �t��I)����9K�;F�>���|��!�L�A���L���B�_Čȋ�������gA��|�A�ĐI�鄰��y�隘��Z���;C��n�U��qH@���/�������V�jx�����6��(y}���(1&-�����=s�>t���;W��&B�(��i�V� \M'9.Wd6�� �J=�\��@і��؎���0K�T9D���W���?�i~htŚ�jӣ~���a9�tFA䔬
��I��J�o��rK��'��.�o4��a��j�+?���p\�73��Y>!��3'B�%l�^w �;�Y�t�o�jd�V�o:���0�"�i��C������y<��ŭ�a���婹��M@jՃ��X]	:ϒ��!����h�g5�I¯���G M��Ln��g��C�M5����{G�� vl_��B�m��z��҆��|�p��ν�gh�}΁9Rmv.��������u�cg�e���@�	��D���bO_DΏ���>��h-{,Yx{���8��e�=jyl(8�d,���:���ӛ"�#�2��U���>���L�d���-��Z{�I�������5��?"$��Kk
T1���0���&����U����d)���j"��\�A���� L9��+���7���ݻ$l����l ]�xz��U�f�+֗�k=
7��3GT��)�r��NW����Z3�=��om2�n��W8����}w�t���)��Ǜ�	l-��Ϻ�oo���H�+����,
^[�き3\�� ����쐑$�	���.�<ܕ��ſ�zE��G6aO����=�	��򾂘�/+Ң�3�Y�� �;(iw����ٱ�
s����&1�Rj3������h1��~a�{��Fw��l1�j��:��iT����"�F����ȇ��; �J�n`U���ѕP���������i��w���0���$� p�f.25�qj@�i���2O��ii:?6o��&��oƨ�X��?�) �m�,e����c��r��ܑw��`��~lk�P���i����1&�?(�f�sG�t[A��h�� 2TGO򗗯�O������
��^�z���9���t�u�t�%��E��jgy��W\�Ayһ�������Φ��D{�_J�ac�+(�=�tu���j�j/۳�	G��G�F"Ej�:�欂��?I��7s�q[(��F����	7Ta�������b$Pҭ�����͇ȉ�oZ	q��{UT�{�[uͪ[�P%>�O� ��s]��H����L!��DWIB�¢Gd����)���M�� ��R�%��ӧ��R:�Hd���ףTf���;C�ޔ��K��>(EJ\�Yd3�?{��-t�(\ �������B)
�w��Ͱ�Z<�	��}�FI�����0˴���鹒?���'�ȷ"���ъ���6ѻ�s������g��`i�D��J_�@#, �5�9��_��W��'�!*���msba�΁�'���Y{Vȷ�H��"�P��?3���» �;���͒�Iњk<�d�m��]��e�F���tn�t�e�{�+V~%%{�,~�[lR�����Wm�
4������@HOB4)dwh��l��p=Tn��ŗp��W=�����1.��9���m�5�% �ˁc����WT©���q�1I�ܓ��+�`��x��Nt�[E�n8X��L&��m��KTjr��4t�Zr��@��6���&)�$�oHj�9$D��0���q��47�K�Y��`̟����nV�y���Z�xE�d���X�!B����t
j���!�:];���qV�V��KCqQ�+��5���!��Hv�t�ܭ�G�|��G*��h�Y�P�>�e�z}ҬK����ь[��X�-@�	!�S+���
�N�H#�8P�g�h��S�!`m�R������.�u7'��o�����5룽&����j�6m��,��4�$�	�	]��v�#���co��y�X��8)��Q��ͱ�V�(8vt�h�H���� ���f%���3vP˺�ZsH�ͥ(TT��.�à_��LW�G�F�צom��#Ak�N�L�c��\7�\4�t~���h�^��}��T����䛽1����3l� �ͪG7�	��O�E���#Кm�Y��I����(wJ��Q� k:�εe塉�m��y�/��<��Dr<���%���m��4���ݑ��W��,],��`(���1�$w�q��.g�p;tt����N�D�扯�tI�3�����?��7S�P��+r�2�v�ы����C�np�A��r:�z����U۠��W~�t�y<t6HF���"�A�
u�1�j��5;w�To���QI.QU'���G�F�%��b�9�ޙ��`1e�d�A��בf�^���ý5�ڤ�ۯ��K�0~�d.�h��|g�j�ǉm~,l\8�Y�(�٫N)\� k�hԅ1ro�7u��l!��}�-M3�y���i���H�2r�m�L���z*��a�/�GrC�����Ƹ<��VG�S���bB�qE
�����ѣ����B�TsȐG&�\�/�vڊ�&����6���Fr�qD��{Ȟ+��<rD��:B�MW��Gcޅ��A4�=�g� Y���~�J��q�F�>��U0����Y2�BF0�/�l>��0n,�"��Y«R�r�d�N�S�r����x_��dIU5#7o�f{��Ob^�{&շ:oF#����:�����gE�s�P�K�����1��G���J<_��bU�-nc#=�P�"����i����Y�|cu<�\*�1o�TE+�H�w0k{1}���_?�QH|��+��������cz��-�A�.��MV����6a��h#�@�H�x���)\����W0�����#^|7	����-C��z��r�j�Inu��| �O�S��Q�I�f�#������C��x���g�MJS �y4�lv�q"WJ�3�O�gÆ�8�l��թ-�C75�Ex|��XV�M�y��A��_׍�/�"*����������w;E���Q %Q3���售;���_W6R���4�V��R\�U�ܳT�D�Q��SH*ܝY]~,��`&��gDVL7�y�\x�ԏ�a3CG��
ۏ�7iZ��J�Z��h赪�?�B��J��#��z�xz��ZӠ�0�ϓ!Z�K���p����զ�8�{�ybrV ����P���P��b#�΍��|�C=��+�G��nN%<�:D �uv/O�YK��o�L�5�����@��HE�y�Q�B��F��{⾂ګ�Z����������K`4ڕ���K�p9A�{��h����@5W&bDT���5>#co��H��/}}�C�L��s����j���Zɹd�Nl>�*�.���L�������j�����R!9q��̀Q;���.C��)��!5Z儬8%E��A���玕ĕ�/���W�g��]��S��������W�6n.�}#1�%�ك���H��n�G�����W���~�p�s6�Q��e�*�����㍶^���*D��M�7׎7��=�Z��;u��!������Y���
�o��v��)��W�8�8�\��+F�%5�^2pE�w�>~sg>׾���B��F7*����\c�இ?��iBt.��;�L��jm�_/�$�м���H��$ ;�K6r�JN��2G��X�*�߬���Ua�,�w� kh�Z|nr�� �\���O=tT���v��#��u� ��8�2�٩���T	|o�s}Y��A�3�,|�t~"uwEySr��Vru��.��U�(�E�C�L��^itb"�a�&���_9(LY)�Jja~Q7��h�LA�5nzMȑ�����w7Q��2��ϖt�P+���W3i5�=�E�_#<xB�R���~��{��9�c�lS4���Ta�띾1�����>��O�U��R�19%�59� xVw�~U���oK]����
���tI/�F}��I�t�d�DQ��d������e_/�h�g������5�&�u=)��|9+K����W���ێ�j���[�#�h��o	@�o�cb��*�^d��w���P3��[J�V�[�`��,�c?o�� �|���z�)E���}�~�R�*۵����������悵��gV��4XR�y�ߒ�W�E �>$4��/��n*�j�ju<�� ��ޙI*���vuy=�9���I�,o��{ĝ���xuz�b�PBic N�H�=�n���7I� ���R�D�<��ý������t �xħ�����Ĺ��f.pH����A=s��ⷯ�S�))��P������MM%��ˮ�{P,dT3�n���l�b�������N���H�ʌ�>�0��4V=J�-p��Q����R�z�&��/Zݻ!E��'����p-w���a7�Ǚ�V�#���;�>�MvS��_�6����*Y�8Ae�#%�yN�F��|�1���ԖH�'�ퟄ}����iCKr����ԥ"��M3��H!ZQ�o1��r@Fi�i�'�|Σ��l��q���	�[��ׅ��I�C��M����è�~�
��u���e�쫭�#l��9v��3���vQ|��|@)�g\g�'\��%�:�+I�k��O�Ճ�Y!�W�W^^yu�Ru�P����'{��F�5��	6�]s�d����
���l��;�>���&Qچ|}!���ڳ����o�w��4��C��Bv��T��l���6��n��wՕ��\�����y�2�`������oX��uG.q�y�����0U�@�N��'w�V��YsFm��կV]K8����Ї�W�\�_Dn�Jrop�2j7�O �\�Y0@V�g�����F����#��u.�,P��/�={��>=zQ�S�Dѣ��/;w4P��}v1 sCt-?�	����k*:ή�ם����ftk<9v5a7�TΥo?QEWv��J|��c��c$�d��m�VN���?�����µ�X�Td�,���>ӈy� '���x,[�����s�����g�(�,-g���Tp����_����᷹���wy����h�������]�Jt{� \tY�2^�2����s(
����
��c��*�W�)���ս�3�:��*WR�j�@��+�e�w�y�!��*��s�*�'��/�8X^�J��x�@��X�ʂyW.�V��ɡ�'���v����{�uC���..)�G �-�6���L죮�q�Ch�Y����(��V�}��@���pב�>��\�m���1y��H���"^Re���F�O��<�cS|/Pv����h1_����|T9�݄�łA�q�~�},$H��aS������3>W�Ǡw���������=P�.��	���P��|����(�g��)���j~����^ڬ�����#����;ys���#��>�!%?����x��d�y����#�3�.�!Z�8O�����Ir��j�TJ�Г:�`�������d�yߑ �����RT�Ĕk��邼�c7zY�܄*٥z�fN{����X-��Xo�o� �E3�eٻ�ڷ��Y Z����g�R�@��Q��Lr[�'V�D:�o����\|��v@O��[�a���-����{�?��g' �P�/��型�k���A��v�1��<$���f��f}��p:՚��Y6|C�|w�Px��"d�k礦�� ��j���}��!a�H��r+]	��5\����#/���h?�GY�@���i�]&���{,�S��7,d�ro�@��b�~���SG�BW ��ޭ�Z+�䳒���g^�9ҁ�	�\�j�Ę�$Q���!|	Q<�@[��'|0w Uޯ%���?������eW4r�!�c���8C��Lv���/ў����J�3���B��M��M��>~������2
Y-ǬK�����/�����B�}O]r�<�Z�,�A9��j�"p�	S��f�5�d�+���G�<�g����$z2�����#9�O4JA����N���5w7�\[�xO����b�m��L�Z���=۴�M �́���W�܂u�qV����喧9�ʝX�M*۹�2n.Ff՗���dY}����Akr��F%D �5g�D#M�0�Nc(Wb,�Q��Suu�6W��$��v���y�~��b�z d��b��V��F�`'�3�Ler���}�@�˵M��t�+Oa���K=h�8P&�nQ����¯��[̇燼�����v?�⧎�������.r٪#3�	�`����_��fK}�*�D�ؚ�Z��`8��6�����۾ �_Ӵ����d��X�@�f��W`�ڍEA����	�b(C�	Q'Q�ּ}I�����M�y�]+�^��|ɦ�D��c����7Hy�.��!����/�mК�g�)[8���Uʾ<X�C��ٹ��Yh�Z�6�������(

�"M�Ti� H@A T��U:�N�MQ��Ti�K�t	%*R��Б^B'%���꽿?��`-Vr�̞����g��7�dM�F�ٛ�x�a=����JX�;v�"}�)�1�q�}���7R���� ���1Wf6gX��s��̬�������������F֯�h
D.0Y*�(����H�;� �[�!�"Wf���#ǰ��7b��@�\����C#ˠ�z����_[���#��˄�f�����M"|Y'i��f���~H��rY;�v#uN�g�;��{:i�O%�@�O`S�/�A���:I�j�[��ԍd�ەtC5\��em���	���׷৿� V1��2�@�\�w5�%)�7��ǵ�.L��t!�d��Md�A/�y�my��tM^���z�غYH��&<�Rǥ�O������=�Z)�'+���V��]���_"����p��ّ���7dA���I���{8�	M��#���e�4�D�H]Ha�?�	} ��s����KN�m2��C�o8��e����IM�
����s��d�f_����8Y�����TC�64K����3a���
M�x�{�¸ϫ��Kq�[`+�e�*xL (l���\�<��¹ύ���c���Y��Cl���8�)��2���n�Z�ل�OV`7ֵ�#�%�:K�}D��o������?�����f���?�v�Ԛ�lXXL؂�"��M�M*QV�C���sv�
ù���������̰͡�Xj3N���:�눽��� |5�]��kcS�0Jk���G��R4�@�&43�,w��ǁ��H74�ݪ_II%�~��D���֫V��I��#Z��v���?ޙT|(X\�a�h�tPL��O�p�ϒd_����|H��IL�����~�1sqq.Ka�w�
�?�-���_G_�-���;��z)�����Dw/��<��2ui���s���F�`A"5�Z$��軇[*F�u��U���'�Y���$�����۞A�7���W��E�5S۟�HD����1U�2
��3z�<�ܣ�+�"�%��؝��0�R!�!*w5���-���D�H�|�m�C��g����f��+�;�+#�Ko�;��9��W(R�7�|��L�'���~����V~�Go�;B���w�o97�r_�V����Xb-�F%.Q���Ԙe:h����t��.�������F�mY ?�7�����9��������]��{�G�L4��xӄ?ޡ�#����HXL�ʃ��"�|�{s|	��<���|��2�p�A;��J��?���YU�t�f���m"�~_�ܣ��yƞ]X"v�I���&�{B�D.t(~J[,Q�9��3��]��˯�I�_�n�'���￥�A����i�1Js���>}:�J�w+��1���vA���/]ߝ�\^�Ѵm����$E�3 �JE#F	޵�G���#�$�ۃ�����v�
Y珞��C�.�0��R`4b��Ai�?[��қGR
3IXҙnF>T@ kh��-!�s9W�ʂ���nj;�B��гZ�b�6387�}��ɥ�]g��\���5T� ������k���}�3�뉉7�CAlla�~:��>����9��I�
����H��|FM���+�y ���vF�����G�z�Ҫ*r{���d�j���ۮVј�͟SA��'=\H� ����)�/>�dh� L\�pyφ�R�F^{���=}��U�d��L	����Z�<"A�^�����%�KaT�3RrMҽ-�Q:7�u��0d�&#��>|�g",�J�QH��$���j��|&?N;�l�8�l��BmdݨC�9���e��L�=���.����
׬h���z�1p�b�^�*�TEI�z���(�����]�����Sa&��?:"j�S~z���^Lq�����f�V$��-@V��o��:6���IUٮ&�l�Χxo.�,g.��KJ)YWNZR{�g���ݚ���K����0-˷�S��#���]��>�~r�s���d�O@0J��ʧ)����E���P�(ߎ�����ƚ9�\d;1>��U����7�-#V*k����@]�6��J�� �k�b�?z������@�˕
��(��BCyyv�v<\�;3SCR㖚T���*��d�W�^�a,|���6��|�!~�Կ#Hp�y2Ы�]�N��[Q�މt�����������n����.F��M���Gj��~�����rp`����Yf�e�+)H)2�+�cֺ����	ɹ"��,�'U�ń�	���K�bRR껬�T�3�3�!��9�=�"#��J�Ѿ��gA~�� ��h��&Zo&NvS�8��{f)�c�"�m����xd�;u�*�ZUo&LAc��sZPU�k�ի8��U�/��e�k.��#�-}SO��I�+�H�<+���?*�E�ja��&|����>R(��@����/�
��M��G�bT��a�1
xG������a\�;{B����-��T��`��Z�.���l!R��i}\DXM���O^���|�G�Ÿ�z�K\�����׶ Y���U�Y<���X��}K�o��{�nNϑS���R� ��ð��*M2�����G�>1/t�D�����5n��8��d�C�ߩut��}���u�r��(���ETu��QX��>r����̹��������eZ�y���l}ڡ q�6���X\J�N�E��%�;q����)Ŵ��U�ai��Ѳ,ң��Ri_9��׀}?�49
L��I~
J���j�B@�X>��| �MVē:�e����:Q ���TAP�ſ�(�@)0A�3TFhb*�w��T"2Ê��F�@ %����k��j�c��pw������]��T�p�k������\D�!��e��3�J�/>���,I�����V����V�����s.N
�~�^�K����:��$�d\�{ Ѱ^�Wp��35�	��n�6����I@�1��[wZ'&l��
�i��R�#��I���
��}���H�Ns��f�P�M�T��})�9���6��<6����PI�+��ґ���t!V�7�q���b�[�9b�
p�W��0	5�4��(V3Ы��c�L��ǩ@B��J��HS�b��+�`����rGzu�Ao�����EV�[���ڱ���8`nD�JJ2q!���h��06���!{>��C8�Й�%�#z�m��WuL�rn$���7C-_,�y�_���ٟ}�,h(�ޡJ�D��$K�b1���
��� ��8��k�ٳT:_�R����=���Ǖ��ҩ�3):G"5��>{�b��D��^g0P0�ʩwE��6j�vo.����__]�ӗ�� ����_�)h���������f_z�ˬ#B��w����_�V�F��׻~Nx
���~�:��]ӓc�5�ܬ��_�רl�3v0��m[z�c�յ\t#��2A������.(}�{Ar�W`�.m�f#��8|5i�؈�	fP��h�?g5���[�n����}L��Q��>q"�oOl{Y�6iW M�n������[�Sn&<�����0�,(�w�K�"�!�k_^����%�����xj>�8����)*��Ŏ�!>ViF�a���8҃����'C݅~�#�AF�hP��B?�*/��d���x�$$aO�1~�Ƽ�5P��ݺ[����&�>�?!���߉��)�ڛ��S.d���e��]T���1�a�EZ���ڀ8�/�R��Uv��f_������&q���scc�FL\��W&9��+�`Z���}�?�[����5�F��p��9����=]�Zx_>�c�H�L����Q���zd�N��]J�����kO�GYa)��%W�^���0eE��Mq�s���?�B��;��L�[��+�::�TU�C�A�t�YO嶠����1��������C��p��]�n��>++�I3�H@��#W �$���͟5{$�3��X�<%�[g�'ȳ������fe�3�Y��J�X�@C5Sr����q:��#�)�_s,$軮c�e��O��#!�OC���@~����g�F_���*�LV����O��1x8��%��5�x��٥� �x��e4��o��ɔ�E�d��2�ۅg�!�
�$}ewE�<�~�(u�ϧACU6	�
9U$��Z�2�z���`�Ե�J��ZO�-1E�9~3���e�8,�̇�4�GƷC^�\��]���"�2e\i!�cw�DXж�m���z6��+�e#�1�(���J��S�t�JU桞	����w�eV��+eb0�fϋ��t�7��.��v;~�������P��_٠�k���3|O�w��#�n��w����1�����A�3/��{7fPL*7�xO�OB�]�	��k��ǂ���Q�����~�@����?`C�#�ϡL{$����f�d�a��l����66�$;_=hgmd��p6h[�><T��+G��L��U���D��\�C'1���VK���Ң���EPT�ǔ�1ۓ�>F|��{iѪ���V�����ď.���w�<j`*΋rչnt(1J!	;��U��*u]E毪1����=����m��w��8q`u��ұ�1���3�
�֝�����=pV��G����c�B"#)讍����S1w���(8iH���=<r ��#������y}�^Br/�g �	OϨT�n�(���t9����Zd{��1}��fLWQ?�'��ExO	WZn鋫���3�k�kE�E\�C�������yI���n�k��,����cq��6�kn�j�H/\d�5~7���b�2:b�aY�C�0X�GK�2	I�y�ژGC�U�1F����wF+PMD�g�[����>�~-�+WA^�p����nm��F󊙁��qkC0zZS�/��g�q�g��m���K�����������E�az�pIp4�[�>3�ȗY�+�Kֵx z���y�Y=��K/�i�D�����ްze�R��pS�ޛs���*|�Ki��Q����Q���5B%E0�B2�z&L�^��*��r�>�o��Տ&;9��7��ʅD.���HXNTЦ�w<�!,JU�Q?;�o_��ξ�[ho�����RL��*0~Z/��v$�h�/��LK�~��y����]�]�x�������X���h��ױ[U���̚u�MJJ*���o��Q�vkyf���Dj!�(�^ږl�~q��
�O^%{��!Dcu�5u�0�s��b;rϘ�T$cs�s�q��X�i&5A��vո�.nf��)�x���׼p�������oW'(Z?�e���R�+{3��_�v�^�ug���3��9�{�ub_��s?¨���&gt�ڐ����,��D �A1�\/Z��A�G����p�j���v��q`}û,٩���$��~V��D��w�͡�)<5OC��VX@Zs k�7`���=�s�c	�F�q�)�`l���n�B�8v�X_l�!��q�,yi����܂��/Ȥ�pض�k�h��at��r/#��8ɦS���G�~$E���pU:�y��_�ՙ�Q?f:zCz4���8���%1���ߢ:����^�Y��k�2�޻���q���E�z���^��o�Y�'q�@_'`�e��+�g�̽A^�N��+�p,Q�ѸH�n'��X��o8<X�F��դj�{ p	���o��^��}9�WKry�Y�s�<�-�e̮!	��c	`(�D�*�����^Q�_��O���l�$=�]� 'LG�@MrM���a�$zQ�dڂ��'e;zb���rߐ9$S�޵�QC:YHr�H�j���\�̊�_^��I?�k܍��V^0��սp�3�j��=�3i3W��Ɩ�Y�#�T��u�����L>���ۆ���ħ P�%��G� �m}����ٽ��;P��*�f�� ��f���ւ;)6Z�5y��5ҝ����ID�?!
=��2rϑ ���A#��n�>t5Y��N�Ǯy�fU �4�� oI.�k�2����0�1�|^4�d#���M�Ď��ŷ���?\�Ν
���T�`wM÷;��c׈�n��L�F�=6�grx�b1|�X���e�:�u$Lf픿-�d:�nsx�ki�G}V�9����y]��^��̀u��ɦ���+��.�Y�n��*0#�!��xm:H��V��3��jڬ�׬�@�<PC?�x�)�G���Vv����k������a����Tr�T��m��_�[h9
܏$n��"�1�����u������zi�|-Zt7O�K�ѳ�^������w�1����LXv�\�w�6_�|�7>[mѝ6�pv��7Ǧ��O�6�h����G:Q��L�z1�l�^ppe��6�[����_I��!����wf)�Ow�*6s����:c@Q��*�pu�R�q�97T%\7��3*��k�#�K$s���M &�<��l��{��
�I��v|���J+��{~���$d����WD�Z2u��`@�2l�s����!���X��ZF$.o�<�� ��c����r�W�t�]Bq��]~��
@̩�c��2բ[c}�pL�%G&�<mX��>b��i��o�{��ìj����yI^,G��M8���fLY>��7�Y3��X��r�Y}l�6bhX�_� x�H\�v&�PRv��U�(�Ko<���R'�٤6XJˢ��tX�^��{�%��j�mP���K��~_^۔�&JJd�UÐ�{�YE�؞1�y�����{ls���`O绾[�A(��`S/w��)��0�T�5	©���d��P'�xQ/�|�qM�]��,���o햧�,?���}nUD%���� �ׅd��i�@�j������Ul�v����.�8ݹY�h5�ly������*����0�����"����ΜSm�|���\^�����e.���#z���Z��g� l_�w?Ƌ����}�_\E'����ujG[!@g�e>���y4v0�@��E�!��� ����o�"�ס���.R���"a]��i5#'sQ��@�:� ��1���S_�Ѫ���Z ?v����3��Rs{e9 ���������5�Ua�ݚ]���a�{���{�W�M�Ɇ-��Νb�x>q#�b3�DiB?j��E����������v�~��{b�2 ��"���S�)��%���C6]�^G-�V1)mTW��PO��� ��n��	�Aca2U�l��Q�]6��Q4	Ja8�+jj����Z>P���a�3�e�;��x�/���j�M��"���k��������ydՕm_L���%*rHo�O�e�/I��B�f?�7��慣��jMѶ�����1�{d�ľ��;��ם��x[����a'# ]kn�����Y<G�������栯�#ꝼyI��+<�P�*�u��J�;�e��1�,�M�P��!��`�"�����G��.��E/��Ǖ�&#�i{�⇘���l�1���7����Rj��B�<��s�*���
�iEAT�q?R5WG�J+����z�[��;��%��M){;����9�� Q��8�����8R���{j�jg�Xhx�zY�X*ird�f���f�2�݌C�txk|�eq��H�H*�K��N��ER��56ퟫ/�g3yOW�yhN3��9[FX9W��@�������.v"@0pR��P�KVR�B��#����o{d�f�^f���{���̄ ΄���`��޶z���iNqA�̨?�a>���-tZ��g+�H�h���1d�MO���SO����BCz�%�"
�I�͵��'��Wg�`����mR5F���E�M����=�	���sM3�
��z��[�Dyq�ԃD���5d�B58�N��A�h��AJk!@�V�P/g�p�3�����Q�]M��$�n����
T"Lb��&�^;�v@O���$lZ3����� �i����<8���է;�i�,���D�SS.v��
��~+.����[�U1l}��a���>L*z�T:cD��~�!!�?��)ErO&�c>zH��1�1w�W��'���l|�i�U���N%�����C ����4�i�Fa��M��s*��I�mfܨ?�I���R?�Ǎ��o��W�2T<����W�6�B����1.�)>)������j�+�8�����rt4�m��7��{#�����g��$t�ua�U��$&&[4P�|{�Ԝ�
��ExͰ�,�1��pY����~`Nq;����g3[�&!s	a����"�ړ���1:�죤�O�@��z����>�������%�����������u�L�_�֧�hy�h��)���_)�m@{T-C�1��@<���K�%�'�r_@G/��
�uSǸ���'`n��/4�Ϣ�ו9d��mw�������>��(8������5�?�^�ZЂ�~Ƥ����א&Da4	u������(�0�e#''�=�<�AL�j{s��h��������פ���:�a!����8�U�jd����2���[�>r��>��p͂m��3�Ҥ�_����g	�&:��_Bs-��8���m+A��O��� �{���hE���ʙ��S Y$7��#�T����*����Om�<��N�w�=���Oh7�**�S?��S�����h�t�u�]�ڝMd��0	��g�T�B.�|XϷ�*�-���i�f-�'�6�|���@.��~RRd�	8ۑ\�L�/�}��`��\3��3ui!��xPd)Fe��%ً�J�w`%�o)��0��O*�[���b滧#��rw(�o��x�mDe�*��V<+�Pr?<r���y	�Yf��`� Z/7�5�78b�Y��/�}���c C�j���bk��9��Sr���ߝNm��zo��-�kx�g��j�}@WI!T�^yMι9ŷ`�ҾǈO�ݼ�ǩ��ȩ�Hbe�3}�&�N�~�T��IY�I�U�.��FV��d�3��?~֟5jfP���3�}�B�t�8&��%=�L@RJd��;���bmW�L�3�?m�8�19��I'I���.s[�Ƹɹ�{[ghDwa�����\$p>��/_ɖ���{�R2��
+�v@G���a�Ԥ�{�u
���$wߙ�?.�5�tn��$Ff��"�����כ�R��R6{��%}�9���>�:ѓ<���'�����Һ�)��<t^y��Xy��|wC�RQ�Y���r�Q٢'�҅g"�o*fۆ�a�:F�o_[u�7R	:q���DF�����FOY������M���,~�M�N����4��#��)�D�?����7H߶��i�v��x��H�'������+bKy<��b� �-��=xt�w�f�݋��|�jO �d�(�J��f������$�
�6������3oa����'(�G�
1u�~Ӱҫ�_�$�g���l�8�����iO���d=�jK��\�ޟ2@�����}\�
�^��I�@�G�����4�,�����Uy�ظu@����YQ�1M�5n��|?��ܹ�w�~���Ei3�ٵ���A<���Yqjf����rTp���|!p�OM�/���s�!I��h�?⹜�Ii��5��O�g��m^�}:0��S��Wo��h�8BN�p{�."�)\�\�~�\��_�EU�_Z������ɽ$኿�]�p�y��a�uU5C���א���
��q����_<�?��|�4�fp�����6,���6���7�f���M�WI���KO�3��;�ƅ@�ZΘMS�B���G�ͧ��BTP�Bt�R�n��㮀e~�[�:Z�����S�g�ULy݃��ܢl��}�LX������o߰£["C��Xx�Ӽ�S�޶������ޜ@�qa)>��A4_�:�3Rj�"9���W����8�;�y �ሸ�dlz/�x.(xXF��$�g�����9N˫?H)�*��K*iP��=J���.�E�~�sP��2K��*,��yq�Atuw��y-���K���?���6Z6%�h�Kԍ� 0�؊2���br����;��h4����%���νtU������jV�S-�Gt�g�'xyx����sd�[������ f�@����^�Ƚ�ޱ�M�lWR��{��$]�e����,��/�L:19��u:�(M�JG��]��7�̡�	Iױc��cDm����=]�v��2�gϾޔ�/��'���Ev�$����"�͝�5
��;�j;���n�GNdQ�ǲ�}Ʌ��EFX؇��z�DWt� R��XP�ss_GwQ���|o~頮�\�r���QeĈ��g7|eu���ͪ��hrw"��$O����o�6-��9���|
#���^�'�J<!r샇�I!�۔�㵭X��\t�Z�Rn-ru��Z�PS�ֶ?�N��p@LR�+D
���V�r��F�Gj�#�~�QBOC���u�__X"�ko}��^a��ҋ3~R}�b9G"�:���Y-.�/�
���rn1��U�}��O�V��P�lHI������ia��1dN�C��4�0����ȿ+���x�1/��o�{>����n�����γ ���!�. :
���qiv��mI�cse\v����0�Z��#������]O������Uw�*���wD���>��<+�2_���8$�r����S!����6s똮�]�L�uRӉ�g��y�R���N3��*��+����\x�	e�D�.��/_D�6>�1V ����_��Vw(ex5����5�����!ھ�bX���z�æ<�����"D�^q�w�=)Uc"s�2�K ����熮�����a2Y�Y�F��ҽ�d���H�����o����<[�l���@����³R\�A�|����[f�`Пژ��3�a�_X/�훯35���lތ�7�_{��	�!�P:��ƫmz�5ޜ����ę��J3��Y��qm;�bИ��!�J�����y6]�[Əaw\N˂�}���cִWS�*��R�Fe�ROm0����A8�v
���C�S�$ڀZ��:��w#C}�]&�w}
�.��Jv�O[�G3}�y9�\А��@�r��5�.��p�)ʸ8���LG���N2J:Q��z��x��B����K�$��鋏�tg(6O�e@ժ�W[��"�nޥN'�Æ'B�%Hq��5sHFV�	�Z�r��W:���G���~���@w_���'�'��.-݇�Ws`	FwNi����mk&���s�!��T����Z�+�wJ�a��!5f�9`��L�����r1�������bLG����M	�Em��I�`mY�=\�j"M�1�=�*������'Ģ���Û�|��}3���@Ձ�X�W��۶^[^��u)r�l�>9oԢ�m�p>b[���A�z5�x��-6��Χ,����10��o97q�55���YV�����s��߿G��Z>//'�^�1����z\:F�m�F�N\w�eOZ�Eٗ��]��Ʋ���r2C��U���U�����0(���e%_�HV>�_0m�ۺ��u�ߠيR��ǩS�+�^Ʋ�3P�&��|��i٦�:��~h�D����/^X���T?�? Pz���oSNlF��XS�}[��5��IbE�[�W��ژ����*N?=����g"J��/����D|�ΡE�
�D֌�Q@{N}9>�.���,�Kh��ŧ�N�����遁2x��2H���S�~_^OF�7*���N=�ۿ���X|
y�;�470�����U�o��/6𨉖�U���Ț�)BM�9��� ��Ai(c�d���m7�P�?V6��4)��΀F�D����]���`�V��G����ccW�	�L�g~n/�9k��<(��~]QV���>�Ul^jZ����)K��c%pN��׺V�\ ��u�8�8Gg���T{mVO�o���RY�T��u�׽Ʀ�ʐ�U�P��˘N@ͅM����} {�K��z��Xj��`�ÔV�l|��{'�yWBOG+G%ǿ/�⟆q���C 2��C�f F����a�%g5�ӈh�����eK�'��g�{��V���N p�Gl1������H�e��ӗRQ����&�&�߇B����4����v�)7�ZhꞄ׹���B��V�y�n4�[4�����3E�5���z>��+���(�����A�IM���d<nޔ�_ܖv�9$nW�K�弊ԅ�!�� I	��;6e=�8� ���E�W8`��rxy��HU�WzDW���ڌfz�3�\VaS>h�(��^2b�
1�6'�I���rwܐie�1+(B�D����0t�!���q,
 �°��g�9%����%fF�ĸI����͢�I��~����3C	9j�e�1Y�kE1�I�L�)O�w�mwk�\��
b�IU�=[p�I��)���̀��?~�����ҙ�T�}�Js=3��Q��;��w��U*֝�Ɓ�5�M}�r�&�\=VT��:�G�ĪfU ����98����y���B��aWrU$�{�b�~�<���	���q��u_�ʳ��2d�za)�@�+���2d��5���A����%���a%]�2q�L��!ZT�5'��Pc�^P����pib�tǓ��y~щ��)�Xu�����=(,.k��ri���C�6��g*�����7����0U��Cbj�l�8�!���O�Ւ�MĿ���.����'[��+)<�����C���wnU���\zqt-���w Z�]����z�C����v|���X����d��Ӻ�?X c�J9K���W����Ze埠W����!f��T
�8ݕ����K�T)�(#s���,��|L��_�R���}d�yo���d��o�q�� ,	��		6��ح-�bq�Z����,e��/��o������9��LN��G�O\� ��h��������i��q��f2n���T:�q$�L�n����]����k�P�;d��Y�L��!��`�˵1�����CT�d�s�1�����ʓ��1`�pD�(�Z�}L{��S=��r���*mz�ٍ1��~
Z�LQ�.�$��\���O��-��sJ�uN�9?��B�wdjs^%�wK��u),pK�\�f;Jr�d@��%�_Oo$&s0%���7_w���)����83ߕ����᧞?�a���MD��5�[�a
�>��_3����S��P�+%Oh@5t�,�"���YT�l�ӓ�ϖ���.W�q�f���U^v@ؘ�'V�%آ
�Fx��ݘe�Fi�r�}��&L"��ah埴9C:�a����k�_HA�"R�A1�D�%�g��i/�~׏蹷�o�S�nX�X�D�DX^6Pd0�2р�����E6�'�����h}x��K�Y��|��}ã��^������S�hה,GC�h���ag72��$Q��k������W��Í�͐��~��>���t-�>��P������ͭ��b4}���`��i����H ߦozO��)%�Df"�?N?1<L}��H����?ZD���]�S���#u���w�!sCO����w���{,ɀ�8�m1e�s��] 1H�x��4�;��JRmN��-��C���.�:ZB��0+�����Ζ���}��B�z��d@|?Y .<���0X����A�����&�$���I ��Է|���Y�MW_��:���q�
Q�@��-��pW�)�=�qF��+���;mmg�+`�q�8=��U�\�f��x#+��ӆv{{�Z4Yya�����kT�(�\�n��4�Y�C�p�����ՉB�RX�.�歛�DU1���؏����
B���x���.O�ҍcz���TU�>�8���ۂ�~�n�1%}�r���R��b�-c YoîX� ��J���q�>�/����"�e���o;i�h�����t��'=��׽�{�ލ%�b@}M{���x�}�n�8�j��lGH!�]�����,M�;|�X�Dm~x�a'�#U��@�<\�ۜ�Ih����[~��3��#����l~��H�� >y�h ?7U�[�R�o̫�`��Z�_��L4ՎP_���G#�������Z��\�,o�H�4:���_v-5Z�C�>��琶A����}t�gN��ӌ����?)J`��З>ZW��j0w�L�'�Q���@yZ��hG{�<���&�:��eTG��ꄂsr2�1n��"1�U֏�go�X"�ʹ�`����1P_�
��U����̖�z��wq������q8}�ٮ�9B0��e%��C�8zs�n{j̴�v%òĀ?�綌8���z���<#� ֭�Uq(�8~���]ϳE���o4���cm��ʥ��g����X��F���ؐP����]��w��"\j8"�)\ s����-��m�b�&Ec�U*ѓt聁*�E��Y4�neEbhM��Q�V�{4��>Y�Ɓ�cX�@���Bd�zN��$���,H1%�&o�w;�Y���a�f����%������=���3p�j��(tAa!R���]�?)��O�I��K�5�!�Mt)��}@׺�k�y��Sߒ�n3^������Ϧ��(9��6�-~9�P����&P[-���#ڋ�gq�>�nx�� ?�t�j7��_���������P���0��9�6Z)����`/����	j5S� >~4��όD"���'�9�`��[�ͦ�l�
4��N��1R%������`������"*DN�b��Ӳ�9��i�*PJ����׳�.�M|J�j?Ē�+�������]�N5�w_�W	b��n���~[G�$=��N���T;l(6��v��7->���M����{XN���bW�7�!��Sl���1��1����1�m���C*#}RH�m��L�3�K6�H����UK��W���ȳD��~�>"�L���X���G�̓#�~m�ߵ��j�&��)�Їcn6&4�$��)����$��S2q��S(�p2�F�e�y�s����Ly�B��[_��<1"���P�c56���˱���=]K*vM�ln<�b�˘}|J�ϴ�R���2���9�B�|�k�Eqm֐��+�H6��=����<m4�O�9K�	��&v1�[3<�,<Q�M�ؕ5����ƶ:�˵f�YfߥpMk� ��9*���ĕq�ƺ)D"�Z��*�����S3�Kg䟾Ҥ�y	�W�1>��6X��US �z�dF�d�uQ����gΞ1xYt��I��B�+Ŵpm������r�r?�_�8��热�C"Gw��/�Û��.����<�dU��5�r#]T�����u!�X�����+�?�)����\7�(�2}�(�f��b�ɗ����"�z��9��0��%(}���z���ҙ�9���Ⱦe��ϳDh�C:�	�i���P�������=�2���|����@�c��2��r�O@��{�U�۫�,1n����
�AZ�c��-ȝ����W�̸Iee6ȼ�3VŽz���c0ETx	̘�l����a�E�d��>;;��S���#�u�x7.�0��ڿ��,M_�� �ha���t oF�kvtu?L1	���_�� �d��S��c8��>���ܵ$����&Sp����A�5��m�����Ϟ��t#��_����{5�ʅ��7Cz�qc���ݟf_���	���=�"�,�r��)
�r����qI[?�L�t"b����3��PN���{�2���»��-�o��5B=�{(4�W]�^8	5M�2ċ��˼
�k�k�U�+�WSO=�$�8�Ş��n�+3�S��}y�G@��A/#��N�2+k�s��/����Ҟ��1xᶘ�R����b�{��P�� �-\@�A�~�βZ�����AW�F�yO����ntjm1��~Q^} �����W<�ݻ�(L�Y�10�I��4��Z�p@����ۜ)XT�xx�SW�+������T���'f����
5@�1��:�[��[_#ԳT���0٘[��:���+�MM�ؙ��!J�=�2��'��a��R���Oܾ}Ҕ�ɋ1��^�M���⬘��	:Ө���΄��ζ8
�pa�OT&5yfO�
.�@�5=�#΢NU#��yH3�$���c\� ���O����T"��[m�M���~1ao�Y��^�U�`�8L�Qr"}]?�{�0��\��	�Ei�_�Ɓ�O�gy1�~��������:ޣ�_d\-���r���I�[)II�e���|��G>vc�늌�j�k g�]j��)�љG��<vy���E^м���)���k�9�����$�UḼ_��'�^�na���'���H�R�M�._+���K���t�+��x��bG���\K��g̣i��k����$�B�CN�rM�U�o��5=����$,�P���H��d���i�KJ&�8�D!�s��o�����/�L9�B�&zE��/)\_�}�L?S7	k��D��Bx~B���+��L���,��
A�zH\d�|�p'�P 9�,��,�:���'K:���;[Mn�#9����De��5��0�G���;��]���mS�p	��R�EV��u]t�����t)˨L����O��3�ŵ�W�JJ��6�n�NoL����PG�Ԭ("B Q���A�S�&@w�����;��l}٦"I�\(��ZU�eiڨ>cB~��1t��F�ͬ�k<���t$ޡ����:����3՞���R��KhZU�Ϸ��{��#6=;�=k�͊(�<���*�92]�]�uRYp-�OF�u(�^ӑ�U��lg[�N����BDp��cܧ�əe�9��"+�k�����'�Ý6H��aF�i�ن���&���q��R�"D�H���1
�I��l��8rj�Ss�6��`��]I�h� ���| Pi�j�3�G>�Ã��;W�� Ɠ
�];�rc}�����C���8J4'�4ٚ:`1%!5�|w�{v;�)�Q�x\,���£8�#vc�SAy��N��|�uXT��>�b
�)�Cw*��]0���P"�0t�e�1�#��-�;�^~?���u��pf��W��^{�����ipZþ_Q������f�@ l� �BHy�T��
~�!��`��1��5�D� ���p(�E�}�ۜD���E}��i\!=k6�"��~z'��K�w;bm��PX!xj+e��'��o����}�ُUs��s�<�I*��jf�J���^:��k�
űx��������a����hԔ����t_sd˒�!�#�oP�F����7F�X��Y�[��SB�������uW���2��U��c�ԽZ�U$óA\W�{�9��_�F��o/�&��ȁ%ډb����~���i�8�[n�x��\�|����o�މR�ղ��Z)�����t��v���nΌϛxc󚫿X�Ș��u����d����k��$r����F  ~�_fZ�I1"�on_4K�>��j\�������=��=�oAR����������4ڄ��zf�������H�%Zw�����H�g瀮݆ ��m��s��?I���$ CɟA4��!8?}���a�g'Ҩ�?v�)7_���}{Y�����w�}�~��
<Gq���9�P#�?wP��?�>#�:�Xo	�.o����5�|kM��Z��n<�' ��Ub������D�V�t��;�׬�.�q2H[����M���wW��ݖ���:�=�'�ǎ�,���*��U��:�z�D������pC� 8 ���'ׁ���Ɍ�a�a���1�.k>����uKZ�A��x@�y��7ҼCm|@q�`u �\�r�/�0�D4�����<(��,,7��+�ETԀT�[z�������j�i�䢔ȗ7��r�&A�E�}�&�!�#*��p���/RG��ev�s���A�(��^b���G����o&x��;r�4���+��@�;xL��	�ʉ��xxV�Z���~0cPa�e�"���1r,8}�:U�N'_G����^���'�E��Y"UԆ��L�͎�D�wRb�$��B�	�J�E٤��-7l���[��q��	�g��ǭ�����^g,��@��`�V��(`��6kf�N���?!��s�ch����2�*z���,���u���u��w%�gߌ�^~iAy��UM3��
�L_ނ�s*xR�>�BE��	ԩ��\�tQ�V? 鰖I�=@�t��o\@MGk��� ,Nm�{5߀�������9H70�����wsP3�%�fcz�~a�͚R(�^#�"0�M���އ6�꾍%�k>�H���5�FU���t��.� �O�sK���Q-��^Op�_��\�m��
�sh�,�)eS(t�����H|�)"p�U��|�Ϡ�r��柷IaG�~~����J˽A^�t��4�f��ZJ���{��[�59@�Bz��%��Y.�`z���� ��"9�N�(�<̟Tu,�0����ŬX<�|�\�54O���|[�9�[ګɅ)��3�Zz	=д13�L���ejo��m�cȰ�|p�}m\���Su�"y��#Um_�-X�xdd�yxG�3w�t�"$xۧ�?��*��e�F�Li��2��2���z�ϼ�O�v0��г��-;��O`��>�^�c}@*g����F��W Fv0�
W]�<z�;�*E+kl�	�9$����;?��\�Qƪ�\)k�祩M��m������E�'`�ٝ�>��d�1==0g�ȧ5��MU�y+U��G��]��{�I`d�D�5���M�
�&X��}��NLB;��b)t�j�����	,�WW?��{�{�y't�i���|Է0қ��6L6�x��j�޲%�<(�ȴqV�3w���\y������ҟ_+_�BV���D��	���`-����ҁN~���!b렋�y���'P��s?�{����W����.��0��xk�1u7�.���d�&)���O��<,��n��\����̤�XI�F�uT"����uz�7���YX
d3���z�:ǽy$u�$�{����g������ޗ����cf��H�>pz
g��0�g��1s�{P�un�A)E3ը�/�g%Qg�Є���K�^��t�J�ET�ݾ�����-�@i�4�+�f0
.����߷�Qψ�d&=���?�g�AghQ�eV���;��y0�AT�6�^�� �j��I� ��[:���<P=���K�[�ܶ������]1������ǀ�a"b	PpEq��/�T�� �2dƞH �efN���m��-�XEM,-]N��k
`�}m�bV�U���X�ca�h�6�PNǒ�X��������Y��i��JH�L��D�ekqܐW�Z��^�)��"�4��)iB^i���b6'7��Z�%'�ģ6��4���V9~%N�]�{��t͞��-�.�/ףU-L<�������0�#~j�X*<GuRt	&�z�'���tغ������u�a���y��8���l�W�H�W��\ƞ���="�y_N�C�X��߿�w��{oZ�g!��7D�y��+4O�:�G��ZE�G��?)��GN�.~��|R~פ��Eq���TP�{��"����x~ٸ�V��<��x�<ѽy#1}l�����%�	Ij�%�
�`5NשA\��Fޫ�$��h�w�B_=TQ��px�t}�h�f�����Qhq�LLo����OKb���r�-����v�\	ժ8Ȱ|m�x�Iew�]_��m&�K��&��s�8�w��M;��4��m�����)�R�b<�7��H�L*��|����a����2*��Ff��С�A*C��F���meXv��G׍v�����W�	����HK!L����O�����W#�|��ɑ�f�}���*����f`���߲��m��=�\1�i�*����V:�FIh���#�9I_}jŭG"�sv�I��Y���Y]��:
�u�S�6�ꦟ��@"X�̣�Uu���-ln>S��/�1O�[�4o�_��n�0����gSOܽ���k���B��e	D��<0�lD�C�����!�@0�Z{�*�y����@q/��WӲ�T(m�d�>|Ԓ*{��2�����ț��W���%���F哙�������݀�I�@Nʾ�=28?0穪�oqN�v�ʫ����5�������ޖ���Y]�����������2?��|��dH�Dh*|�冏��f�`^ܜ����l��O(tL�d�=�AϰW{����{(�	Ì�������2�ָ��z=�E�`�ɨi	w҆U(��n3d۶�6���C��uO4��/��(�����z���=�#������j�w�������������2�˗�TYw�ފX�pRv����J:|�U2��2�\["�[G��" �;�R�:t����0�����\+��]�+92�\|jYH}$�p�گ��{�Z�oNⴾZ�����=��pNo���9m��[ƭ�rz#�9>��w�5�i>���U��r,!�����>��(��؆B"�BP(�l���ˎk���-��m�߻@ R1������fN.��<�r�Na��P&O찪:���k��ԃ�,-^���;��<�8>�i�pX�urO��M�է�{o��ʕ��FJ$�w7��_�P#n㘯�Nϲ�1�O�	Xw�v&�����r�|�Ӭmf�	�FO�R����>�V�$-d�0���+����\p*@�sm�_'*��b�����<ڡ����Cw��'��B���5?t�#nS�k�y����6����\��Y��T�I�Z[Paʹ��Q+c�h��B~����SZ�N���(�~+\�����:*h�v�T,y�QiA����[�$�6!�R�ˌs��F��ꮔ�!�N�臷jFGWW�1�7���d�#�<�v�!K$/�o��$�I߼#�>@��YQ�n��jq7}��0�@Ϲ��uj�i�j20Zn� ��^��\��_bT`�!q}�&Ⅵ�.�P/���RՌ�ԫ�F��c�3D�N>�OaoNII��_Ҿ�-(*����s�KiE#)�J`sli���Bb�ݓt�	T9+�,S,c����"�tO؈G��E�N���`O;�H�T`#�m�����'��3Gk?�׿�D�$̥o�爚�)� u���6R�ĭz��|�-b��ȅ?�n��3ۋrR���Uw���w��3!��Cc��i��FZ"8�-hs4��i�Qt���P{|�;�s�>"j�s��{�p��{�7հ���7NT%:<��4uCh7�܍{�� �I��^I�������UK�##�I����<q�b�H��ĵ�9솳�H�i3��{h�L|�;�vɋ~�I�^�hư��%A�}�h`y���ƋA{Q��tJ��0e\�l�ۼs"q˽����j�RGW���X��?6%�FE�Џc��dZ��+I�jZ��2E�~8��<a��;�� �R%�K�~�����5�iXb�����,c�*���Yi��P8^�Y@�D$�="� �Ms�GW�Mc�3�VS�������;A[��>Mh��������$�����M�-����^垞�ˁ���\�0ϓ)��I�w5�C�����g����2��x�ٜ�"�ם�\\}N���G�q�M3T�h���r�+���1Q��R6���i�t�K�B$J�ڈ�܏�_��TD����f�m
��w�X�Ǟ����W5h��[P(p/�PS�{x���7�(�Ɠ�ԏO�Y��tj	D��$�W6��|�_�(F�M��qr1???�ZfF*����k��ER4�#X�~�JzS���~��h�~�����)�$�'�I��<����i!,��˵��"��@��?-x�~=���u�,��܇��<	J�Z�]֘<keWo�����ʪl���!v�EqB��t�$��R�7
W�g|��S<�9�����J��i@4��8^k?����=E/����E���>̄Dq	�F�)ЎʬX�.�}�/�Ց_�E>�~l��9]���nB_E�)>ݞ�)_���jF�~���4R�#�qi��*s��W�� U��ZC����插�ڄ�7��Bm|�P d��h3jμ�RҪ*��s���Q`��p9��Ĝ����e�����úr+h��{�Ay�#�	�Z$�wږ#�������(�H~���5�cQ���)7��� �`�-|����b 5�U9��,Z���%R�֨����V� ˽3�&\=����j���@F�ˏ8���f����ٽ�Q�S���&dE���h�!�I�xi�󏛸��V?	m�okDJ������:��cY�8�~��E���B����$	w�XAb1�@��o�oN�V+i�!2�K��f��c���/��{l����_!B���d\:�Iyug�RWt���Q!��`�gS�]'>	���}�Y �����^�u�	j<�'(Y�;y'�AN�ʢ��
4v,�m*_��SG�҃��R���zmy�Q�õ3�,�4޿�h�y�`��^�L�M�<�����[5��i3=���ZA�|��������:߁Lj#�F|�PM����ޝ�r=L$��Ғ�3����DOHHKǍWuz�ϮB4�aNT���T���ξ5
��U��x�{����҅֎�#	FM-t�~V�&������ǡW����^�b?hq�/v�Slw��ϠD�3'so���*�N�-?��������v���P����Y"X�#�o�ql�D'�<�'����E�� jXH
��W�l����N.1�E�o��y���%qS~9D�z��/�M�Ѝ���_࠴� �v���=�#66�-V/��;U~&��'$[v�Hk���T��ֽ⥭����(h�c"�_�~s�fW�#`JU.� � {� ��Fkթq�@��ƅzMyU?�h%rh�_=i|�#/���p�mu`�o�\�Ax�?6�����״�� ��L�w�ވ�"s��/t�T'!	��=M3.�F��Ƃ�=�U]2��l�뿜 �U	�2�E��`���h���p�-�a&}�u���c���IY�?���}�>��_A��<v!��I>�ؼ��$
�9Q���t�F��g˫�2��������!�E7@oPoc�qF���Z�ͦ�4|��$���n}I�}yU�6$�e6�gWH�!�5�.l��D���_p�o2�0�ԛq��_��`hqw��2X�G���"��
gV<;u�+��|�w1��s�,N���(+9e*�Jߝ�ƿ�^^>��`x���)�<��i\�>��~	����E�{�w�$��L���( ;r!��_Gަ���(�G.��h���~��������Y����) ���hK��C��Y2��[�`��iC�2:6���;QF�^��9��^?o�h���w@�ʲ����/�3R T��X�y���l� *M�MM�ɋf��/r��0�-U�`��g-7'�b�ڣ2\_�.ʺt���u�h��C�yJ�/~c�&��Se[���3�U���@[��xq���p!w֧9x���aOht%��L��z�I7��������/�;�>1��o Ǻ�B�ٗԫ�G�p���G�P/R�l��
ܘ����?�S���TU�����u�o��:������g�����`{;_�x�Ga���i۸tv���Z�2&���e%��c��<����XG���7��<�<��g����D>�&��"YHe�?X�^Ä�fM�ެ�i��vp���Lq��,x]�%�|gnQ���{�<q���ñ:�A����xDh����w G�9�����E<g���Ī�j�}�'��38Y�(��u	�jSy��'�iX�1S�j���7������#lu3C���Q؟��L�ͩY���U!]$��=�>��h^�97�5G�,����w�/���t��i���{���!��3�.��Լ0���d۞�+�l�H��:�J �R��'閯��4z0�j�毿L����Nǯt��|a��%��s�U�g��a=??^t�B��Em�2R�Y�"�X}<FM]S*U����}�_[T[��P�rp�?ā���ԋEs ��c�8�^bs����
�TY��y����Ӱ�1X�X�+ZO�gf��t�X�}��
U�a��-H�
����Ze9������*&��_�}�5.��� K��X���R�z_w�E{)���U)!'Ԑjc�"������gM%~�ܛ>����!j���.�;-�/4���yl` 0�s5�g#!��l<�������s���u��;��ȩ6S��&�Ϣ��-t.���¥-��f}��혂�>
	��h��׵4�+�B�!L�ă8��c�[�x�N@6����4Mv� nw�r1�yD����I^r���tZ������@Z��2���8yG~p��DgH$&�D��;�R
��l�ѝ�/%8;O�~W��&P�<�d�jcy��͞�~�hA��-М@�P����hʩ?���6�xT����7���
�s�e`:X$�+ד-9��V���8ƙ�����ƤD]��p���iX%��7Ҷ���ܯ� ���	�$�DҞU#`�Uw�/&���R����Vr+�D�/h��!'�Gh��|�UZ!ur���%5��>���n�1H�"V�`j�{�8�-y']$�G���Q�,���jNw����Cro�8����I�t?7��׏ꕣ�%>�l�6G�
;,f)9u˙�R@���&.T����#�M��0�/41��-cyx�.)�i���^!{�wAu��7�1<�w�Hn�w3��Y�\X�[�a� �
"Ó_�2"�J �M�4, HV��K�Ze=��i�c�"=pӬ�N�g�Q����d��WuO1+�Y�3���V��}���O�'Gܗ�=`Nf-�cCC��G�[Уh�z�l���J6"d W�ڧr����|�k����V 2���I��dp@�������ʋ�(bWl�?5������1��|4X��>)#1�r��n,Ľw*#�خj�K��)E{�R�LO{�x�����d5���`SS���oN��rw�8���&Gh��o]l�A\;<���?�|i��\��]�l�E�Ȳ�wW��Ȅq�{�7_�嗻�������Zi[?�6!ӽ������utL �kډ�H=L�$��z����^�R3ڟ*fs�kn����0��U[�M�u�]�;<6Nq_K���}��%5��f�~�x��2/[zI�oP�(�q�֙n��4������".�)#wXL�|����Us�����,�;�S �o4Q��gƕw������4���J��JmE���Y�q$��RUF��`4z���i�@��y����>����jPS���D����!���N�:NkӲ��I���(�.�ɾ�M��`�W�k��&,�z��F"�:2^���t3C"�gNϟ=!�=<�yH��[����3�׊�u���Ť9"N��{G��׮��~QQ���vT�1xG�--�+�z��a�jLN��Q��z�oC��h�����,eQU��Ґ����'$\��~�kw�q��k���ɡ�PIH�'���'66`�6R|�����X���%�wo,���/�x�Ori�<�P0Cl%�������nkB#�vҦx��E���Μ>~�d:��g�F�r`IX&��#�K��ק.;_W��hU/Q�xѴ��`v������u:"�:KQfT�(�((�v�"��^����Lt�7�7x�x;�cR���9��<��7C�uqe��n����m��E����hu��WCT�XSJ(�5j�b¹�XNrd8[>>5�?���I.����1����?�'�?C�|�5&y��f���W�\�fJV/�~�p��b踩���B;�t��6�����W��������娀�����s��9��F���{�^]�H����J^�ڹ�ǳSj��P	"P����}���f9��֯�|!'�(O�=!	�=L��X� *S���ޔߣ����8B�?�~ɺ�������a�ת��vt����˧I���,���?x;�>�9@Ƒgx�%��*)���53���c�u;�GA�e+��U̦P�7�z΢�|S���N�����4Ŵ;(�|`���ԒK@ ��&�$Ú4��!Vm�������w���dK��|����QyL��Z������(	�I\MYϝ����ͱ�D��ϴ��\]-	!�P�)��vCO�#���c$��59��^�չ�z}C�F���~�����+�W��^a�3x�Pz  �JMu���I@ק� �^ X�q�W��d��0�������ځ�����[uv˱��9Q)^�>����L�bK';�������w=@�����%�Q����&֓G#�گFJp�Ƨ������@���ə(MΓF}�n���X���&1�Y��XW]�hWZO2�,�X	�Г������<���hn����7�O3�[?$��|m/n�](K6Q�PaGW�N��g0u7�}P������Z߆��}��E�Jx�u?cd" �U�U��%�ci�<E������4m<&�-��n� w��Q>$��Juc���u���?;�5�kM�@�rMO��$�h�N��/������� <UO��-?�*����ʬ�h*����֋a ]�n�������2�v=���?<J�I�)��R:e2�D�y��+]�	��&�6�X{|��A�
E)&3�������u���%���XY8�J�VIC���r_��mq�� �ϠXePW~֔4Z�b�hjxT�e��T�s�@�����޹�)^�H�Ո^�T	�m[$o�����kTm�tc�q!��%�79U�9��	!:WX1ߧ$}���z�^��'��o�C�6�Z��M�?��j������!2�##�T�9���4��XG�rr�MRD�Oq{\�������� ������N�v����!y��T���&�Vz2'���{c\��ʏ!�T]Ia=q6��ÐЭ����HN��^0��3?�������#�- ������GGN���P�ċ!ǒ�_����_�� r=�7���EK/��}��rQ
y�Ƭ,���_cK;��
��w�)��>��0�(��%�����������?��}�#G�(�ޥ'Mދֿ�,)9å���W��\�3���2�xgbd���;E���A�>�����o��4hM�s���f�k+��Sa�7����l9߇-#���_3h�<m�a]�]�p��?��Loҙ2o��;�Gu �u�������7P*ï��8o����h'�v<���c��VI���+�](�Pʂ��.���t��wx�F�	-R%h�&x$�_��D#by�
�Ɍ}��h��b���Մ���<�F�K��v؈�~����ua'�/6����H��4�_^N��t�Aߢ��6l���1��k���I�F���J/?�o�I�1��g}�nVs����zMh�p{����ƞ��vg�V�������Ĺ�~G�5�hs�J�t�KZO��-oʕ���X�_G��Jv�I;�&4���9*C
�'	�鶢�olZ�є��D�Po9�}���6�r�y�NxE�M��������W��G+vg�c%� P��P%?������I�yGY]]R֩�4Q�W�� Ǿ :^F�4l<|�Ȍ-�6q��y|g�f�a�'�ֲ���)P�e�v2�N-*�!5'A�(��yrgǱ�[;�{q�k���,�Rʛ��i,���b��!�yd#^��q*3�����N�5�ͨ	�������R��e����R8ѧ�FR�8��F��Y��N�FW݂���2ʡ��� ��&���"W� �R�$�۪8�8e��E+����
�$;�{&�)k�o���jkGs�v��d���y���� bb������Tz6���g�cT��gP�
���H��$�G͙�T��C����]�T	$;)���޼�������fx��QD�j�u�1_�ܧ�3}��F�����������YD�p-S^Q�E
��0;��I�0vB7_���� �=�'��W=̈���p�����"��#j��E�{�}ף[6=k����U�얱Eg�4K��wZ�R�{��GI�^<��	�y��x=�����c��VUI�Z�=�Hy�U���>`��7�-�Z9��t@m�>鲨��ƫ�WjR�9 ���;�KES�L߆����o~nXmُ8ޜL,�;�[A� t��4�{'3�YWe���_I[�fڙ�F�No	(k������8��_q��o;�˾��.�'&�SN/	���]�3﹙J��56�Uv�-ld��5�J�F�+���AN��{�����,F��
(!Zm���r��-�<�x;�[�᫳Fb����FЦ�����zN�ͧ���I��V�	d 87@~.8�
�Eo��÷c�����ی�`����t��$0�&nN�`�����Q5T��Yڨ��셜hd�٣N
���'��n��Nu�*J�s^���D�"l�kPt�6������^��02�X�y�W��(��H�ZML��e�9��������/���hv?
�(w��g˸��]ɣNx�<�G,\�/Y�/j�͖Ve���ۣ�P�,�#j�,��p ?�+�$xMy�0�!Ŋ'��Q?���J<�H��;Z�� j������/z����*�B��JJ�������3�m� n�熳\��@F܊���E����;��s�s����f���PS�n�k�%������j��%��r���|��S�W�6�%�������3\�iy���H�|]R���Z0%a��%h�~R@Z=O��x�'�y�Ϛ�ƽ���(|����[�<o�X,��)P���&H�\bL���J���H��a�萁�[~�U�.@����٘�~� 	��[ �D�����G&I����+���w}�cq$n�i{z^=��Y�"�z�^��yi�'1��
�߳�6h��'�3������������
��F���hrی��5��ԗ�߸YQB����ϓ-��6]��$��?6��툀���7@���^�����v	�I A ]��j� �m����Fl�Ou�l_c6����X�uᅏC�!���$@����������z �u�����^�{IM���T=5h�K�c�������9�\��b?�`�[|{�>�;��mz�5���/,��d�[�{�z�<�_��b�?��z��`s��q�4눺v�
��o�)d����}B�6�����4:���j�艩yS�=/�O쒚�"��G&�R�VP,�X�ī���^��/Vb� ���Y�auuu�c�k�z���ZI�F\0���u5�󏅑���e�f,U�i>+��/����'�蕧���ܬ�1�7j�i�ܓj���8�c����d��в¦I#�LĎ��:dd�L�^A��?O�Tt E���Ѣ67�ZZ`�~,����n�t�����E��ӟd0s�������b���t�`H �iq&|zQ[�9���7��(��d.��.��v���==��T��ӑ����HUe
Jhc��XN}�u?����Z���g ���v{d��O����8K;��%��C������u��
GU�����X�A�/Oy���د��̯ou"�;�R�ݩ��F�}�杶��f�l����޿��9�����rR?ic-D������߿;b��D���7a��Fdb<���^��Ө��o�@ ����cpC�|�dP����?"�h�'�5�V�����#TT"��lF[�l5�")|b�����q9�ͅD"���)����IncSY�kp�
o�+��G��]߀�`���GHJ u����H��'w��m���:��J��{����4�q�����'܉b��y�Gƍ���Y0*�
�-#.�� �l��(��Ps��� ����@���k5��R���[��ٲ�@!�o��%tA�jٵ_��9��@��ِ���7�FC������xY�D��/=7���[Kr��R߆�=���+L��{�a�ૌ&I��Bn�e*YU`͌3�e�y�ڝ[���2o��%���,�.�ѧd��Ju2��@���z�⬍�ܳ{����FFF�����ݶg�o_~�c4\N��E/-�u��D�V��ݖ�CÀ�]�#N���ԏG4
u1��+��'+��*�r�1G�a$��f���$�����^������|cת!��W0�X��5�v)�������(2Z�!�������7GӒ��:�j<�m��v���o��cJ[��"�+/���);�� ~���-��Λ�S'R�5'������a���,�ܾ
�|�~�n�G�v��q::�+���݈$R����%+���|��a!5D�Ʊ.E���b�h�0�^^?p{�(�w�zk�ǎ�Ia�'#��9����8�#Gt�=",BW��4f����nOOO����b��#��q��Hy#G������ ǂ�;��R���)�~�/M2�ģH�y�hJI\'��ı�
����s���0������a��F)�ƽ�r���뺔���qOHM���܁.4��gjwW�hi�r|Ӆ�c
�����x;2��
����T�5*�}E���r�|���گ8i+��Xf۬����~I��E6z�a��i�9x�¤PF�*�zh:T)����/
\�Qq�%Ḋ|di(8Ypq�ݍ"��-��\O᝱E�4��7ں��5Ia�{����$'&h��K�MY�#��&ץ���]����Q;8���wP�zz�;éU��ǷA�BBbq�\���86���Y�̀���}��[��s���#��B@��i�\�VS���]���P=	W���ӎO���b�D�&�S�wD�J��ȬL���R84w.2kZa:���1��CH%��(��/�K��<�+_�7��-K'��5���K�`�r)w�`6�EK��e�;Q��́n��N�#��MO�'8�J�������g�����G��)*s
��خuz�&�v^�y��t���PıCѦ^./7Fo��N�>������.X7�(�VP�t��C;�z��ه7�8���T�YmЇ
�^�]N��B_/EFM2��8�w�%�Hn�l�RI�z�/}����{ƾ[�,����[e�� &'g]�p~#8���-������A����SCDo
�?'��i9���������h��l��K>�~Xb����n=�ݙ�`e��
1n�YCP�qbM^Q�e��^@��������Ԃ���Py?���F� �a���d}��߸iKC��F�A]ُ1� ��G}5^ӏZ�y1fPݹ��w�7�Iz'���P��ͱ�"J:�qq���/�<*w���=b� 7`K�4�_@t��{c{��h.���WQ����� ������Xp�E�h:(��gea&�w����a{�<�7Y�����
�p��O5Ep]�f�Z���qc���(�d��|�sKLJ�^{������T��۽;���,���+J��[N���U&j9�Y#�a�K��W����8�cG�ZWC��L�L�����D�;�
��������%�r
��})�.y�n�T\kY�$��蕮�>��eD��`����΀T�A���ȈN�ѐ�,�����]��kK�`0έ�wc�=�H���;У�7�di�����
)M^��:��y�@���wK��� !;Y-���3���M�R�_mE���9��cw1hE�l�c��&(p!;(}�7���̾���NwB�T�6���3�}�9���l�{1�	��p����U���o�-��*2L��F8�zE����}��Q�����3��A��H��ɐ�7/3#�7�<�7���7�Wn[�c�墧~�Fb��c��蜐A�J��A���=;�O ���׌�/�����jm���Ƙ�yR$k��pdD�G����0��&�ZL2h�~n���,Ȳ�������ȇ��\D�F6KK�H����Z�߃~y|F!?T��߷D-x�f���)馀hdo�j��$����L�;!I��r�v�y`�3���~^����G}���%�~��g���-�m�S;w-�/$yϷ�3~}$����Hw�
u2jږݠ;9�(�A��<U���>Z/ol��/����n�ofi1��ᎄ�S�d�2*�7$t�ň�.�uu��|�3-K*~��@����'�:������3�_ٽ(�D�W�E���0E7Ň���K�mm��Ji���79U�3��|�1O��9�QЫμi�J��R�2N4�[���8y�;���1<����Zvv>���B�C�8�/
��Iv��U�1�J�?���NGww�7�����A$%�Z�c�����I�I�&D��}k�a�����oY�7�K��2ە2���F<*�.����d�&��k'xWǒ/��'�~-�+�D
���b��=.v�O^L�׀OY�}�d\&��+ϟ��n9�]j^��$��I?SD��@��[�1�b�h��{�3�Sz �������-�� �H�A�%雡�6/?���VG�P�����X�%u��P���Ts==�]�J�%��l��`��+��z��lc���K g�� q��=����5Ʊ8Ət��ރF!�(ȻGk�W���I��W\�R�Z�C���I�ő�8��~Z<'$�ۧ�HlA��}O���=���NP�����T}�m��;���]��Q���3�G�q�5	s��u����b@:(��w���}�W~�LQΦ �_U�O�e�~��R>���oUZ���G�;���mXF^�����	v�;9��d�Rd1�،���s0����>�l�{�9����61�+X��OPiP�M.0�<��煱f�`�6�メ{#�/���#%����ea�Y7rG���ژ��w7�*?��=~��}���{�C���MOW���q�;ƒ�S{�E�k�\�Z��{�����D�/������"?���؈�L�N��R��n���̱���������lC�`O��� c�
3>���a��YB��~*wfR��>��0���g
Ȑ��0���uT����Q�����7[�.k�E�?���Rv�)T�أ�Ц=�x��-�khk�p��.���(
��	ץ�z���e�����Nx �s�j3�bO[�	���ʺ{@u����`�{�`Y�Ɓ����T;��Ų��t��7@���	�}ԂA��R$��$!�Ձ=>���ي�B܎��R�����G.'�`��;�����T����_���{�~����p�?�i� L��ّ��.��{_�ZZ����`EDt(���<<��{�t� ����Y�#WwoǮ�,l:���n��e�2�}�{�1O�������U�� �1�չ�pO��v"��H���Y\B��1i*��o��W)E�=9>O���vS�2�bҀ�<�f���ٖ��&�J<J�At�\z����C`u����_�Tŗ��)V��ꏙ�q���Y��U;J�[����yY�������:ݣx���V,D��D���`-�ٷ
E���.$G��ӊG�_�@���d�gm^zşΔe���~X%(�m�q��:9�(:��1,a	%�5��Ef` 9��;�ή4�U�΀	}ko�{��&38�����nD���GpA"N�D�w��a��eG0@��.7���]*�dZ��L�G@��#������%C�}�?�j'��Ԕ��4(4+���/�����B�O}uj6����V�c�`䄜�1-�"zi��Ar�j�����&�?9�2�����g
>|Lc!�M��_f02����f�{����D�r���Z��2G�P�p��o|_Q���
 %���8���@%zy�
�Dh_��O7v_4l�ei@O�>s�A�>��l{2?2�vqb���D(In�"��`9b�Y�y��2F�̌�F�����w��?2�*�.j�C��t�""(�(�1����tw"��-�9t(H	��]�����������g�Y�f�=g�g?����;��=M��пY�3�8���p)���>�K�X��/`���4�N�B��hJ7L���kkR�t@O`���� ļCy�L�n�2=�tݖ
���X�SrA
�q��@_SGh�[	�kp�n儥 �y�[�p���Z���N31s��K��p3>��7�r� D�3�Ni�g��*��[a�sԷ`	�:�K.��Ӧ7�ؙ�a9������V�2�+���N 󵻮��-�Ȓ�q&浆I�1�&FwС_�4���`<�V �)ih����0 -la"-��2�	$ue-A`#V�"��h��ş�u��l����l��Og����ωԴ�d8x�4��Ϲ�6��(�O��GJk;jFF�DQ{���7�(j������J��ׯ��][ �>��""~�	�^僬;�� �b��*�JQ����gi���`$� ��\2�"AK���UX��pҔ��E%�ӉU ����y���V����-Y��|�D�7FFϥ�����a̟���@U��N��oqt</�u�\��ɕ��q;�u�7���@<�gI)�12v�3�0h76���@���Iʉ��}�㲂�#���H;X�u��dJm%%gb��
�A"�߂Н4��&��d�G�FX���ޮ��� ,�v!��.�������?i�K&e-)(�0��>2�ު��28����v&�s�Ǯ�����N�B�1&
S4����CȒG��lDT-@D�5���?�ft�P���T#���?c���3�,�'���)�lll�f�V^Rb�:*�a<�WTOվ��p�o�$�/��)I�;�Upv���D���h�~hk����u�E���&�)d^ܶ���*q�W�l��H�x�HT�ؤr��u���Xps8y�W4k��d�F9�R.���-3�{\ �I�ф��ݭ��&���{$W?]"m
c�����uI��^��b1Vod��^sh]۞�=�5A� D�7"v�:�[��9< 謪�t>�Fw�⍰����֯@�,)�<���%k�K$�&O�i�E�������$����p��ی�z��Ryh��_�O)b����gA�?�mu�ڬ��Y�;�����l�y#�?��Ӳ�qi#0��tjv�c�1H;)R\�y�(z�Q�0��~�F��V������F�Д.m��h��T7����
�܀G.�4�)k����ԑoZ�D$T�1��u:�
�K��=�q�������d�An�1�8[��H/�Ջy��M�q�wn�*ȹ= M)��`�Z#���΃��
��+U��l��'C.t�c���v�!}<:��S��PE�'Y3{���00����zU�Q>���S9>��,��u񒈁�#�	z�&��#��K$yx} �Cu��T �E�}��,�����f!��1	p��F��i�q(|��Y���C���c���L����!`W8�0]��ݻ"a���<���ӞA^(ݨR0Fz�~UM�9.�~u�ԿD��U$��u���L_/�I�-��	Eq/o������A�vʵ��̜!���WA^��t
��Hb�Sf��S��`�w�@�=Ka\r~�M(����3:�&7w���Z���A����0�b�A�a4��G��`#sA���=�˗y<�oR$ڜ�_�Z
˔��@a	C	T�"3?��E۬���������^��9=�O
=kE�(�I�@,��8��k����BWv�*ʐX�>����'dC���ԁ�,	����!Y1h.eY�����TN��t^(oZ���W�o�7D|���\K'Q\�ٯN�<5c@��קp�\��)�%�sZ 3�2�2���EOc���b�7O9�+�Eq-�[��(P�N���h�ڀ�-cu��{��# <Ȧt�c���V5�a��v��+u<��A������L�H��Ì���}��,bGVV�¡ѓ*��H�ƶ �'U��P��m5p����
��&ᆇ��fO��o(�҇���>��|���L�n�=���j��L�c�g�"���M��+'���Rვ�Է�2F��y�l��24�G;��o���W�q	f^o��h"cw�'��OQ.W��L�?5�͞���n����p�݉Ѡ�X .YyX�)X�0G)$��h���А�g���uHZ;��c&0V���eGv��n�qx�@;����gz�f��"&y@���}��˼J3�5DA;���D���Xb�_YYֳ��㈏���4wT�!�6��?;\����6TЫ�b�Dw��[p�W.��Q��:%Ќ�wz����:(�y,�gi�	�.�g�e?�Q����.Tڞ�)j��_��:\�E��c]%ip�8#��[4��6��jǧ<�k����#��nG���!���%�s����T�AV�K��%�[��K����i�;$��N��QP�i@4�!�����%b^9����>���/��Y���kO$�aC-��
�us��yP��S�������`Ї�1��37�41���(CӔND��hC��GɳF)�/4Xէ�
�}(:�G��`���Ȇ��`�$ {�DG��"��Rn��<!�^�Cv�=yɜgN�Td�!�2��4n��?�2��ݸ�}I�M�٠�1��(v�����q 2��E-朇2�#��v��Dɀ�g,�әW����X\z����퀿�`��2�mĂ�I@�3�1_��$��g��)(�R�:�+���G� �3��W������Zthp������h�U$`S����(��u|H��OI���i����0��іC�Z��٨|%�UP:*c��D��pM�̤ٓ^x�ݙ�z���^���<ԃ�t�Df3G��y���`�ܩ���'ã�rY��D%��$с�6}��I��&yt(����Ҙ��$��)L��O_ IC��Nw���E�W�P�x��(v�!��7�ϡB�`��[lIid���R���$��U��a��]%�;�V�`]�"y(���G��5/{gT��h��fP%H~}Á?��1��~�
�:�AW�����3W�V��±�;�8�u�Ջc�
�4���]�i��l��|���`�����7<YE=�W�m��3Y'�Ӳ}{��ޛF��`O��6�ĩ��9?�����|��{���go����g�Mۘ�=�S.��Y�"� ��L'.�	to~o��Q���.9� h��ճq2?\:�6�-��̀�nV�ҩ5-M&aE4��ecY\��Js��̫�d*��h]o  6�y3��S�d���} �����:��W\;SeVo"k?��%��FGYId��$�k�7�\_��C�k��&��OH�6����l�����Y�S��ڿD�A�{�ŢP	y�
�k��m�m�o� ��\U�M������]��j�[��tāB'mƛG�s������ �Z�m��f@��,A%��F���Tl���-������� �U��}
�O~+����-��_�C��n�c���t�?�H2��Ьy�R�����#i��������UN@ה"hC�o�sP;-�zUx����lOC�C���t*b?M�CZ�hI^�0˛Eyq��� JSƲ<��kl�l��3���iH�����xQ�|��x����OꦝV.�~��D��^6��=���f5?�H��(/X�Xɴ��׀�
��6��{{����:�A.�;���T�Rvg����׻/0U�,E5�j��z�#>R����e�1?{��[����@�a���"t7
�kXj+6	�e��1�J�T堨�xy'U*�~gj5C+ۦ��r�_��7�4E������*��m��*Du��Rڊ�߷�*
������9�;�>}A��)�t��]�}�����b^<�edE�]�����6��.^~�.�j���閪�l�����BK�Gf�)Q��WO_���!?�җ��W��8��}v!��\��]O�aG�@$�����/d��P�f���.wv������V���EM1JP�!G���l|n���lu�]����4W`���ЫT�(��|��C���D���Z�i0�xl�����#�@c��u�%\������h��m�ђ�����cù�4~�B\ӣ"��K����An.Zr�е}g�mE��x嶓Ik�Qy6�K�/n�<S>�O��6���jn-�k�'�3nZ�D�b{G���},�Fwb���T6Mp���ZtH����*�����VZ]�.1j"��S��Ҧ0�{2��*^͘:���SnDXH=�뺚���o�J��WO�q��lM�5�T���3+z����!�a�ɹ#�3����i���B�� a}��{���ʲ<��fĮ3$ek;+�3�GX\i�,�y���$��2r͵�l�Ml��eޔ�c-�,��"'���'>�'���`��r��X�]\u�n<�ʅv���d����.�OU�._�L��aЌ�P���\����I��0~�oD����*ͨ)	�'$��\bVɔ�&�?<���YU��p�~LAn�o��,�r=��g�����~��#w����Y8�3I��e�oL��Z��6bC�ױ�	m��|-�+?-q��,�ynJ��]��)7Vڜ�N㎃���ǰ���i9X?�ǫӍr7^���\���.907���}�V�R��1���7t��/֙��N5z5�߬�9�s�����6jO������g��qE��z��m9dS���|��<J��g��;4;0?�;�5��Rj��k����/��z�.��u;���l���O6u3��Y9�*{�T��"���H�������O=�:k����d�)�FE)^��g�����E_���f�
Cڇ��ӄ7*��V�@�^���t[�5H'2;~�#O.�\(�d�n&�.,ze����/���lUm��;��5=�p������7\�/9��u����\���x�%��,�
z)H.�ܺr*1�ko����E��=Hq{���D�/���z$l#��~��%v�����ɻ��R��U7抃��UR0)Iй�}>n����㷛jLW�����S�0@��N!]&�b����ܺ
�����e���,��p$]��6�k����b����<�s��{���&�8x�=�8z{�����h)�`Tx���M���j�=�*I/�9|Y�Y����M���-hI�%7w�]�{������F��ٯ~�!����'M�D;��A��,����4�듬4����-|ų��0v!��qC�ӊz�\slC��Ɍ���k����D��:�_���vi���*�9�n���t�ʏ8ek�i��U��W�7��w;"6g�~��ByMxY�������
?!z���1�rխ��O�0&��������;<|�ߵ��,t�i����&��x��T?�(~��O�?���y6�h]�U�����5Yh5.���u�aW,���|/����~���M�h>��g�7q<4�����6읢f���2[������΁��M�T�T4+��BZ�؇e��jE��~yB�Brkn޺]�yg����;A��ˀD!���l�ԶB��2J��*R�#{�OL���߫���:#�c�]��<k5�Vu;Y�o�dfoJԟ�v�+�LIm�N��6�T�mtܤJ��	����(��$�T��pNJd���I�S'�Ӟ���	ɛ��y�}:�	P�Z��}kL�-�6����/TeK�zf,B�B]n�'g�$i��i(�iC3]�����"��}}��ࠛ{�ݣ�`e�n'9s�Ҳ�5�O�.ѧX,k6�I|�\����P[(yָ��KE��C��;�w+��"��k�w�w��,M+)9�v��>�/�Q�@ls��ψ���7��H���-ZCrc�gc2s��J
ئچ`7��K�:-��͗'��nw��O^d�����z�R���'*��'�b��9�
D�v����&,�oK�ZM\Mئ|ڴvwR0�}�P��U<�?�K�l�����Ӥ�-�m�0�};]0������|��j�RM߸�JH�^܎���/�U#D�	c�so����N���^\����!ʠOJ�+��3�+�B�jZI,�=�B��g�%���%�`e�ϓ笺@�1�����A�9�Nr����
X3xѶ]���
҉����p�i��<����*ʃ�3���Ɓo?%~��C����'��~���jɵ`�}���Db���� �3���-�|s�Wn|�=\e��Z]/X3\�9�*�xZ���t��dv�Q�!�&��"�\k�!P�����cJ�]����j� �t1r�_b�O0�yɷ%`EC$��C��#N�>�k}��G�v=�d
��j����kƀ%E��x���i"v3'����lbҎL_$�zR��tU��v6���B>�u�	�k=U�RA��Y���j�N��y
�d+,e�C�;71�@�oZY���V(���_�3��F���]W�N��s>
^�OWJ��zH�?J�i ����&�7��u�ӫl/#��i�RI�)/���������W��;�
�T�!����&�m��;R��1�^�:��3m���jM_$�J�����b7�r{��	s�����dg�➝m���wT��.QWj�<R�����:�[���s�׊22�\u6��&z�u��C��!�Z�a�ڭ�׬�V2�DL2��~�`�Dcmd���x��j�JJV��m�A��g�>qЮ���A�%�<+J��4��d1�T����;����#(A��	o�t�[�P�آ��v�=;� =f�S�c� ���eK]]]B}�e����;��<,���?��H�4�]7�t4S�*�y߄8HW��>�-_�9+�n�n �wD�|I�`���M(��P��f�,��=�����ţ g��]z��:�T��)�L(�й���#��Zm��Z�YF3�R%.�t�$����ox���<�Ļ���vaa����#�'�[g�p����<,V6u�/���c�F���9�?��`�9�R��O�3D�T�/WU�|Y���ϯ8���4�&xq�dTVn�%�s4�&ك!>��Pv-|Y�@���R%��[��?)�d�(�"h�P�����Zs��}=���9/K~�P(p�B~����^��V������fb��`y�ZqX9�E�<{�c㦥ܑQ����Y�k��J�S���vt����pҤ�h�o'��yq�ٔ�uA�?���"�eX�����B�o&� F-Q��lf^�Ą�����b^�����l?��ߛ��2#5f��ϰ���d�[�n_�q����g���o	�)��k��i����TߥS�z˃��ȴ�]H��kR��C~����R��.Lw�p�r1�n�(ϼ5�p�1�2v.�0�E���r��\X�S37=\��6��+
������Ԁs���B
O�!IØK$�W1.*����X�y<�ߪ��ɇKьK����)0��gs8���*�1LAڂ�s(X�)ʉ	������!�c. <��f��o~x���ל>�QBN{C����D:5��ۭo��3_�Z#�¦��U�X����cd==��N��d��'�u̓(Q�}r���F�΂��$G�>�۟�8]jm30�&��͋�����xO+F�h9����H��PWw� r��H�J#=(~}$�zX����ky��َ[g3u+^�f2\�l����H���D���O�>_HY/	�y%)��"q�1\j��t���+v����j���0�p�
�x��5��B�"d�nB����|� %���ma����QJ�c�9�Y�>/%�WZ�I��N�Ar,�W�{�7�
��7v�;XSG��p{P�L�FUUy��9GI|��W=�o;W��MVU]�[H +J�jY���5�3��O��O,�_�ct�+Y�@bN� ia/]��DB�̛{�=?��]�L�9�����qD4u��D��զ����_��(p-�Z\��i���H4�f��|��|e�3;����&u2��//�yD�ESK$���p�?����;�+�B.��O��O����JP=E����T�B@K|�]p��{�/�"B0��+�umM�ݘ�:��2�fo<=��4��]����z3�F�D/og��:0��I��ufhZ�-4NA|�Dή/-8Ї��YG�.�~y��}�'ZҪ�y� ��M̞ne���M�2]�Y,�9ӯ����xp���*g`G΋9�������d��8꼯]�e"WQ�U��V$i⎋U�LѓF�	�ɗ�u"�:훅�'H����0�k����y"���T��Ά���ʺE�����^�u�W�����M�ҭe��M>:S�����F5/�P^�}�a<2`�jy>�$`�A�y����'�l~LI4���?ރ5)qϚ�ƃ��}��H��ø/~I��	��s�c@+�<��N��7]���,����I3)L�@�oMҀ��o��� %Ƹ��q�����bٯ'D 2qp�>�����s��g��&�v\PKd*aQV� +E֐nB�uvYv��z����=$Ǧ��Wm��D2�XJE�$Bˏ���U5b:��T	:Ҵך��I�v��H�u�:~�OOM!Uz�ۮׇ���ekNsIrt敃��Ba-���x��O�k��[��ᶥ��F�I��s�F����I�كn��om�%b�濏���ww�Z7����i�JY)���m&����RF�`@�l����K� ɫEY�#\z�P�����}�y�.*��ݘ� R%����b���ű��Vޝ�{�&�ca8�0�>l"��Syp��⒐<ӡ~g�a�}����?�}�2����.�⥡�;]/5]�mv�˞���vOS.4���a�'�c�NU+��J��wԅ� ߸b[(}CO"��Q2H���[Ti�:�����[Gݎ�ٖ5W?~�I-g@/�̴eZ�0LHY訟i��ۼ��'��sg�ٍq,��v~E,�+��QU���̀�B�_<�pD4�˳�T^|/��oI��v#�d���&�_�C=��n�-@Çۧ��N�sX�$F��vtڽ]%��v�h����4|4'|x�u5ƨmh�/�@B �T���h�)?��`v�{�����붗��0g"ý�١�D~�N'"[��3	��yG���c$���8X��HY_���-��bi��H�O3�M1���������L�@��pw�fmsI�'��mt�V������$p��0�5�7��R�N+Lh}C7sfά�=cV0�F91α����1��y2ʸ�`˔)�<X���w��3 UH���a�j]��E���;�H/?~�.��D�e�k6u�33�)։��_"U+���_≈�o�Ϲ���r�4a�����j,��f���$,ƀ�&?�{�hms����4�o����%�l�� r���$��u������ �C��4$�`�/�V`������0���J�Xi%��] E�b���j��	C&Iްb��-u;<i���씮�w�G��g)��b�%>�?�V-8�oEe�8���TiUW�����iS{y�s�Ѳ| ��(I��1Ka�s#��ú��u�.qpD�K8VkO��(��J���;m�5��F��-�W[���ڞ� ����1��ⅰcB���;\�;���p���O�ķY���� ��&�9� osg(��+�PX7&nB���m��Rƽ���`8)�&_�ph��P�mr
ɘje�U�����z���MOg>�y�>t֝�2�-�W�dVLv�d`~'�徛	M*"^	�Ģ[;��1%M�_5䚯�rκ��%��$��}��-��ϝF��0���;��H��m9�b�4��<L7@�q ����Y/N��g��c��/�o6����p3��/�g�{�RG�����_�}�*iSÇ#� �>�8��G�\m�Ux��o���}�񘼝��B2w�%���������Mҁg�
^H��&��8�
I�ڽ�A#�Nm���V����Yn��������$�K_�����I(#W��-��X9N���$�x���#�[�m`�����\���L�D�!�)-��7�`W�lSp��E,e 
7�����DvP��\:��3�ݷ�r5�hX�mݟ9�L��&�.,r�!�~����h����Zn:�,BA�L*h�w�5kx��._'�~�����,F����R1xl����9:�b�5<��A|���)�P@}`��i%��y'\�����~�Ɗ��v�G�ӑ�8
�[�_�q��0Q\1�Τ�8pY��"A�ѷ�1�}�-;s��>�oRٗ�"���L�Ԉ��}��]�ҵ�Å�L����@ɞ��u��:���`偐.���
^���.rrU�с(����j⨛;CT�7'��`��Y�{�AQ,|�=��8�=����gz���}��?�Eg��kZ�M��++��>CJ��,�<͓��eϝڀ�Y����Cڿ t_�?�/����V27���蛠�:I�ɿ2�����ÚKtx{����}���-U�i���O��o�B�<_�^�*�^E0��&��}|��7�VH!��
�y;t�a۴$���CB��j!��^ŵ�m0�\u"�WF����%Q	��2�b���`�����ZC@�*n��̻c���~�J�&������ o�M�v���乕7�4�4��*��7X=��H�g�LOl,�Ws޼�����N�y�|ȻB�����wS��S�+$���MS��g�"�zX}#N�&��.>�7Qfѷ���߭%,,;\R5w==�4���T&p�D��g E��m��)�܃��*�;G�г��4�S�n��w� ;xf�������������R��ϭH��߃Wb�'=ɞ��3�;	���]K�����*7߼A�jr���{}Y�?�h�
Mt�8��A�Y�PC2�[z.�f�
hi�}�X����.^c7��6J�1�j�/5�^���?�
��Ws-�rg<����|S�dg���^炌?.���3d��L�� ���5R��0��J.-*HOQ��߳ �V�y*F���`׼��]Y�F�aC�#dƎ�
�-���Dd��mw:��Đ"�a\�����	HХ���à�hH�\E}����>��:��^��;d��{?0����K�tT�8���RXbX���R^~D��%}@��|�9<6/�S��|t����PuY����<�k����wݹ�u-����ʳ��������e�*�p#�+��������4��7O���Z��� %��|��U�52(e�����]�(�0�
���.~!��Sbi����+1:٬
�U"k���[����i��o�~���tg�y�In߲Og�{�_oWԝA�~��,��]_*�g�,L3j�o��+������nyr\�#z������O4%��eFl����ݎ�%שN܊5 �3�X2����B�)��rvj��v*V}|@��|�4���ʀO�a]�-�(g�����
=�+��q[��y�?w���r�7߱>�S�_�M�▸���va��S���0!�w�މE�u�������������&�{l�������M��Sd�:^i�l`y�.��΋���@UscUՅ6zL]��ip�g8��D�aTT�9��"�Hm0{�o��8P����� o�4���pHr,7���?<�����@N�KA4T)�(�)�Tvj-�=����b$\]��V��_�u���o8�exwTzF�j��ko��7IS��Ƕ��d�	����Y	��Z���'�%�5�7 WˑM����Or��R�gW+
��~�j���$.ϼ3-1���ET�S���2���4@��o�`_E.1�>dU���ע_�tjE�ѧa�64�� ͙E�R���&rRЯ_��(��s��̬"�=�]�J$�����b����������� �b2��n2׋�)+~y*@�����������5�����_��Q\#rh�Lre �G��W�2�_[[M�̱9���A�|!G��hf8(,�KJn��q���g;o�.�O/
;��~�vw�ъ���j�-}�!1����ʦD�bs�F8�{��w;%d�e��bg6�k��qR�a����D�)�ښ��u�E&�xe��δ�k���{?c���FzZ��>���b�z.��w�d�]#ųӧ��["���9��0�=��!�8�)L�{��z�ˬ����+tc��]L���t;�z��O?��C��,�%�H!�:1U�ID������Z�NW�I]���kBQ��0��� ��n�	�잇�Oh��X�a�B�jw�܇Åtț�(~@3Ø��:��Ix��ͣ�`�~�j��vX
����ǒ�H$0�>ȁą�c�*	��V���F��܂��b��]���v�i���|�/��Ϥ�)�\f��]��+m��t��򫕣#0:���
����;�=l@�_�4k`�O}�5�����%A-+�١���ƺ�����Gz��J�P�wHO�dv�-�'ꇴ���":�� 1�&�3E�L�_�E:���ڑ��G�I���7�W';��E;�gk�I�<r�U�a���6$f���kU�jk�_���l���b����F�1�ī*�"���,w���&X{N^bN�<�I����;t������ٽ�D��aP/��ޘ�n��/�_<~ I�:��b��][0ùC�Y���
��?vwkb�'��q��F�K�<<;[V��f-�.*��O�$�"A�r���[�>���5�E��K���a��g���9LR����KoƇ*���E�~gV�+��f��q
�^�'c��N�Y�Wm҄��ᷙjܚ�bh�S��-��+�԰��`����9�r�P��(&Bbj���!&?z[�S�� d�r���� Sk���Q�\��BF�N����3�p�ƯVN��{�GψT>�����y&�~���_D�3�I�`U2����G
��q78����;���Խr�2U8��!T��X��,�.�؏�9� �MX�}�k߁���0�꺕T�F?:5��z��8�|8�'cYH���(*z���Al.�щ{Z���+��g�!,�Y�G��>N���㒑�6��,f[�1�\��W'x��k����펾m�+\�A69l5D�XL�<Ƣ{���`A�I,q���{8pW��le��J�y���x��r� �ܽ쥟2��(ş�g�1����ګ��-KVX��Y=��<.I���t�o�SU#� G���I׍��y�uI��Z�17F��3�c3�$�hA�	�r���"�݋�:mMT�%�E������_Y�~H
6�K)C�<�|s���q߄VT��T�n>ђ�K"�O�O�����ǎ�
�d�ր�Q�uJ�����dqߤG�灐;;0�����΅k�2O%�h[i*�|�E�qQ�f�w����7���tǂ��?�hg�~@�<.s�x��]��Ɵ'�$j����/�ğh���;s�5����,C�.)@OS�x����N2x�q�F�o-�3@�J�B�sv�=��m��MG���fs����>_y�h�33h���>E³����t��!�%�&�~u)4�k�����,�Ā���`L�A��&�U�p��.�?`�L;��JAy�١?-'���[鿿0#��]�̎޽!�ǸL֥ {�?��D����O�0U`7G���$�/��8�Vk���K��?��;s�[�`��w��`��uQ��v/}�(u��ħ�7&)��v(���P�4[��*q������`Ⱦ@�1!��_�����;��ޝ��L�Q1��}����RQ�ST��S�\��V�J�V�����8ӡ=i����cc̀�#%�������Cd�g�l����w��O0BDu�]#����B�?؃����z��\s�
!.�r8����^���ƭ�d�I�j�*j3�k��3�W�?��L^)mLA~_�s���P�s|� ��@�G���[%� 	�z��ɇUV�q�����w��vfZ}�\����rԘ⍼V�-$�v�[2@HB4���:t�6���ƙ}���2��o�R��{�b-[�֨�%u5��������WGm��Ӽx�?@R+�#��(e�,$=f�����T�5nW�� >11�f�����_�c ��)�����V��Ԙ�eڐ�~�h�����4a�3���H��&,"S�ƾ-9����nZ8:>N8�f�2x���lOM��Y�^���tTG�*(}w�����޴�C��7y��b�K��#��Qxq?�l���$a�8�S���i��r�5Ο��0�	>��H�k�婴=-�F�tl���}焏��˻c��.	9�՞��Ͷݗ!����= iiS��?�>�BG�~k|�N(���1��T��8U^�zМAFn{��4������,���ûhę�^��ź���	�޾7�۫�(���'{��s����P�גo�7U����+7]"�#O
��ٹ[=�N�1]_�}�G�:[K�9M�]6]�������4V{<������xE��V�
�;�Ī�k���?W��BT�RN���5#$.���������/1;q����;�m-�q>�'I3�M����9�k�+ ۝ �gvѦ@����X
�&��tj�:T��v�7ʌ�7�w�L�����E��9�Т�¥���|�SLn++f�{��x��#ά����C!��jpx��}2)Q��f$�Bp���"y�iG��@�iLGؐW�,Zr��j���˖��/v�}�\��x��S>�}J�Ք���B�Z|��a���)���J�O�jw��`��A�g�����Uo���N����O| 	\��/O_������N+,��fعi�+���8wNaH��-)���ݍ.@��׿�>�hxm׍4�mXu��tG*�ˡ����yO���]����=��a����Lf�E����C�>N�h�����¢w���D�R��<�v�Q���^��~ΐQ^��q�����{�?���'��I�r;;��K�V�گS�,!x�	;	��#͞7�*��DQ�b�d�V���C�;������|-C�Ǹ�#!R�^`��"�σ_����FG��>��&����nM&�(�72�#�l�l�]E��)��_�n������f���dt8da<5����`a3)��_h.���5�c��<�k3���Q���H���0�{�	6��,��=b	��谱{��y�?P/7g6���ѧ��������e"���<p��t���͑i��!c��l�8�����">��ĸ/�����O?�A�\�%�*p����4����b�c��9��U��U{��=���G͹�gc�߾�8sV����Ŧ���QMsR�Ǭ�xw}~D<+����m��x�+F0��:/뼒tU����]e;��',�l��Tx��׋ʳ �hD��U�n�Z2��]�Vr�L-/+�`\��a:�2����g	���w������H@��M=������31�;c�2�e���/>o�w��228l��q�y
l+I�:'�Oם]7W�"7�x_=ڿo�f�7+��z<�k��R
��XF�Q���rV����67��.妚���=m����-���v�N~Q�
&��=��x����y�/��!}�&#��Ӷ;���� �7����j�*ߚ_���Ƃ�I(�yw����In�GZ��j�B|�s����&G�]7��;�k�}d'��'0�q���jS��H$�z��(/�0J���!� ��>��@��ţ�_^n8���	Lk :h���.����݄������dq�߷��~/<I;U��9�D9�ep��a�U�/UMT��s�zH��������_�!Y3R�S��� q��U�0~VַoZ�A�q��x{ժ���*����D�+���ȝ��F�Cآ��}~��<[{�pY�o?��<��a7�J>�W�m�@{�xW)�q��	7lj3�:�.娶
��U{����՞Nߟq�& Gm�Xd����!_G+v�#���Lu���/8X�#��ϱՋ�|+Jv-,x����)�Q5��6I+~�"�֐���?�/|;��U|P�c�9�X�ѵ^�\Z�.0�G��#�����w��u�4�t���G�L���Y�r�*BѮ)�ϖ����F�w�ucYΧ�G��X3=Eǫ��Zs|7��NOħ��rd�T��W	���̛GYkbȡ���G��K�T�����@z�Į�ޗ�!j���m�K����ad�n�K�[�g~����l��z ��5���t�s��~#��V;�.q6P�>[v'�x~�9�!��m�a�sk��$��ҪN�"&���^|����r�nۆWl�7@���ur��=�[&��__�bH�|����˞)�B�+���iC�yr��]���%�!'o�"��T3��+���y(Ý^��+�B<`mffZ��Z3gۃ|\�O�[��z��~]��99���+��\���j�<��1���;B3�$$�V��n?���@�p]K�r��f�������q�	f�����y��MS��wE>���n}����I��T������7�)"����a��͟?M��_W����g-{N��(��&Mi���g(�����w&GT��FbX����Ƈ����7"Xz0�v�-�{|�e�kM�~�t5X�>a�ڶ�+9"+5���x��L��/FT�`~�ɕo�6���9���կ�g���Cy�!���X�C۵G̝�7|�fjѱ):%���2���Y����)ˎ����;J#�}D���ra֏v]��!�搑~��A�Ǒ�a��%����i��k^$}Jʉ�k�p?;i#�j�N��[0���xX�%������u��P��a�;'��佑�����$iSg�d�S:�݂�D���7h�3t��x˰(��}x(	%����I���N���$D�FR%���Cb��5�������_f�X{�y�k�=���}<SQ�qe���	��y��d�,��{�CT廇 C�`�F?�-�Ŀ��@�ߘM@A5����sd
H�{�=��<��i>*���U�8��/�����.݃�����1'��	u�ů���?��RGZ��.�^@}�rD�N�f�s*ty�b+:/�7o̿͐eK 7-���q4��*~YT���8<ST�OE�Y�l{�~q�s{�,���w���{��2�z���P1�̜��K vY���Fi�qb�I�%�"V���}"2�ȫA�?n�0)]z$6������k=�*���6�A��n(�=���Լ͋{�ۯ=I.� 4�R-��q�yo�8O��{JO��@e�c�W ����yPk���z�Kҷ<��{�A���F�i��%��]��C��]̇huu�_`,zz�w�~[܋�l�ް�3lG$��@��5k���N���]���N��`�l�-a�D��厈{2����E]j\-�MC%�| f�s�x������v2@�Z�����94�a�w��,ip�?i�bru��x��Y�B��n���L\�z��m�U�����_�,�=�_)S�k�@^l��J�H �ŉ�D���"�����֟��E.���0����L�*0�����X�����r�6f�H�2�S__���������%���r��
��9q\,����*�r#�	����e�}	~+�pi��ww~.�͵�0�Z>y4�ꅰ�N4����,��b��}i֏:�k)^RRJ�E����* i���ˀ���.I5��w(�km���ѥl�8؄�g��i�����v����&W� ��֏߻�.5� 5}��@���y":�^e�5cq��tI�c�������6]�> e��j��J�z]'�
2���=0�>¡��/�=T���֘i���Z>m����
��~AV!�6#���Tzw�աU]"~�?;`CV��ɫ�z�߃���浓�>���CJ�c�;�&�.���a|mC'gq�4�$%�He�R���B�}��Ê��[�ؼ��ɻ��>���5�J��O�epS�Z����&��[S����=������=.(�;?v���nV� ��f��>�)xmM���p������3W���z5�gd�.q�A�ZМ�������%�v��M�^�}ڬ!F~��Q�s�Az�h�Z@�|Lc�CGcQ؅�`a�L������>@B�o��c�G�!oL���!�{;�C�4=BF���=���L�CS� �˷w6f�<��q(�����@���c5I�ſu�MA�J��ʪX_9�k�`����O��g¾�1	�cZ��"!�����E(#�ӍW@$�����6+>I^u��H n�]"g��M���y�&���&b�н���} �21��ώ��Q�'��?4fSS�]��l]e�_���߹K0��~3F��Zc��~L!���o����ϟ�&�a�g�ҼD�q�Hx�5v��f
���fX�Ni�{���~\����%MD�h(��~�0�nc��1�(�o���7�;�ɨC`����F�Jkk�[=�����ǻ-M/ߞ1�-���{35\(��4ɿ��.�#;�wq�l!�!>A�%���a1�NRfz^�>��%���i�m��:��ViA�'�B�`�{���v����SS����N�s�-��}��3=}C�]׆W͞[��7AS�we[Ʌ#.���1��;P��/&��M�����PG{�i��6�tT���9ة���BJ@����-ĵ�Z.bP��1�\�o��^�wݍG�6�R�MO���
	�B���s�a�?-����=p����σ~K�On�^�R]
g	\ރPޏ�h����R��A@T�Ҽ���h���}/-܉U0����@�����D�������5��PQ��ٺ�Dw$�j3�F9�X�^ x=�ult�9z���Ed�t�_(g���7_�^m��_8Z�	8U�Wf��&f<��o,�����u9vO�d8q��nj|HRC�P�^�"ꅏ������e��^���Vٺ�;,��O���V��p��Rh0�$�'^��*SQ�[P�|�� 2������������A����}p�:-}��j��g��JWO�*g�����{���7g�T��/�~\�E������x����c�/�1p4	�!V��GLR�3߯��=T�5�t����!���Ӱ�vj-�����鞃
x��ٿي<�����-:���O4O*�h��o��&�����Z'�+����(`?��%��Lt��G~y셫w<>����rq�]�V��<�:�Z~]��|Fu�a��0_GK��:�.ྕ����	�����i��7�Z����8��
B�����p��B*~�-B��W^9�{��b<ϯ����E�H��Fg(�
L����F ����+�a����q7�;�*�����߿{�e��{T���3�a�3���CŎ�99��Q#?o��8T��1V*���d����~�G�����ô�����R��k����|��zg��~�CN���iY�X��W�߈�bآ�����̀2��cS22��n�q/�@�\h�2�(��C��B*q��4�嫏�I�/o�����s6���߲������7Q�S�D@"���3������5S���b��KD�|�����CL��`��My�le�6� �V�����~,���^�3��|��I(	W�(�X2^�#�
���a�LN���i�]��������)jm$GG'UT���&��E��v9����j&���(�ԡ�ca���k�%���8[�4���	ɦu�b���uI�}��X���w8���s��"K=�ℊ_X�N�����k*�L������%�O(r��'��!;�~
����F�ơ����>Q[gV�.�54�km�W(8�H���������0"��T�b�G�@a7�k ��j�c������B��5��fO�pnv�V%�k���#Z��ϗ�/Ʋ�׊����x:=���>-+D�6�D�',�����U0��@�ũ��9�����% ��@��Ϟ���c�E����4.�Uijs;�
�S�e]���d������%Y��K,���r����̹0�X���g���~r$P}tL�6t�z����F��,�DRh)�).�a:�h���̴�KkE[��C��O�$599��)��QQ��z��}Z[�/���߇
��ψ��M�M-��8��jSˀdg�z��k�м��U��O��/�)�N��U�q��`��S||�N.�+��I�k���y��A�p�@�x�?e?�A�H�P�r0g!��v�U��wly��E�E���Ԇ!���6K�S�'p�j�XN}R-�����&�e�2����?�Ķ��2Jb'H3Zہ'�1��p30Q�]�}P^w����x1�%Ym������R�[.[�op��ZEX�_�!��k�u`^g]$M韈oK�Қzu��E�vYf�����O�S�_l��#����b�BitO�m�q����1dY�f(��W|Xe(�_	�E�!���@Ҽ3��d�L�n���\Y��b����ݻ��e�9�r���8��EMgn��LT��<��o��Z����v�n��mn�������h�n��KUѽ���Jcme�@8Х��nj���GsD�C��w����݌�p��1��jz_f�O�`��V}�;������:E�G��g䣖��{��Ű�Hъ�� @g>=<�S�A��m@s2h�9쯪�;�y5�T�J�{[�����U���n��9o�͕$����N|��͝��bx��>�x�{�u�no� 
Ш0%�c%��q�.�PϕiP5���1X_VAM����.��T\4���أmQi��O�4@jHr��l?��R�N�	dX`tM��oI3��_TT�/�/i�* Ր�\<��d?وT��Y�& ᨰz�;�7o��\Ȉsʟh˴���f�Px�$�jQ� �C�.�I��d�����8�5���/(����^�m��%k�%he-�(��
����4��b����-�b?,"4�i�<�YYE� ��ց"l�3���^��Fdi��6�����Q��x{���T�g&�E�'�{�^�й�Kj2��-;zl�kӹ(+g�D�
�HH���%IsfQ���BQ���%�I��F ���$k��k�S	&�J��w�\鼦����Mx�̴Y������F�4��Ƒ�HLM��3�4��-�	���
t�A�n>#�f1S��]7��ee�Zm��)J���獫���;��	�����[l8]�p�i�!� q4�t�'�\�07f�Tz<OҪ�F��1Va�{;��G���+�ws~G��'�:	������~ d�c�|VQ�su2A�28|"��f�ғ��x�1s�(Usɕ
8�y��b��qH~M;�_c�_hir���)����z�����b�3�^1�V�/�������H�}����WRv��~�bc��YQqs�*���<J|dF�~�GJy��i��2:�JV��F���m���\Q�
B���T��%��C4���u��e�K;�kSs��x6�ʾn�D�"�q�$/?�����-l�mc�!s(^�
����@�(���+!6�G",��r�{�ΪX�g��BM��Q����$�s�.�m�'�x#Kw�>dL�����_�ջ��@�4HG��&��� �Z��{ !M����'��1[g�޽p൫�dM�9J��z���sB���i�vY�?�PZW�'_��W7ܽ!0����I���>{��]���u,��O�*�b8ȤR���	�<<�I6�şD[��߿΃��o.?��x�)@
�e� D�l���_��X��n�c�0�';T�l�&���G�I�ˍ��{B�~��Wk�ɛ|$C�CR���VߛL��z��}VG�����"� ���N���]�
JJ>��x�<��A�Eh��a��g	��K<��w2�yG�o��T��$xt���]��퀷�_��K㳽�d�EwK<� �n&%��i^C�ɬ�
E��?��DE�����8Zor��x��>W�/�w=-_�)^�L�f4�7^6��DK�!抅;���ıh�s�^�~f��������e���[Ӛ<x����t��3p5������cHEE����:�C�$��������'�Zo���ņ.�U�n������~;�[=L]��4㣢�{kT!!�iR�5���{�g��QےG��}���F����2jR�a99���2�)d������~��ʬ}L��|�lMʤI&n���-hs'k�,X��W8V=j/|�V����mT��g�� ��
b
�I-�{�se�����ݧol|'ūEޡ�Z�AM����r�\�����֡J$ΊcH����?�,�/�n���;���1'B�l�ׄp�I/}�HNނ��v*G-�xg��D^ed�9��ȍ?��h�z�KlZ�LI�[#!�I������5�_�<CK���P�7v�%(��l�����xs�.��|�m�6������B(� �?�<�K�܉�X��Ϫ�C��1a���9�P���p�3�pVW��
Ǎ����c��F���	:9B��iT�f�,��a^���@�j�j i�u�0���Lc�0\N;��U�DY��u�X���H�*0 ��Ī�y��
I�fÕ>���;5��Y�u��`~�|��Մ�uj7M^��cT��i��}y�q�ˎ�>�k��c�%m�����mĬgr7w�uI鈟�r1�]�o�vtD�ڼ
wl��P�%E��*Y{�U?��*"�ˇ�ԉ���'.w��*�"��NϚi��t��,�{*Mu2b)�8mnۃ��h#��v���&��nX z��\�Mr���x���/�β�k7�.n����-���17�=�t��j==6�� �1�n�nꀌ'�v��M� ���M�'�Ѱ�;�\�a��bR��!��oJ�������ԏKX�}�����5j@�d�-����e_�Z/�W
�8� ��r��lJ�9�/w`m7�_����PQ�#6�"�C.�ڛ�3��&��]ͫ[t�r�X
�t\��陬h��A�7���|��z�Z<%��nxF.K,�
�?�q�J{͞��������S��Z��\_�v�I����'��{!�����YH ��՝�wD���޾u�7��>
��	���G�Z095n�8리xI*�+=�>'/fP����Q�be#Zz���o����_�@'Dӱ���E�CAk#��+��J��%K-Ty}�H�x��[���2���H��]Δ�A�.pQ%嬠���L5*� �a���'q0�7C�>��������e���H0+v �*��(\x���$�9vA?���g�]�NC4��:���{=�&��P���"��(�Ed�yN������F�ئC����[++b��nٓ���_���-���C/t'j����+-�l���;�����֟&����h(4_������Z�n����%E�����h+��+\������6���exq����&�`����-R�թ�>3(��`��&6־Wק�φ��c+*�[���Qd�*��׏�� h 4LB������]�>2v��d$S�y(��xd���/�9�"˖���8��I��!Ĩ׶L��Mpdf�3+�梻hp��)G�b���POje�C�Ғp�)�(�p��T���l8�i��r�Ɉ/.y���������kj��;R/O��~�qn����C��\�w������UU��>n>����
x�Z1&,����y7���y:Y`�2|iñ��]8�ǻc�@N�������;P)i溟��<���ل���,W!��z��+�:��$�K�B9ez��nɢ��kN�o.��@�vb��@?W��(���ϟ�-R��w( ��{����݃7!%B�@_�E���N�fg{qcqd�*^|��TYdl�� �CK�:�:7����6%P�r(�t޼K��nY��|��ZP�7�[����c,YP�(f������2����c;�����y�zL��h��"�N2�t7�U��r.A����Z#��=�Ũ�wqX숧����}Z��;8����n*���f㿶fd�5�����\3Q�&�V��}�3H����7�m��YM�	����S	��ۣ Hi:�U��㻉���՚�G��p��;�#�h��c#��&_�����
�ꪍ���)�r��G n��ϩ:A�/�M?��.��:L�8��%��K��X�_ƌ_�@��-E�2M�N�,�~��9f����9����W�m�)S#2͝�??w8`:�,�!�#��i�2�'HZ�����N52�9�T� �%V!�/d�KO��}��������;k�l��1�
�$px�V��K߰�ĉ��]V�*[[�_�U�N�7�G��S���_�d""�c��;�G�A@�?Mz��o�����PQԦ�@!
L�$�������U�_z����?nV"��M��M���
	���a��)!=����wf���ťPq�{�W3��c�0Z9AGsg�tr���03��Z���Vr��!�	�3I�&��(�VS=I)����'�<z�0&/{�g��e�#��T�i�5���;xo�cHFvܢ��PW]���[��**�qF���C9�����S6"N�F�o��};3_W_g�@0x�;S�����cF5�UM�,J� ]��&���F0�I���֞T�5Uǎ�aG@��h������G2釩J���ךq8��R�D��R�V�?��D&W_�=����-NE��x�9�"Ui�1�����*a��龊�y��w���mm��~P��i݇ԑ<L����]�-<T����Z�a�Z�.MV��.����)~�w��fZYS���a~���m}����|Png����{��r>#.$j����Db^ʮ���+b�L�C��s�-T�D_�:l�·�+��������S��ח?�_������//?�(��sq��9m:>^j��{�eY>f���{��U&�3 `q#���K�^�?L�>&~�0%��[�Q��t�p,GZ��[�x�t�a���J6PuO.b(�] �)�zbc$;�����qV��)'��'+NE�̏�.�O���.&�l������&�܊g��c�S�m�EQ�!ٽ�Ө�A����8'�mj;t_����{Sw96?[Qc�����<��H���cz*~��L�@�6�D���SBR��Bp����-���?D2G8>۞`�z������x�֐�������Y;�CE�P�Ʌ=*��~3��ZU���!th��Ӈh/��~3�⛐�E@˕�)��ܽyLԦ�!ir����k�Lyj�$���@�a���nH�N����!?�.��v���R�۾��Lt����~	xV�!wb�t� 	�)lӞ6���?(��/���]������ǘ4�Bx�����y��"��<�����UR����J�yO^��|����؋v��ϯ�r �m��1�fd�z٦�泥��Qf�
[�]�^�bd��'b��o��=��Y<�e^-���.,�e={F-��(�	��wk�8��J�gi��CC��������M@�a <����vz���.��ܼ��N?�J�ϙ��mz��$<�b�X��	�����4��'�#�7e�$��z��qa�Dr�%�śP\�s��=�C�a@x�_$����p�C'�I7�� D[���Z�) ��1����݄� ̶F����z�W�~%����J�$IUى^��b��Q�R~C��*��O�\RR�,m������<x���ykӗ�mY�����K�lb~f�������!��+�t�AȞ Hv@<���ʩs;��H1��YT4EÄz �9���Y]%#����ݟ�x�YT���l�7��Z�p�Z��n�g�H.t��1	��"��57���g	8��u�\|�����ԤRk'��\(���gsS?x<�b�8FĐC����#u���u���D���	���ނg��m�S����:��@M��t (�c�q���D����/�v��x����^Jj��r�����d�O/��v�Hy4$$��B����e㑌�Z΅Bm��c�q���{�)�x�����J�M# Ԡ��~���p�}5�������^��/��
��w�l����soKߌ5���ƚ-��M���LԂ?�jU���,�=��8�REL�}̓��_`�$E���]Y�ͼsQ�#�i����J��z�"�'�Nf7��Z���Cr��w\�6�M�o����d���-~#�
	���S�=-r�O��\�זFb�A?%F��V��cW$�y��P� �~"y��)�)i���]o �ƾ9��)R9� URd5��_���E�1h*��"����L�VM��Ȗ�?�9{y{v�� �^F�� ���8�V���-�{�����J^��gN��D���O�%��P�Hc8D0����]*�vT&�'99�p��|�[������.��u$/��'b��'ʣצ_~��������;��J�e�x��2��}	G^C2��
�:�:����S5��	�q�>�����ʺp�+Q���&ڲo��x��ŕ����C:���"�=!�2Y#k��n�3K�~N\'�U����w*$UAQ�V&͸��Q2h����u����hMCC�`���"gK�- ��Jρ�1B.;��)� �xdu�S!"r���ױh���=&²�y�۫Ig�1m�H�o?�>Z6�6���$�C��>�`߅����rkj�A�ƈ���5˼�N�7����G��ޒ��,�\�J�h���Em��l��z�]gܑ���Q������ԲgB"�爟'[�`���޷.ֽ؋M����U����l:`� �<�PUEeo�Cg��}J��XS�B)�p%�ت�+���.���c�y�
/j���W�&�
I�[se-�W��Y�-r�<���'��.��G�,).�R�Lm�Lzs"@[Ydd�҃��w�`	��2�.T�#*R��/�Jd�p�����"Sōh����W$�x[�7�K��2k�:H��1d�P���V��W�K�]nE5]Z���R)L��`�@O�:��e~vz)���-��ś�w�
����]���Ne��V����H;��Ѯ��5��z�(xA[m�Ϲ1\���:�����@P�Ǐ}�ư����ouX�5W���J/]?�����Y�-��;��J�?5��/��	�����w���|�������W�᱁�o��ފǠM��>��0訑�n�k�ߙ� �rS��6��g�
�+��N�pQm�!H�H�?��?i��C�����o�������Ƈxۑ��.��M�d|� 3d�Ԉ�1��T�GO�����*�<��@��F��8��if��yB`�`�%�3vDKq���������@)����F�A�/�/ �Y�b=��I�~��1�j��2<O�ax���/�D�ZWO�r��R˟63�8��)u4����ʗ{�;+`�:;�jP��)�[F��c�]����L��_h����i|���Me�c�g��y��e�H�Ȕ�aǜHπE/E%YvCۚOZz��X�y;5��R �$������; ���|�����z����ejє,����N�2uAEEa���N�|5e݌A�:�p�ڐV��������C�&����AA�U�#���S`�B�W<� �|�GN��[�~<.T/D�sB�	W-��I�Ѩ&���K�0�/���['VV{f�cõ ��,��b1�N>&]8t�,���!$�ϊ�{�(����vYW��H*������� R'K]I��@" ا1N'�a΍@3�[?e��E�,��ώ�EKH|^����G�{|�օ�gRa�'��GX����Љ��R�m�ȼ�|hbG�Pb�u��Rţ~��,lA�ܗ�#�$�N?��������u�5Av�x���*U�9����#{�֥A���-'Y~����3ao֩eߦ��3�g��>4Ξ3�`�9���4U����p�E����NG�0=��� /����PPa��5TӉ_��N.��!ɲ��,R!������O�dfɼ�5���t�q����#E�l𻄠\�)�a��^���1R*�jl&�+]$�ҝڋ�c!r�"dO=���S�O�I�T��x��P�����	�~
�]��VV���q�Y���;G�q5�4�4��{n��{��9��z���n��?pJ���ί���e�:��p�(9����խ��]�������tw��;�;CH ������z>Gk�f���	Ǜ' �/�.B;ls�<f�wU���v�H�����NȰ1*&�q�����k�<S �0���MIZ+�أ|q� +�O�{�)��"phD��H;e�i������ho�$�����q�`�۳V��ѫb��/h�n�EG�%nFҫ<����JլN���=���*���x}��+8��V^K�ù�k�~|�u��rESu��� �d�)]j�r�c�ݶ�m)Oܹ��MѼN�@�Xpױ8t�+<�~:g��	a.В���߹�"�}zEAc����SG��~�?P��0�x4���n�s��jCE�
�af]��0�'7���4�&��N��{�p켋�rZ�l�7[�߈�V����x[���5�M7`(��X����n�s�A�^��:���-�9��MX��6�;v��� ��q;���b��X�4O�ř�,1a��tW���*ӹ��f"Ω�� Q_��`�
�d:�+�-�d��Z��H!�E����dd�e�~ر�y*����C� �� >
I��uVj�q����[	\�[5���V~��#�:�a5�;V*IV�/��R������>r���v��s_Ϛz�9�(��=T*g�`�J�-z.١�K��ʲ�����%�l�׿AB�?�<������9ekL��9ۘ�YG1�7h�SK�w�VC�x�4�uHz�G4�A���S���n�H{|QG�&�I*>�)�b��1'aE���ZޥT@��.��i�M�H!�:
H�`��]������:��f*P�{�A�h�ef�ϐ�Gfq���f�|�k�"������T��l��8;m�Z0�z:B���U�<��oqt�%�����f��U#�B8��<�:���]�&���,�q���!A���$'6�/��T_��	i\��;��^�pW�E�����}v���i�;�s7)v����m>h0��#��IxD�`Kz���i��[c�fJ(Y���e�3*�إu ݩ�큶����T���f��]4�L=qY��CN�)W�Mh쒣W��!<w
I���=>�N��@�����8Y9�,�odġ��x���i� T����_"��� dD�M'
�b�d����'?�bK^��X�%���>���
�F�D�� &��7�ct����,��w�(Se�'T�Y4m*a���H���X�s��ɱ������GB�WN���=))�������_������hN�g�v�)��}�p��m+y��TV�@xR�˚�{�%����&��J��o����c��"����`��h���57��
�v&������H�hx Е�p���E��	��*V(�$�F��=�_��
d獫��h�ɛ9	�o�k~��S���5���l슎)_' W��枿�DZ<g>�!�mwø�=R��N��?�="]G�qEk���x�c�:ſ������9���9��+bЅ{8j`is����E��כ���:�M(apA���4N�SX��v����;��뇧 if�i#�,��܀p׳�s�Q�+�J��@��sȼ�Ũ�t~)�Ĉ"�_��L|EBs�+v��*l�"�������)5�������0������^WF۠�
{+��q��%Պ�Q��=@��[�g�#��:�_��D��n�Y����<�j,��1屾��W_��B����y���� a��8�{�ㅪ5�S��x�'$Z���������knKm}�*���ۯ���tYN����G��N�\�.t���y���H��T咐�6���W� �z�Ψ)� ���z!�Q���9��S������ ���u fTmf��1�6gc��:��B�2�t�h���T�� ����[|Q���F  ����kҔ⩹����2��DD���K 6�I:s;C�pu���=��3Τ����4Ʋ�ڼ������;)a����N���F{�b���t�?~��ӏ7~_-���J`�N)1aIa�rk�W�Σ���#�Ց�C�{j�o�/�f$G���JՏ�)�ߍ�!�S�� �H�ɂ��~��k�p@��z�,���=p���ot�ڦ��r&������&e�X��R��/4�Ps?��|)I�Ew��5�!Q�������dS}O�:���7���M����*ץ:V:�g�l��pm6n(���
Z���n6������M��>��verJJ?U#�Wy_4?~3�X�l�+� R�S���m���� ��o�A�y.� \z��w�����/��;c� e�<2���?��@v�t�>�*;����`3���h
%�=�h�!K	\��ǜNr0o�Q�N@;�mtU��7�%�<��5����Xh��bz�r��؊�ϻrͦ��\LV��u=�"�؛�>)�Fˎ�\ީ���y�ĺ觨"^{������U�a��{���scf@;IT5��B����Z�<���n�9��e����-��c�K*)B^��3_3x:PD,M�x�4�<��Y��"�5���^��͇_�E9!���w+�j�~�"��[&��B�U�́���N�SK��pJG�\2 ��;u�W�/,+Q��_�a�i���3&�;�@8���nM�[���Q���v;Ld~s�߇0f�� Y�^��ϯ8�FK�����>Q^��4B
	���ri�l>Ύ��01������Ԏ�������P)��'�ߞ%q?:�����09K��ka 	pT���fcS���90%s���l燘S�7y�V�T��&��w���	�2�F��?8��u:C��機��W�g�9�m!N}�X��)x�n�C(�/z��5|�w#�����ۙ-���>�s��x�'�l� �>+g�u*����J�Ď*��kL�.�߼H�Y|k<>џ�,_4�-O���ӊL�����ֽo���켖����0j���x�xc�@w�+kb.�L�ql)O�	�����䪲����j~�u���¿����U���J�����v1��3��)��@P���i�{<�B=s`"ƣ\�)������d�X_Ȁ�:�hI���'��nx���`�⅁�q�'������@P�m����������H8��꧒�n\������ �e��"u�]()'�)��>M`[��<���J��N��,QC�?�t�	y�.)1��U�<��2�x�꿉�f�~���2��)~M���<f��M,r�x+���|X�<�#�N6W��!�Բ����7�R5�!�%��/,bz~��ew�&��,)��hQg��| �=�t��fu������Yu�(��Va��,p�gQrSj�D��S�dO ����&�x�6KN��ŭd�R;�R�OK7��5�	��E��\��+I�i���sƧ�cvK�@eF<븻�����o4��l�<\.0�x,�h���G���'X:��>r��ίNV��(qrl	9����=(P��˚a$�ݖ==�K�U0i�ɮ�~��M��~��k�P��~B<��L�Ma�`u�j���M�xY�m�y.q�0�gw���܈T�A"��@)��h�/S����O5ڞm~=�~���Ţ�F"�����9�^W�&��R�*���αO���Ѽ,�3�Zܴa:�d�kc��)�.�J���'�)p����N=�
��Qh��0s�b%Π�hU}I�Df���Hf��T$�v|�����BU�tlUyy��h���n,�)�XB<�R�Â��%~���sl՜���0���o���47ȃ�≏�����gcy��k����xd�ㄬD*T>*�����v �0:<����-�}IK���xp��8}¨IUjލ�2AH�i���7�@ڨ��Kp��>�mj���Z����6��<�=~�Psv1���L��o@������t��(��~R~LDǴ�5|��4�Ns�����pZ�3{�hF,��Ue�n�(�S��ڜ�>��r�ۙ{Vu�!�Kt�ll���ࠊ�%+��IY�7@b��}��t��'ǹ���'���:4��Xd�(]����+�:�8x�k�Ǿ �
O��z5O�fN�^'��$�7@��lW���&Vz�6���s�ǫ�M=�j��ʞ��{`�7Uvj��&���g�YWW�=��(|���+]�g�%p�Z�&2����b���r�M��W~�X���?M͍D�C�ز4����_����w��o�U��!��|Ͷ�ס��fB�n]�5{�R��%��Ì$�U�;��O�w~�����!�N��Hl`[�yB <�`Sl>�h�a�>�m������F��S���	0���&�Q��@�MT7���$�x�����#��D#�vQ�r���h��f�X����3G���WN/&�(�*T�a3
��O&r��N��_Cè�c��:no T�M�����cڹ�f�"u�݈*�j{wi��ݘ�3О���M�q��%O_A�����)W�W�;3�?5�^��/��'��aD�2j��1������sbYl�8����	�K�3����|��6o�����`/FO�m�S��5�|���#��P����i����3_�����Y%�������9���\�9� �<�2����_��b�9��a1
�O]<��]��F���OW!����:L��A<�#��&{RԸyd���5x��AGF�q@h}[���&������E���&'	��[Y�cV�`�ϰ��N~-?��I��m}}��~$���?'A>]}�v�t��+�c�����fps߇ñˌz�{:����cm��bw��/��?� �0/���������:4`��J��xX�����߾�<�0�$:]�1A���c���8M�3�t������v^�J�b��"E�G;�E��9�v�ޟ�y��5Ϸ&��~k���>7������A�f�U�ء�d;�~��]�Q�<wA!����>$�w�8`��w�u�k:�yZ��c5���t��"Ǯ��q�'��[!���Nii����oN�%B�j���?��I����p��m�୻��(Y��W3�b�%��"f�Ӗa=L���#E�X�L?=�j��w�.g���S�Mܓ|��=�|՟��H�90\�0������l�a]n��*/lx�f"��)	���D)K>������s��o����W�;@�ʵ��?��23����\�������S����ǋ����Mu�ӁE�̒�*n^f�U�g� d<<�.8���q����j|0�mZ|�DeG*��kӽ���)�_�m�
��33Z��?�~i[\ʪ��$ {���џ���嗰,��R����@_��v��Qkt��E��x�-��5����	?�`�~��MN/���2As����qb��s��=AJ�����5#ǥ��3M%��d�o���f�y�M��_'%	�����`'.�Z_�$F ?F҇>&��
<%g\�J�h���u�45��lv��ϙ����+ҺÚH�n`Ul��ʮ�,һ�*JPi�z(J���"�&Ā����T��[(�����H�&����y��{n���s��Y��܌���E��A���05?_M����Zy�U
R)Tw����J��zX�����MI�]�:�' 1�Յm�����UK4��3Wmm��#�җA������7u����{�XzO�^=����&h��^-a7�����^�҉��RHξM��d��n��l�����F#i���c��9�fČ̰Q	[�vI�d6�n&����a(��J�#\A�쪣�#�9q���Б<���ۆ����2�i��oO��n���f ��G���}:]_�4A%v����v�3��r`��"�n�-9���ɮHK�]Y_�{\��l�}���?�䔮#6���Cc���?�9hqje�h����wb賲m�����L�獍�e�̀�*�g�[ѯB̽VY<��`DJ^��/�.x[�Q����`�2$��Pr%�T�T��<Դd�hw:z�0��^j]����36���c�5��1D�k��a��E����w�a������b;[�,漘C{�!d�<�$-����"��Ζ�"5M��1W�3��A���� ��PRJRW�R��o_�`�T0[���_s�K�^�hk?<�J�38p���̕�������A��y)rw���B�6���}�Jg:���_�^:˹��b�(�kn&�>�V{OP�g��=��4�(�-r����ݶ�S|�1����o���d�j�:7$�[�3r�u�ebC\���B��^0���3�[����.�U�C���G?F�D[�t�)}�E��J�ʱ-\�IK˃��.o$X�	 �K#y"5��r����#�Y��7@ P w���Q�:�s<i%�
�x��z��M�A�3Y�A^���14�4�""޳��gdĈ�*m�\�u婩����~��>Ix�J�S�n�S��`-�X��BT�C65	��PE�
�P-�C��k^�S0T�[�P�����
�	�=XQ���Y(����n�,i��e�B7�x��ݶ~��h��<q�^��VP��ɹ�u���;���JJ��>L��s�̌�e���u��z��+)c�bb����L�k״Ld��URyn�F�z���A���\�n�[D3c�$5U�UZ;஡��=I��Ŗ�	��m�o{1h�R�i�1���֧bb���
��*���/�qd2d��b�2��� ��ͯ�K!0��C�,�u	0�ʰ_$ �z�/ �/�';n�ۧ�����x�$��������.�9�t��iﻏ�Kf�b]yi������Î>K�`E��
��#�^�[��ʠ��m=����}M&�+顺�F�y���7���5�q_e��?b8EZa8r��MA��X}xV]X�-����ن�e<���x��6x{���ZI����C�+��3V�v�Q	x�����o���3G���,W/{���W\l_�~ �P��n���@5H�Q)i�(8G
�h��y�E���7uK7Hs�����V7������c���4��ְ������&Ed�G;��P+�	�!����"�r������&�a͘���G�@�=�S3P�%�]\v4Ys��r��V���Y��{�UAW��ٹ>�&J�3e��S�τ�㐬9]j]u���P�/�N$��= ���jt����g�Z�MQ�"[~�9�O�6��5\�k��D�K��K+�v�����Z�I�1|I�还�W�R�l���},��������,ƙ�ѐvA��e�L�U�f��\b�0�>�(Q���I�s,_V���+o����jȉ�hZ):)�T�o��ԯ���Y^yJ�L��v_�ŋT��FE��.��������uT('�/܂k�{��h̗�W/i;�F����H��6x�;��]w���mıK���R�Qb9Ci�%A�ؕ��5�ީ閉K�t��.��.	���0A� ��?��y¶�a���X��7_ }� �)����F4),埔,s.�}-��N#W-�@�d���XIN��J["�رOl�d6)�8����=5l6}$y��s^/�}����y� ��ȚDz�|Ժ^�H�S�ŏ_���s3xR{�Oa�b$�������}�h���D���@7���@wh-=L�ZX���-G�l��K���%@���ћ�`� �b�cb6�5�G���w-v��Q�H�"�B��i/��GJDkYޖHB?�8{
XǝHY�[�Q��W�'��̶یJ���o��-�X����P���.x��h��ingܕB�b-������Mn몛�\�^EP�(?�G.��l�;�~���_�LU�<�`g���֩ՠ�ȹn����;S>��h�}����9@
-�Z�)�s�e#��w^�w����@̪#��Y�͂녘��6zS5���������*��>�@[�2�I�X��,X�`[���έ�D�����t����s�I�6^G��_�}�X�k�g�W�Oi�jZ�� ���q6W֞��x�]ظ��U��˞�����a��11�s���N�K�����x�Ͷ�@��k��[��^���&�Ԗ��7�yI2�N0���Fc}���v�͋�w�%�0f� !� �Mj�S(hӌ}��8�-��C�AN��a�@g�o��ܛ���F����x��Bq|�دZ�L�a�_j�M��T��(J�K�6�"y��cV�2��1�U�"���c�y������?,���oH�R�������T���%��鏆�v�v%�d��G4"����d��Q`1��B�Bs���~}D#�i��ZյjLC��}-���V�`� ���  I	���nn�'�N�V!���wn�}���]&HlA�q�Ĳ��.� g�!���N�ae�l�7	���ޙ��"�w��HO{��`���]r%����U
B�l�kو��k�	-�<s�a�;�����_��hE]�����Ϙ1����[�\ڬAkT_`!u�7/��/)��f����s:��8��
�	fm�M=�eb�z�eXO�¨��.��y�%w�ע��z�Z% �����kn�f�&
Zܩ働�a�e&���4� �C�L�3°����T�2��xkfG�0e��5;=����:��D��L��L�,	�E8����"��Q$?c��)�w��=<��X�Qj�9��B;�	��=5�.�,[SF�gH#�~6��� t����� ���F,v�ݑ���9��@��f���/�d�[�l�WCLs��?���U�}L�"�g@HD��N�t?�䠺$��oO؎j]�#}
c�]��r��d���������R.Y�dj�@��ux����m('~�Ψ�]�<2�܅�}E�(qu� K�$�܃�{�1[G��}ȋ�&.
\�}������N�b������>��	�ӫ�5g��d�/��Ď}�����Z�y� H�F{��M��M�2쿒�������+�aUaZ��ZfD��iUaͰ�Uʑ^����"�G{9m}@�����I�X݊B�~x(� $}r�X�Ѭ@���: �P�v:�6rō�?��V��)���5�z��R��{���0pÍ���L���0T��JCx_X�@,�)��8�])JVHZAU��DV�4	Y�m	��֥���U�> �u>�lul
�����Z_Q��B����*��>��%��qy���i#�����W�Gĭ�4U��������Ό�;���AY��|��5���Bp�\�$��Io+?����l]�ab���Q���>4�oOފ#��0$���� ��Je�W_�'ς���*�[Z����:p<�|�^�?�(�7[����j{|����9YО;�4r	lR�'@rY]o�|5g��3(��;��k��B]���.ӛ:�QA��Y,g��kX�ѹ0r����@E�ꊮ�&t]�ó��g���{�nz:Ũ≂ tCxy>�Q<�]�e[�MT�gGA�,�X���\�r�+ɫ54�Kp�O2�Mi�K<�r뛘��5�{|Y��us=��p�]�+F�͛L߹ߟE�Bb������%g�m1���`8�V9:<�,d���4��$5��l?�A}y��> i��q�<�<���.ۊ[��c��eԚ�����l�q=oIA���0�U�]��R�5�����bH$"�:�ӿ�ʎ�Z-���q:��r�3�ЙP*ڠ����+���W�d�X�3%�^Α�>��&��ki��8R�?�6��qS^�ȟ@19Y�����+�,�qŤ@T�
ڤ�o�,
�W�h/
�|5a5�-ꀴI6��F�7ѥ�� ���:EFҪ]��_�r�ᵷ����(����T��b��0�ii��edK�a[)x�)j�H/���9V��g����6��w�
0��=�#ɒ�H?F;��`��BO[!��֌��+���NM���]�n{��5@q�#����A��*㌾*�pҺ 3Pv�T�	1�M�sG������{����g�!~G��W暭mU�\X�P
,�4u��p,W���θ��gH���̐�	U�˽�>��c�	����������wq�u�k���X�b-	E6���LlE�Llb4W��k8�3�i��B��7 �3A�O��O�Fq:�<�I	��He<��3L*y�6V+r
������{q�7�R�Xal�<��F5����G�pR�PMhCR��:�D�TM�#�/����K�<�j���di���k��Y.�>�˘[6�}s�b�Bu�G�~��#��T.�]�)�P�YW>74Fi= �����O�S�5!��KgΚ����d�F��*��VS�՞�";��	^<�|7�	i�X:}��H$<rUf�	�/�(���M���O�=;��v�!��yǘ�y8�tJ~�->�+5������s@ׇ���2za��2\�f��Λû2�w�>�'*�? ��g�M��Z��z�^|�6Pk�:�	KVܸ�:�7��v]��~��Z}'�.�>������Y��ȕ�S~M�gf&��0�蟳�B�������v��ݜ;\�᠊'�E2�6u��6'�:/�3�o��A�}6������m�I>
?V��Q��y�w�(pG��Ju]o��MP��x{���f��,�gJ�頁�_u).&e�t�X��/�жe]�6R�9d^��q	��r�,!��B�k?z���^f.g���n�G!S�n��ʳ���j�i�)P��Q����r�â��X�PyGz�i^.ɕ�ҡMD-�ݢ���8�XXT���-ـ=�Pȷ�k�� �����7��PK   ��!Y����`  [  /   images/fc6d97d6-a1d8-4630-b4a2-8bef38b47130.png[��PNG

   IHDR   d   -   X���   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  �IDATx��\tT��޼�QiԻ�PA	���b��[l��N�v�����ݜ�g�l��8�u�u�u��F�`0ŀ�$H �PA�޻FS���4B`p��q��#kt���������G\kN��G(�B?W�k�}�t��E?��s��n��ݕtnzw�Ӊ� _�d'@_�l6�t
4�C:����j��3�A&�D�G���1:j����^U�>00�Ŧ����胃�[AK���FY
��F1D?�*���0z�>2<*�p��󆇧F��Xen��^��2��Q�����d򄗷�|������t>>����6�S/�Ԑ��ޣ��@OϠד��9��p8�ݭ�=<��&���e�Fړ�c����tⁿ���p��uw�ႃ&���� f[��
���+Ve!vjm�7�������"19�5LQ`����ǽȞ33∩CB���/�����Db�F7�}���>���P�_�J�����8Dk1cɲLb��8}�{�DO��e6)�%��-����;s���L��;��:,�{�|����;8��$������E����L(�?��u�x���h^��"����X*N_�?<�T��t���G��Z<���$�`���7j�q��<��͢H$�.�a��2<���E�,l|CC�z� �
=k����XT8]�R�U��;����<u/MX��c;�����ˁ�����O֢�d=��@z��6�@ىP���w��l��w s�B�w��$����p��?@V&Y��'����?�BkK� 33]��:��/m|%zz��ޝ��e'K�{a݆�bm��BV����}{<p۝+�����F֌Q(d�����d1�ٹ3�Ghà1U�]���;�����CGkP0+g)V���[vczJ|�u�f -�&,_��m�� iZ7	O����,�=oݸ	S�I9T�1q���h�����jFp���B#���g�c���[��b�����&�0[6BϦ���CHN2`�r���l���>R�F1�[�ۉ�L�o��?ۈ��Q,]b�֭v��葖҅g�ڄ�(V��c�6;��TbP~��f���p��v��"g� ^x~1Ɓ���a�N;�U�����l#t`�Zv�&��̷���An��끽�2}`�";���"��7 )�y��eN��a�)x`��E
�8�z��w���,G���(U���Ě[Tlܼ�A�}�8S����Ik�Ӛ?�{�Z�u�*��������|�Z�~ˆ�V�F�À�
�u�	�u��,�@{s��ی�?r�9������wۈ'e�O#*z��-=�-��QzԞ���8\�Iww�#<��/�p����13����G�O46�PN��!����� �2<���*w�F]�9�HnjI��[��S4�F��x��o�}�F��9ȝ81/σ����J���R;��,X�'W7�AG�{#m�0�E��ޑ�`�E���;`A驯����%�mqa1������%7��Qb�i|_�--qS�JF���"e�ß�UW7Hn���q+������#(ȅ�3K�ﰢ���g�Qp�8�(Ą}����r�2��SPT��Q�e6z�AF� :Z'2��HƋ���I��S���1-AG�b�446��eV�[��ԩ:���b��4bz32�-X���)JAe�s榢�����p/����T[1sv2�dmx ����Y���H���G��^�|���E(Ng�н<��Y3�hvbl;��(@�Ҋ��hHoo)��+��|�0���&�0bq��6!HH���d��.Z�W�ɏ�v���
�5;0<b�=�^�p��z���L��D{N����[w�I�]��v�l��(�xU#�t�5-��={=p�Db|�x��d����z��,���Uথ�Pt$��\�<K�.2��(����B�;ɂH���13vG�

i"�78�m� FѠ)(�/B�4�՘�%Kc%�9\��SFH�p����'9r�bc����Ś��W&Y�q�#*�C�.�M%�>]�QQa��-!Xuk��s����b�U��X}k��x��|Z��)8]i���f�(.��*36J�(+��-krIV��XuAb�q�zM�쳕&��9B�:=�A�b��u�ƗxPM�C�Q���K(S!A�Q[[��rs�:,�9O�X���LW�ڮ�����ROMn�"{ɱs�U.̝�C�ω�D��҅g�܈Y��iI�h\|"�<��&AM�W�۱aJ��rc���M��Ĉٴ!;�iC�Cx��-��ƚ;�q�Ǭ�x#��_nAh�?�{��k�W�Y)�lv��y\b��~��w�oX nI�!N���;Bn�!�?^�g@h������"��)BOV2���ۋIH1��Y:�F����W�^^�LrA�y��P'���~y�&'Y���/DmM�y�$�Z����1`�T�_$2�I���"���'q�����G��#Y�#	�����8G�٠�^�A���n-�$�tٹ�ZhQF����B.�xB����TU6	]p6�y@FS/��-��3ol����thI��`�^NW����O����>��N����/���y�D0�j�W���
:�:��ʁ��*�F������in:���7���Wppfm|�p<�f:�s��ێ
_��e��g���*�;C��Ƈ�&�c.���pD���ϗ�3�ƫѵ���ҹ}S�;(����}���<�����O��J��``� ���$�2����� ��3�h.��?D��>��&4��T�×il9-ͽR�ȃq�	�նQ��C���s�;��c�RAA�$�
�܂��[����	C}J�|�T#��+j��왴Pܮhp���*�4�\m�XK��j1)���'�[#We���@.L�qU�M��a�P����{ ��dY������5)�8%�(R�c�tw_V��eQ������F�Ȍ��7�{0=-J\١��^��ukʗ0{e���+Ȅ�]�[���`�:�5���2s���\�|�e��6�]jY��{�����F�|Ė����u�(9�8
�a�f4����o���j��q	��zlf���Ȩ �,�X39�������' ��a�5��PO���BI��s(����ŗ\w��&(��gh��I9��Ж�+�'_wcXIa^*�b ��6tZ�P?}�l��+VgP��3)��{�`�����~��FF��8݄����t�mm*N�:��v���S�E ��E�1�U��ji�$�F�{1H��F�-�ɾx4����+lq�Ŋ>�S7ç�����J.��������4^��`�H����)��+qH}0!^��4��nL�L�Ŝ�dXH|���уw�*,}#�*����|�DV�e�p����a#sy�~蚖��1 ��ʤ�9`��lATL�d���
6!�`��5����~�=�u��������]��>o~2��%�X�a�$u
��Z���8���kb��YƵ�c����q��1����0�zbp@;�<[�,��O���'�l��w`��,-:	��?o@N^6���JyN��s�0�kAi����CMM1ҲnEP���1nD��<֤��q��G����>�V�F�#�>����ЖS	�>*y��,�m[�cf�}ؽ��,���!"�EG��������I|�ᒃ��tknU�8WQn<ALlv�v�Z�d+�J��zzE Z�� "Ҍ��~)G��<������[N�0V�� 2����`ܳ.[7���>��WV;�6]�Y�Td�Os��1z)�ݨM%���Q;`C���}*{�h�_�MOl,��P_DP���yTt A�.��iI�(o!q?J9���s��>�c�*gNbz�"e�y]lhGXd&}Q��+�$;�{�5E|�Z	�x����z���!�2ns�x����#�5���('֣c�k쫤�<�`pJO\�/�ir��.�#�?�PV\���X�c=����-�O�\���<�|I�?{j!~�ě��(��OȒ�Q����M#��v<�jF�� |���	����\��5z{���9(�⮻gS�݁��R�#n.9��D�I�?�H��CF���"`v�ArAY��������獦����w��ݷ����o����/v�0���o���}�P�N�iqJ��,apc�޷�B>��q�%.t���Y���(!쁯�l��,ET��]����U2�����Rp�8K�8Q^NҚ��ٳ%H�u	e9	)��;�Xrjv�Z���#������%�n:,Zg�~N�c��gYAYq���='�|p�7ٺ�O��~��G�ط��˹���1yj(��FY��ش�Nf�JJou�,;K��Z���
��Z��������[�
���q�sl��>�� �g��<=B��\�Mˈ�����N�%��ڱ%+�ʊ4��t-.�ݸm[�i(���u5LO�!+�PV���V¢�K(�k�\�5��o��ri�}�c�e<�gq���c��MÔ�`t�@8��%	� _�߯N2�=�	��(�(Cj���t�QY8SQ�U+U��0z�5UGYl�>�"����o��R�5�����/O^ aۻ�\�k~G� ��;��d9u�(<24*�^.8�hJM(+��/$2ʊ�U0u�(k��b��w>2�o%�gAX�i��?���H\P�͆��
�|�(?o��ߴ�k`�����n�ģg��_��x����P���U�&e����f��<PI(���F$��0�QV����z��)��ЁN�t��]`��B��F!��
-����5�cTyv��K�^�{��|���V<�ʮv �e�]c7�9��-�Ύ>x�gQ�(�P�A���PR\��,��Z�6+��yP
��p@��n����~w�݇��/rNM�0��t�&}��wSFpi�N	�«���F����iBY?�QŐrs�����P��q���E��)fn��E=��1w?	��.TW�~D
�gL^��X��̘?c(�T�E���O|���'��c�҄��#˰ck�/!�PVcC�g.vl+�g����%G�0=5J&��ű��,�}_KK���P�Oe8.x{e�eDPy��i�t��y�`�*���X�ͦs��;Vܬ�Ty)Rg,�tb�i��z$�Z��"�0˵��Zy��4|Di�:���O|��nv�ki�>r����?Kʆ�
�3���.��_�(zP�I��K9F��`m1ʊ������	eM���>Ϥ�x�!~�L��XS(P]�>��7c}l$(o��Y�c1^��5�g#�jW9�1d�]�dE��3g��Ȳu�8<�K�x��$�s��<d��K �Ok|�v�Bv�*�[$�iQr�s��`RX��h��q�`0x�l��W	�*�����K���>�@�̾Z��h��c�L]XP+&x�=���.ŷ=���_�~�!��{���EPo�v�}{�����f1bb)s�sߺ�8�Y?Gn�-:'���戀6�w���I���娮n%�D��_��r1��3Υ�z�H��׻��
�`���*Q���2������ʻ��CH�/0u��HH�+,.�����z.��2��r�����gD�gv-4�,����b��9 �3rc���p0d7x����BZt�V�>vJ~�����_��S���K�x�tdω���G��=8v�Ԓ2=B��?��[�WU�q�j��"?�}R�O�{�Ճr+>9m�(p�|#�W!�`�\�����{�6*_�fjw���)'����1k>C`�^p�
K���Ƹ���*sf� v�|I\'�E�~�ң��ʡ���B���Yj\B�N\��n^N�)c���o��p��t�'o�_�IY˙In+`�)��9(�z[�\YMI��L�3]�3�ٍ�X�!��B�g�FU��}ߙ'�ow��f�s#w�y��;�\�௷)�Wu���e7R��@��Ä���H��/{��F��|�\ǃ����QԒ�b��G�܁��kq�9<��	�o�V�[�d���q���T�����eS��*���Gq�������$7��������$��=Xʧ��*��������_��^��@�G:;�v=��,�\-u_*���DmM�\������>�����&qU|]S�����8�✉����EP�δ���v}-D� 2g����o>p�O�E�Wܾ���m!���3?�Մ)ɰ��x�t��K�k9�X馃��D��G�Lg�r��Mh_IQ'���&~��W~�������.+ٸ��w���y�E#��C    IEND�B`�PK   ��!Y����#  �     jsons/user_defined.json�[s����
����c4��%�d�ql��S��J�j�"�:''���rt�p8#+����`Qd7��o ��x��e�����ǘ�l��x2�9-�f�9��V�|�j��G��/����^���ݳ��|��bv�Z/��,ͯK�Fp��q���1>�_�W�&=�Z͋�ί�d<����HT$z���!5%^D�+
��c���rv�ڎ����Y������D�"8�Ć�4,
�����G���l~2ϋ������tvuy�~=^��<ǌW�1���o�.>����hA����%Y�g�\���I<[-g(׮|`q5+��nv�5�j*���ZY�@������y��X����r�kt�|*���4���6��JX�p-�Cu�3������^}��>fx�,0΍��Y{@���7��ج뻭e~�-�V~Ƿ��˴\�66����|��-�9fIr
�F'Ns|�2ؔbH)��y����b����(��}L�h�[{:����\��6��o�r�y:�Mh�g���˯����sZ�ߘ�OR)�<��f�d$d����w�>d�(0��%���
 ���]���ŎA�&#Y�o�AC���t�����	XY)��i��o��ɹ�q�h��%�a�q���ys�5�	0m+�C��~�ț�*x�
Sq�\L�j���:�h��hPa+����d�y�6	��A�JR�`b��,���k}�jWz�Jh���,NH;��|�n��*θ�d׉�C���S��M� ��JN^���>�"w0�	��q��c�@��q�'���w�(�׫K�d�����d�X�31J��37������u/G���~��zu(w	*%��&10A� �adB!k���%��:w���QDB=�t!�'V$F�1!�얻��|��B�FϫGxv&*Ne�0lRLC��EWO���C��~I.�!g�(���q	3	�5�(H�L)�q���1|J���7X�`}��}�����ϋ��W�W'T"�gF�ёp�����]OD&���p���w�.C��;�*���s�r�����	�F��r61�R����4�?�9�T����X�]}��V�j
�.�,���:<�7�V�s�eV��X,"�h�����G�:��r�?n(�q�9�Ū��C`��)��\,~v��X�\"sY�$P%�myI|Α(4Lncb��k���o�ͷ�����D\\�KΝ��Oo�\U�.誶�O��o�ǈ��|*�gW�2�������{)�d�N7_gJoyG�٥[����	t��$���S�F����N���<�F�<z�	'w��D�<dEЍz�YI�"1B��E,/hW�!�QI� ��8�E��X�Z�3ţ�]T���<"VY[)�U�<�;��Ͽ���~���go�UZ헾�v���ѳoNO�p�_�n�Ev/k�v���v��,^���~��Y������w�,��xS�g���6Ylg��b���Y>Эֲ<�� j-���]i���Vk�-������ -&
}��C�0��4�M;kh��AC��;�Pm���[�a�nq@��+��h���^iw���E�.ɬ;���~�����L���{����e-��v�}T������W-jv�}��Q���~�bFl�b�G�u���]�.Һ����1x~6}٢f�k�T��K��3�:�@��`H�>:��	�EGCx�:X�8Z�3k�}�f�ޯ%���tV�m9jC��C:�Io�Ҽiw������xC��C8�	o�xC��C7��gZ��7D�>h�:+kA�7��>���6��%��!�Մ���>d�#�,w�1N*�Ѱ�4�&��8�pc8�1��c�1������Ќ����x�{k�H�t��$�%��u�	\'��K�u��Lk� F����g���3IAq�i�濝��Z堢�Q���KHp��p�|9�H;�PU��kܝ���m��;�Jkv",�Į����=��t|���34��kl3n�X��
7
��F0����G�E~ٿ���������m���u߿Y�����������Mw���q���be�V���m�����b����~�BWS�Y4XD��ګ=�6k$�����%j��y��?�6��V>�!���o���Mt*��&���t�/{��� 3�]�����t��tW�u�ް�2��36m!`b�%Lw'l�?ck�񌁘`΄�IuH����?���m���p� (���O��MGu>3zj�Z��<�LR�g�e2Dg`$k
�;�4T3�|�jnx��M�r���rq�y����R�S6���[ݭ�E�$�\������4�O�3V|�T�Ι����m�"-�����6:Lࡂ7=R6�_~K�j�B�@o��46�O`��l�@�?���~�����O`z��m6m<FC�b�=FCK�Д�=FEK�дs�gݒA4U`�����i��DO���1M;���zn����v
�O� ������z����|��$����#c��(�1Qb�`D���/O׌:]_}���j1��lNG���5K�Le˥,'�5q�d"�5�(-P)X���6PQ	,1�2�ՎcB(�b�򲢥�є��J&�W�*����`
t��!�5j��Z�ˍj�a-��n�%xE���K�~���ո���D��Q��.���;e�cx��ķ�@xE����yف��=�@ di�NR;��x,R@���&��h"&QO�VE�μ�7H4�r9��21��92� ��o���8�G��6��K� +µ�*k��<�_�x�������Ũ<�g�)m:���� ���I��!�<�`p�:K�D,W�t�n�����h� !��(F|R�d�cv�c>*��2�VSJ'��t�}���.��ZO�'�YZ���6**�[s����y���o�ty�U �nܝ�:���e�ݡǰ�_��;%\R�g�z�\�6Wn��UP�)L�U����Y�	:[]J�9�G��C:H�aQs�@���$,�I(	|�4�A���~$��2�81La6�#�-1m�:䐂m�64��oA���m�����.g*)"��*��'������?��ϟf�t�UAy�\��0�%@`�-PLۘTJ�	�Jq/y�$a�Nӌ8		��7�2i�h�X���zv����^R���������闧�5�@JC�� ��B(�q�4ɜS���u�V���0/,}��sF�)�����O�sQhe5�!"(C�Ԗ�<�05F�EC�l��/N�&��<Ғ|��h:�;�W�4bT���<B�S&<�����<^9T��C��oX��u@u���jߏ��j��=w���!��y	��c��њKb�-]�B���GԠ��A��� ޣ@P��hU�Ҩvn.H%Dp�����=-5u�Na��w���+Ʒ�vL�A���m�צg��&`"`škl�Ϟ��7��u��|�����l<L��< ��]����y8i��ǭ%�(I%'
0:�ҝ��+I�0B�4�~I*�o�ʟx�96Bq���ڒ��r��u{�����\?�U�e5�_F��b��H8���F��(���{�r��܌�FѝwjMe�Vq_�d��g���6�k�a��tz��/�­j��O���<�?Y�5������mNM�\�poR�STY�Q�댠������f�JwC!��@�k�w9z�>���um�T�H�e�4�r"!a��&)��	�ف�������������������������������������������������V���� PK
   ��!Y
O�+.  �                  cirkitFile.jsonPK
   ��!YG�~��  � /             X.  images/0739a1b1-a163-452a-a325-ab452d55b136.pngPK
   ��!Y�R�� $� /             /�  images/179c08ce-6e18-4019-8002-932a24469ad1.pngPK
   ��!Y�;�К> � /             i� images/277be1dd-7489-4b2a-8eff-ec6391927629.pngPK
   ��!Y�H<�'  �'  /             P images/289c84f5-bee9-42dc-8a56-be82ea7098c8.pngPK
   ��!Y����7  �  /             *- images/2b66d102-ef9e-4dde-8ee7-817842500f7b.pngPK
   ��!Yh`Pҷ!  �!  /             �> images/4b60cb4e-ac73-4aba-afdc-1cf5937e57a1.pngPK
   ��!Yv��� f~ /             �` images/4d249bba-3190-4770-b321-fb8fc027a237.pngPK
   ��!Y8�Z��(  �(  /             �h images/52e5cf08-beef-4b5f-967f-8676d3f3880a.pngPK
   ��!Y����+  J  /             � images/5644ca41-1cf6-484a-bb07-c2f9a6f5b19b.pngPK
   ��!Y}�� � /             �� images/5874d651-dcf0-4a98-b8b4-9fcbfdf83d7f.pngPK
   ��!Y~��k�6 4 /             �^ images/663b53f5-e86a-4272-a51e-f5b809259b46.pngPK
   ��!Y�1.:�  )  /             �� images/8d2526ea-6e7a-4b7c-a99b-0902daeefaab.pngPK
   ��!Yu��|  w  /             �� images/907fdf8d-ea69-4713-a731-45c9eedceef3.pngPK
   ��!Y�Ƚ׌  �  /             l� images/9185dcb2-65ea-4de0-8d42-42cedb1b5634.pngPK
   ��!Y�� �f  y�  /             E� images/96fabd4d-0b16-452b-94e2-688cfcbce531.pngPK
   ��!Y�&�}[  y`  /             o9 images/982accd3-ee7b-437c-8e9e-7ebd1fcbf7fd.pngPK
   ��!Y?S��� 2� /             9� images/99226213-8268-43da-ade8-d9d07cfcec9f.pngPK
   ��!Ya6֌1!  ,!  /             m images/a0acbd77-339e-480e-a1f6-37906f79b183.pngPK
   ��!Y$�8�l  �  /             �� images/aa130aff-16e6-4627-9689-819d55b5861f.pngPK
   ��!Y+L$��� �� /             T� images/aad47697-5cf4-402f-a095-abba84463b41.pngPK
   ��!Y����<  �  /             v~ images/bdd7c0cc-86d6-4eb9-abef-3fcf444ec41a.pngPK
   ��!Y��g)�
  �
  /             �� images/c1fb8ae3-abb7-4800-a199-c8a1e0562abd.pngPK
   ��!Y���]  [  /             /� images/cbec1558-c992-4de5-91c3-4ac90e5ffec0.pngPK
   ��!Y/yR�c  ^  /             �� images/d2af519c-c065-45b5-bffd-6bf239de2b90.pngPK
   ��!Y�GDU7� �� /             1� images/d628d844-ce42-4e82-be63-f5fdfa438334.pngPK
   ��!Y�Y`�1u � /             �� images/d9bcf815-618f-4ab0-b416-9f611d86ef67.pngPK
   ��!Y~��a� ٮ /             3%! images/dc707dc6-8489-41bb-a5bc-77a0670f90d6.pngPK
   ��!Y���� =< /             ��" images/e0d827a2-ee8a-45f1-850c-b31b1c4188d2.pngPK
   ��!Y;��q p� /             ��% images/e9c16099-5161-4325-9ccd-582d4965bc31.pngPK
   ��!Y����`  [  /             d( images/fc6d97d6-a1d8-4630-b4a2-8bef38b47130.pngPK
   ��!Y����#  �               �}( jsons/user_defined.jsonPK        h  �(   